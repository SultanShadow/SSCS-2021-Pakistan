magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< nwell >>
rect -1138 -1138 1138 1138
<< pwell >>
rect -1266 1180 1266 1266
rect -1266 -1180 -1180 1180
rect 1180 -1180 1266 1180
rect -1266 -1266 1266 -1180
<< psubdiff >>
rect -1240 1206 -1139 1240
rect -1105 1206 -1071 1240
rect -1037 1206 -1003 1240
rect -969 1206 -935 1240
rect -901 1206 -867 1240
rect -833 1206 -799 1240
rect -765 1206 -731 1240
rect -697 1206 -663 1240
rect -629 1206 -595 1240
rect -561 1206 -527 1240
rect -493 1206 -459 1240
rect -425 1206 -391 1240
rect -357 1206 -323 1240
rect -289 1206 -255 1240
rect -221 1206 -187 1240
rect -153 1206 -119 1240
rect -85 1206 -51 1240
rect -17 1206 17 1240
rect 51 1206 85 1240
rect 119 1206 153 1240
rect 187 1206 221 1240
rect 255 1206 289 1240
rect 323 1206 357 1240
rect 391 1206 425 1240
rect 459 1206 493 1240
rect 527 1206 561 1240
rect 595 1206 629 1240
rect 663 1206 697 1240
rect 731 1206 765 1240
rect 799 1206 833 1240
rect 867 1206 901 1240
rect 935 1206 969 1240
rect 1003 1206 1037 1240
rect 1071 1206 1105 1240
rect 1139 1206 1240 1240
rect -1240 1139 -1206 1206
rect -1240 1071 -1206 1105
rect 1206 1139 1240 1206
rect -1240 1003 -1206 1037
rect -1240 935 -1206 969
rect -1240 867 -1206 901
rect -1240 799 -1206 833
rect -1240 731 -1206 765
rect -1240 663 -1206 697
rect -1240 595 -1206 629
rect -1240 527 -1206 561
rect -1240 459 -1206 493
rect -1240 391 -1206 425
rect -1240 323 -1206 357
rect -1240 255 -1206 289
rect -1240 187 -1206 221
rect -1240 119 -1206 153
rect -1240 51 -1206 85
rect -1240 -17 -1206 17
rect -1240 -85 -1206 -51
rect -1240 -153 -1206 -119
rect -1240 -221 -1206 -187
rect -1240 -289 -1206 -255
rect -1240 -357 -1206 -323
rect -1240 -425 -1206 -391
rect -1240 -493 -1206 -459
rect -1240 -561 -1206 -527
rect -1240 -629 -1206 -595
rect -1240 -697 -1206 -663
rect -1240 -765 -1206 -731
rect -1240 -833 -1206 -799
rect -1240 -901 -1206 -867
rect -1240 -969 -1206 -935
rect -1240 -1037 -1206 -1003
rect -1240 -1105 -1206 -1071
rect 1206 1071 1240 1105
rect 1206 1003 1240 1037
rect 1206 935 1240 969
rect 1206 867 1240 901
rect 1206 799 1240 833
rect 1206 731 1240 765
rect 1206 663 1240 697
rect 1206 595 1240 629
rect 1206 527 1240 561
rect 1206 459 1240 493
rect 1206 391 1240 425
rect 1206 323 1240 357
rect 1206 255 1240 289
rect 1206 187 1240 221
rect 1206 119 1240 153
rect 1206 51 1240 85
rect 1206 -17 1240 17
rect 1206 -85 1240 -51
rect 1206 -153 1240 -119
rect 1206 -221 1240 -187
rect 1206 -289 1240 -255
rect 1206 -357 1240 -323
rect 1206 -425 1240 -391
rect 1206 -493 1240 -459
rect 1206 -561 1240 -527
rect 1206 -629 1240 -595
rect 1206 -697 1240 -663
rect 1206 -765 1240 -731
rect 1206 -833 1240 -799
rect 1206 -901 1240 -867
rect 1206 -969 1240 -935
rect 1206 -1037 1240 -1003
rect -1240 -1206 -1206 -1139
rect 1206 -1105 1240 -1071
rect 1206 -1206 1240 -1139
rect -1240 -1240 -1139 -1206
rect -1105 -1240 -1071 -1206
rect -1037 -1240 -1003 -1206
rect -969 -1240 -935 -1206
rect -901 -1240 -867 -1206
rect -833 -1240 -799 -1206
rect -765 -1240 -731 -1206
rect -697 -1240 -663 -1206
rect -629 -1240 -595 -1206
rect -561 -1240 -527 -1206
rect -493 -1240 -459 -1206
rect -425 -1240 -391 -1206
rect -357 -1240 -323 -1206
rect -289 -1240 -255 -1206
rect -221 -1240 -187 -1206
rect -153 -1240 -119 -1206
rect -85 -1240 -51 -1206
rect -17 -1240 17 -1206
rect 51 -1240 85 -1206
rect 119 -1240 153 -1206
rect 187 -1240 221 -1206
rect 255 -1240 289 -1206
rect 323 -1240 357 -1206
rect 391 -1240 425 -1206
rect 459 -1240 493 -1206
rect 527 -1240 561 -1206
rect 595 -1240 629 -1206
rect 663 -1240 697 -1206
rect 731 -1240 765 -1206
rect 799 -1240 833 -1206
rect 867 -1240 901 -1206
rect 935 -1240 969 -1206
rect 1003 -1240 1037 -1206
rect 1071 -1240 1105 -1206
rect 1139 -1240 1240 -1206
<< nsubdiff >>
rect -1102 1068 -1003 1102
rect -969 1068 -935 1102
rect -901 1068 -867 1102
rect -833 1068 -799 1102
rect -765 1068 -731 1102
rect -697 1068 -663 1102
rect -629 1068 -595 1102
rect -561 1068 -527 1102
rect -493 1068 -459 1102
rect -425 1068 -391 1102
rect -357 1068 -323 1102
rect -289 1068 -255 1102
rect -221 1068 -187 1102
rect -153 1068 -119 1102
rect -85 1068 -51 1102
rect -17 1068 17 1102
rect 51 1068 85 1102
rect 119 1068 153 1102
rect 187 1068 221 1102
rect 255 1068 289 1102
rect 323 1068 357 1102
rect 391 1068 425 1102
rect 459 1068 493 1102
rect 527 1068 561 1102
rect 595 1068 629 1102
rect 663 1068 697 1102
rect 731 1068 765 1102
rect 799 1068 833 1102
rect 867 1068 901 1102
rect 935 1068 969 1102
rect 1003 1068 1102 1102
rect -1102 1003 -1068 1068
rect 1068 1003 1102 1068
rect -1102 935 -1068 969
rect -1102 867 -1068 901
rect -1102 799 -1068 833
rect -1102 731 -1068 765
rect -1102 663 -1068 697
rect -1102 595 -1068 629
rect -1102 527 -1068 561
rect -1102 459 -1068 493
rect -1102 391 -1068 425
rect -1102 323 -1068 357
rect -1102 255 -1068 289
rect -1102 187 -1068 221
rect -1102 119 -1068 153
rect -1102 51 -1068 85
rect -1102 -17 -1068 17
rect -1102 -85 -1068 -51
rect -1102 -153 -1068 -119
rect -1102 -221 -1068 -187
rect -1102 -289 -1068 -255
rect -1102 -357 -1068 -323
rect -1102 -425 -1068 -391
rect -1102 -493 -1068 -459
rect -1102 -561 -1068 -527
rect -1102 -629 -1068 -595
rect -1102 -697 -1068 -663
rect -1102 -765 -1068 -731
rect -1102 -833 -1068 -799
rect -1102 -901 -1068 -867
rect -1102 -969 -1068 -935
rect 1068 935 1102 969
rect 1068 867 1102 901
rect 1068 799 1102 833
rect 1068 731 1102 765
rect 1068 663 1102 697
rect 1068 595 1102 629
rect 1068 527 1102 561
rect 1068 459 1102 493
rect 1068 391 1102 425
rect 1068 323 1102 357
rect 1068 255 1102 289
rect 1068 187 1102 221
rect 1068 119 1102 153
rect 1068 51 1102 85
rect 1068 -17 1102 17
rect 1068 -85 1102 -51
rect 1068 -153 1102 -119
rect 1068 -221 1102 -187
rect 1068 -289 1102 -255
rect 1068 -357 1102 -323
rect 1068 -425 1102 -391
rect 1068 -493 1102 -459
rect 1068 -561 1102 -527
rect 1068 -629 1102 -595
rect 1068 -697 1102 -663
rect 1068 -765 1102 -731
rect 1068 -833 1102 -799
rect 1068 -901 1102 -867
rect 1068 -969 1102 -935
rect -1102 -1068 -1068 -1003
rect 1068 -1068 1102 -1003
rect -1102 -1102 -1003 -1068
rect -969 -1102 -935 -1068
rect -901 -1102 -867 -1068
rect -833 -1102 -799 -1068
rect -765 -1102 -731 -1068
rect -697 -1102 -663 -1068
rect -629 -1102 -595 -1068
rect -561 -1102 -527 -1068
rect -493 -1102 -459 -1068
rect -425 -1102 -391 -1068
rect -357 -1102 -323 -1068
rect -289 -1102 -255 -1068
rect -221 -1102 -187 -1068
rect -153 -1102 -119 -1068
rect -85 -1102 -51 -1068
rect -17 -1102 17 -1068
rect 51 -1102 85 -1068
rect 119 -1102 153 -1068
rect 187 -1102 221 -1068
rect 255 -1102 289 -1068
rect 323 -1102 357 -1068
rect 391 -1102 425 -1068
rect 459 -1102 493 -1068
rect 527 -1102 561 -1068
rect 595 -1102 629 -1068
rect 663 -1102 697 -1068
rect 731 -1102 765 -1068
rect 799 -1102 833 -1068
rect 867 -1102 901 -1068
rect 935 -1102 969 -1068
rect 1003 -1102 1102 -1068
<< psubdiffcont >>
rect -1139 1206 -1105 1240
rect -1071 1206 -1037 1240
rect -1003 1206 -969 1240
rect -935 1206 -901 1240
rect -867 1206 -833 1240
rect -799 1206 -765 1240
rect -731 1206 -697 1240
rect -663 1206 -629 1240
rect -595 1206 -561 1240
rect -527 1206 -493 1240
rect -459 1206 -425 1240
rect -391 1206 -357 1240
rect -323 1206 -289 1240
rect -255 1206 -221 1240
rect -187 1206 -153 1240
rect -119 1206 -85 1240
rect -51 1206 -17 1240
rect 17 1206 51 1240
rect 85 1206 119 1240
rect 153 1206 187 1240
rect 221 1206 255 1240
rect 289 1206 323 1240
rect 357 1206 391 1240
rect 425 1206 459 1240
rect 493 1206 527 1240
rect 561 1206 595 1240
rect 629 1206 663 1240
rect 697 1206 731 1240
rect 765 1206 799 1240
rect 833 1206 867 1240
rect 901 1206 935 1240
rect 969 1206 1003 1240
rect 1037 1206 1071 1240
rect 1105 1206 1139 1240
rect -1240 1105 -1206 1139
rect 1206 1105 1240 1139
rect -1240 1037 -1206 1071
rect -1240 969 -1206 1003
rect -1240 901 -1206 935
rect -1240 833 -1206 867
rect -1240 765 -1206 799
rect -1240 697 -1206 731
rect -1240 629 -1206 663
rect -1240 561 -1206 595
rect -1240 493 -1206 527
rect -1240 425 -1206 459
rect -1240 357 -1206 391
rect -1240 289 -1206 323
rect -1240 221 -1206 255
rect -1240 153 -1206 187
rect -1240 85 -1206 119
rect -1240 17 -1206 51
rect -1240 -51 -1206 -17
rect -1240 -119 -1206 -85
rect -1240 -187 -1206 -153
rect -1240 -255 -1206 -221
rect -1240 -323 -1206 -289
rect -1240 -391 -1206 -357
rect -1240 -459 -1206 -425
rect -1240 -527 -1206 -493
rect -1240 -595 -1206 -561
rect -1240 -663 -1206 -629
rect -1240 -731 -1206 -697
rect -1240 -799 -1206 -765
rect -1240 -867 -1206 -833
rect -1240 -935 -1206 -901
rect -1240 -1003 -1206 -969
rect -1240 -1071 -1206 -1037
rect 1206 1037 1240 1071
rect 1206 969 1240 1003
rect 1206 901 1240 935
rect 1206 833 1240 867
rect 1206 765 1240 799
rect 1206 697 1240 731
rect 1206 629 1240 663
rect 1206 561 1240 595
rect 1206 493 1240 527
rect 1206 425 1240 459
rect 1206 357 1240 391
rect 1206 289 1240 323
rect 1206 221 1240 255
rect 1206 153 1240 187
rect 1206 85 1240 119
rect 1206 17 1240 51
rect 1206 -51 1240 -17
rect 1206 -119 1240 -85
rect 1206 -187 1240 -153
rect 1206 -255 1240 -221
rect 1206 -323 1240 -289
rect 1206 -391 1240 -357
rect 1206 -459 1240 -425
rect 1206 -527 1240 -493
rect 1206 -595 1240 -561
rect 1206 -663 1240 -629
rect 1206 -731 1240 -697
rect 1206 -799 1240 -765
rect 1206 -867 1240 -833
rect 1206 -935 1240 -901
rect 1206 -1003 1240 -969
rect 1206 -1071 1240 -1037
rect -1240 -1139 -1206 -1105
rect 1206 -1139 1240 -1105
rect -1139 -1240 -1105 -1206
rect -1071 -1240 -1037 -1206
rect -1003 -1240 -969 -1206
rect -935 -1240 -901 -1206
rect -867 -1240 -833 -1206
rect -799 -1240 -765 -1206
rect -731 -1240 -697 -1206
rect -663 -1240 -629 -1206
rect -595 -1240 -561 -1206
rect -527 -1240 -493 -1206
rect -459 -1240 -425 -1206
rect -391 -1240 -357 -1206
rect -323 -1240 -289 -1206
rect -255 -1240 -221 -1206
rect -187 -1240 -153 -1206
rect -119 -1240 -85 -1206
rect -51 -1240 -17 -1206
rect 17 -1240 51 -1206
rect 85 -1240 119 -1206
rect 153 -1240 187 -1206
rect 221 -1240 255 -1206
rect 289 -1240 323 -1206
rect 357 -1240 391 -1206
rect 425 -1240 459 -1206
rect 493 -1240 527 -1206
rect 561 -1240 595 -1206
rect 629 -1240 663 -1206
rect 697 -1240 731 -1206
rect 765 -1240 799 -1206
rect 833 -1240 867 -1206
rect 901 -1240 935 -1206
rect 969 -1240 1003 -1206
rect 1037 -1240 1071 -1206
rect 1105 -1240 1139 -1206
<< nsubdiffcont >>
rect -1003 1068 -969 1102
rect -935 1068 -901 1102
rect -867 1068 -833 1102
rect -799 1068 -765 1102
rect -731 1068 -697 1102
rect -663 1068 -629 1102
rect -595 1068 -561 1102
rect -527 1068 -493 1102
rect -459 1068 -425 1102
rect -391 1068 -357 1102
rect -323 1068 -289 1102
rect -255 1068 -221 1102
rect -187 1068 -153 1102
rect -119 1068 -85 1102
rect -51 1068 -17 1102
rect 17 1068 51 1102
rect 85 1068 119 1102
rect 153 1068 187 1102
rect 221 1068 255 1102
rect 289 1068 323 1102
rect 357 1068 391 1102
rect 425 1068 459 1102
rect 493 1068 527 1102
rect 561 1068 595 1102
rect 629 1068 663 1102
rect 697 1068 731 1102
rect 765 1068 799 1102
rect 833 1068 867 1102
rect 901 1068 935 1102
rect 969 1068 1003 1102
rect -1102 969 -1068 1003
rect -1102 901 -1068 935
rect -1102 833 -1068 867
rect -1102 765 -1068 799
rect -1102 697 -1068 731
rect -1102 629 -1068 663
rect -1102 561 -1068 595
rect -1102 493 -1068 527
rect -1102 425 -1068 459
rect -1102 357 -1068 391
rect -1102 289 -1068 323
rect -1102 221 -1068 255
rect -1102 153 -1068 187
rect -1102 85 -1068 119
rect -1102 17 -1068 51
rect -1102 -51 -1068 -17
rect -1102 -119 -1068 -85
rect -1102 -187 -1068 -153
rect -1102 -255 -1068 -221
rect -1102 -323 -1068 -289
rect -1102 -391 -1068 -357
rect -1102 -459 -1068 -425
rect -1102 -527 -1068 -493
rect -1102 -595 -1068 -561
rect -1102 -663 -1068 -629
rect -1102 -731 -1068 -697
rect -1102 -799 -1068 -765
rect -1102 -867 -1068 -833
rect -1102 -935 -1068 -901
rect -1102 -1003 -1068 -969
rect 1068 969 1102 1003
rect 1068 901 1102 935
rect 1068 833 1102 867
rect 1068 765 1102 799
rect 1068 697 1102 731
rect 1068 629 1102 663
rect 1068 561 1102 595
rect 1068 493 1102 527
rect 1068 425 1102 459
rect 1068 357 1102 391
rect 1068 289 1102 323
rect 1068 221 1102 255
rect 1068 153 1102 187
rect 1068 85 1102 119
rect 1068 17 1102 51
rect 1068 -51 1102 -17
rect 1068 -119 1102 -85
rect 1068 -187 1102 -153
rect 1068 -255 1102 -221
rect 1068 -323 1102 -289
rect 1068 -391 1102 -357
rect 1068 -459 1102 -425
rect 1068 -527 1102 -493
rect 1068 -595 1102 -561
rect 1068 -663 1102 -629
rect 1068 -731 1102 -697
rect 1068 -799 1102 -765
rect 1068 -867 1102 -833
rect 1068 -935 1102 -901
rect 1068 -1003 1102 -969
rect -1003 -1102 -969 -1068
rect -935 -1102 -901 -1068
rect -867 -1102 -833 -1068
rect -799 -1102 -765 -1068
rect -731 -1102 -697 -1068
rect -663 -1102 -629 -1068
rect -595 -1102 -561 -1068
rect -527 -1102 -493 -1068
rect -459 -1102 -425 -1068
rect -391 -1102 -357 -1068
rect -323 -1102 -289 -1068
rect -255 -1102 -221 -1068
rect -187 -1102 -153 -1068
rect -119 -1102 -85 -1068
rect -51 -1102 -17 -1068
rect 17 -1102 51 -1068
rect 85 -1102 119 -1068
rect 153 -1102 187 -1068
rect 221 -1102 255 -1068
rect 289 -1102 323 -1068
rect 357 -1102 391 -1068
rect 425 -1102 459 -1068
rect 493 -1102 527 -1068
rect 561 -1102 595 -1068
rect 629 -1102 663 -1068
rect 697 -1102 731 -1068
rect 765 -1102 799 -1068
rect 833 -1102 867 -1068
rect 901 -1102 935 -1068
rect 969 -1102 1003 -1068
<< pdiode >>
rect -1000 969 1000 1000
rect -1000 -969 -969 969
rect 969 -969 1000 969
rect -1000 -1000 1000 -969
<< pdiodec >>
rect -969 -969 969 969
<< locali >>
rect -1240 1206 -1139 1240
rect -1105 1206 -1071 1240
rect -1037 1206 -1003 1240
rect -969 1206 -935 1240
rect -901 1206 -867 1240
rect -833 1206 -799 1240
rect -765 1206 -731 1240
rect -697 1206 -663 1240
rect -629 1206 -595 1240
rect -561 1206 -527 1240
rect -493 1206 -459 1240
rect -425 1206 -391 1240
rect -357 1206 -323 1240
rect -289 1206 -255 1240
rect -221 1206 -187 1240
rect -153 1206 -119 1240
rect -85 1206 -51 1240
rect -17 1206 17 1240
rect 51 1206 85 1240
rect 119 1206 153 1240
rect 187 1206 221 1240
rect 255 1206 289 1240
rect 323 1206 357 1240
rect 391 1206 425 1240
rect 459 1206 493 1240
rect 527 1206 561 1240
rect 595 1206 629 1240
rect 663 1206 697 1240
rect 731 1206 765 1240
rect 799 1206 833 1240
rect 867 1206 901 1240
rect 935 1206 969 1240
rect 1003 1206 1037 1240
rect 1071 1206 1105 1240
rect 1139 1206 1240 1240
rect -1240 1139 -1206 1206
rect -1240 1071 -1206 1105
rect 1206 1139 1240 1206
rect -1240 1003 -1206 1037
rect -1240 935 -1206 969
rect -1240 867 -1206 901
rect -1240 799 -1206 833
rect -1240 731 -1206 765
rect -1240 663 -1206 697
rect -1240 595 -1206 629
rect -1240 527 -1206 561
rect -1240 459 -1206 493
rect -1240 391 -1206 425
rect -1240 323 -1206 357
rect -1240 255 -1206 289
rect -1240 187 -1206 221
rect -1240 119 -1206 153
rect -1240 51 -1206 85
rect -1240 -17 -1206 17
rect -1240 -85 -1206 -51
rect -1240 -153 -1206 -119
rect -1240 -221 -1206 -187
rect -1240 -289 -1206 -255
rect -1240 -357 -1206 -323
rect -1240 -425 -1206 -391
rect -1240 -493 -1206 -459
rect -1240 -561 -1206 -527
rect -1240 -629 -1206 -595
rect -1240 -697 -1206 -663
rect -1240 -765 -1206 -731
rect -1240 -833 -1206 -799
rect -1240 -901 -1206 -867
rect -1240 -969 -1206 -935
rect -1240 -1037 -1206 -1003
rect -1240 -1105 -1206 -1071
rect -1102 1068 -1003 1102
rect -969 1068 -935 1102
rect -901 1068 -867 1102
rect -833 1068 -799 1102
rect -765 1068 -731 1102
rect -697 1068 -663 1102
rect -629 1068 -595 1102
rect -561 1068 -527 1102
rect -493 1068 -459 1102
rect -425 1068 -391 1102
rect -357 1068 -323 1102
rect -289 1068 -255 1102
rect -221 1068 -187 1102
rect -153 1068 -119 1102
rect -85 1068 -51 1102
rect -17 1068 17 1102
rect 51 1068 85 1102
rect 119 1068 153 1102
rect 187 1068 221 1102
rect 255 1068 289 1102
rect 323 1068 357 1102
rect 391 1068 425 1102
rect 459 1068 493 1102
rect 527 1068 561 1102
rect 595 1068 629 1102
rect 663 1068 697 1102
rect 731 1068 765 1102
rect 799 1068 833 1102
rect 867 1068 901 1102
rect 935 1068 969 1102
rect 1003 1068 1102 1102
rect -1102 1003 -1068 1068
rect 1068 1003 1102 1068
rect -1102 935 -1068 969
rect -1102 867 -1068 901
rect -1102 799 -1068 833
rect -1102 731 -1068 765
rect -1102 663 -1068 697
rect -1102 595 -1068 629
rect -1102 527 -1068 561
rect -1102 459 -1068 493
rect -1102 391 -1068 425
rect -1102 323 -1068 357
rect -1102 255 -1068 289
rect -1102 187 -1068 221
rect -1102 119 -1068 153
rect -1102 51 -1068 85
rect -1102 -17 -1068 17
rect -1102 -85 -1068 -51
rect -1102 -153 -1068 -119
rect -1102 -221 -1068 -187
rect -1102 -289 -1068 -255
rect -1102 -357 -1068 -323
rect -1102 -425 -1068 -391
rect -1102 -493 -1068 -459
rect -1102 -561 -1068 -527
rect -1102 -629 -1068 -595
rect -1102 -697 -1068 -663
rect -1102 -765 -1068 -731
rect -1102 -833 -1068 -799
rect -1102 -901 -1068 -867
rect -1102 -969 -1068 -935
rect -1004 969 1004 988
rect -1004 -969 -969 969
rect 969 -969 1004 969
rect -1004 -988 1004 -969
rect 1068 935 1102 969
rect 1068 867 1102 901
rect 1068 799 1102 833
rect 1068 731 1102 765
rect 1068 663 1102 697
rect 1068 595 1102 629
rect 1068 527 1102 561
rect 1068 459 1102 493
rect 1068 391 1102 425
rect 1068 323 1102 357
rect 1068 255 1102 289
rect 1068 187 1102 221
rect 1068 119 1102 153
rect 1068 51 1102 85
rect 1068 -17 1102 17
rect 1068 -85 1102 -51
rect 1068 -153 1102 -119
rect 1068 -221 1102 -187
rect 1068 -289 1102 -255
rect 1068 -357 1102 -323
rect 1068 -425 1102 -391
rect 1068 -493 1102 -459
rect 1068 -561 1102 -527
rect 1068 -629 1102 -595
rect 1068 -697 1102 -663
rect 1068 -765 1102 -731
rect 1068 -833 1102 -799
rect 1068 -901 1102 -867
rect 1068 -969 1102 -935
rect -1102 -1068 -1068 -1003
rect 1068 -1068 1102 -1003
rect -1102 -1102 -1003 -1068
rect -969 -1102 -935 -1068
rect -901 -1102 -867 -1068
rect -833 -1102 -799 -1068
rect -765 -1102 -731 -1068
rect -697 -1102 -663 -1068
rect -629 -1102 -595 -1068
rect -561 -1102 -527 -1068
rect -493 -1102 -459 -1068
rect -425 -1102 -391 -1068
rect -357 -1102 -323 -1068
rect -289 -1102 -255 -1068
rect -221 -1102 -187 -1068
rect -153 -1102 -119 -1068
rect -85 -1102 -51 -1068
rect -17 -1102 17 -1068
rect 51 -1102 85 -1068
rect 119 -1102 153 -1068
rect 187 -1102 221 -1068
rect 255 -1102 289 -1068
rect 323 -1102 357 -1068
rect 391 -1102 425 -1068
rect 459 -1102 493 -1068
rect 527 -1102 561 -1068
rect 595 -1102 629 -1068
rect 663 -1102 697 -1068
rect 731 -1102 765 -1068
rect 799 -1102 833 -1068
rect 867 -1102 901 -1068
rect 935 -1102 969 -1068
rect 1003 -1102 1102 -1068
rect 1206 1071 1240 1105
rect 1206 1003 1240 1037
rect 1206 935 1240 969
rect 1206 867 1240 901
rect 1206 799 1240 833
rect 1206 731 1240 765
rect 1206 663 1240 697
rect 1206 595 1240 629
rect 1206 527 1240 561
rect 1206 459 1240 493
rect 1206 391 1240 425
rect 1206 323 1240 357
rect 1206 255 1240 289
rect 1206 187 1240 221
rect 1206 119 1240 153
rect 1206 51 1240 85
rect 1206 -17 1240 17
rect 1206 -85 1240 -51
rect 1206 -153 1240 -119
rect 1206 -221 1240 -187
rect 1206 -289 1240 -255
rect 1206 -357 1240 -323
rect 1206 -425 1240 -391
rect 1206 -493 1240 -459
rect 1206 -561 1240 -527
rect 1206 -629 1240 -595
rect 1206 -697 1240 -663
rect 1206 -765 1240 -731
rect 1206 -833 1240 -799
rect 1206 -901 1240 -867
rect 1206 -969 1240 -935
rect 1206 -1037 1240 -1003
rect -1240 -1206 -1206 -1139
rect 1206 -1105 1240 -1071
rect 1206 -1206 1240 -1139
rect -1240 -1240 -1139 -1206
rect -1105 -1240 -1071 -1206
rect -1037 -1240 -1003 -1206
rect -969 -1240 -935 -1206
rect -901 -1240 -867 -1206
rect -833 -1240 -799 -1206
rect -765 -1240 -731 -1206
rect -697 -1240 -663 -1206
rect -629 -1240 -595 -1206
rect -561 -1240 -527 -1206
rect -493 -1240 -459 -1206
rect -425 -1240 -391 -1206
rect -357 -1240 -323 -1206
rect -289 -1240 -255 -1206
rect -221 -1240 -187 -1206
rect -153 -1240 -119 -1206
rect -85 -1240 -51 -1206
rect -17 -1240 17 -1206
rect 51 -1240 85 -1206
rect 119 -1240 153 -1206
rect 187 -1240 221 -1206
rect 255 -1240 289 -1206
rect 323 -1240 357 -1206
rect 391 -1240 425 -1206
rect 459 -1240 493 -1206
rect 527 -1240 561 -1206
rect 595 -1240 629 -1206
rect 663 -1240 697 -1206
rect 731 -1240 765 -1206
rect 799 -1240 833 -1206
rect 867 -1240 901 -1206
rect 935 -1240 969 -1206
rect 1003 -1240 1037 -1206
rect 1071 -1240 1105 -1206
rect 1139 -1240 1240 -1206
<< viali >>
rect -953 -953 953 953
<< metal1 >>
rect -1000 953 1000 994
rect -1000 -953 -953 953
rect 953 -953 1000 953
rect -1000 -994 1000 -953
<< properties >>
string FIXED_BBOX -1084 -1084 1084 1084
<< end >>
