magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< nwell >>
rect 495004 678715 495325 678813
rect 495092 678711 495257 678715
<< nsubdiff >>
rect 495090 678761 495261 678776
rect 495090 678727 495124 678761
rect 495158 678727 495192 678761
rect 495226 678727 495261 678761
rect 495090 678711 495261 678727
<< nsubdiffcont >>
rect 495124 678727 495158 678761
rect 495192 678727 495226 678761
<< locali >>
rect 386438 693286 386473 693315
rect 386472 693252 386473 693286
rect 386438 693214 386473 693252
rect 386472 693180 386473 693214
rect 386438 693142 386473 693180
rect 386472 693108 386473 693142
rect 386438 693070 386473 693108
rect 386472 693036 386473 693070
rect 386438 692998 386473 693036
rect 386472 692964 386473 692998
rect 386438 692926 386473 692964
rect 386472 692892 386473 692926
rect 386438 692854 386473 692892
rect 386472 692820 386473 692854
rect 386438 692782 386473 692820
rect 386472 692748 386473 692782
rect 386438 692710 386473 692748
rect 386472 692676 386473 692710
rect 386438 692638 386473 692676
rect 386472 692604 386473 692638
rect 386438 692566 386473 692604
rect 386472 692532 386473 692566
rect 386438 692494 386473 692532
rect 386472 692460 386473 692494
rect 386438 692431 386473 692460
rect 386904 691893 386918 691927
rect 386952 691893 386990 691927
rect 387024 691893 387062 691927
rect 387096 691893 387134 691927
rect 387168 691893 387206 691927
rect 387240 691893 387278 691927
rect 387312 691893 387350 691927
rect 387384 691893 387422 691927
rect 387456 691893 387494 691927
rect 387528 691893 387566 691927
rect 387600 691893 387638 691927
rect 387672 691893 387710 691927
rect 387744 691893 387759 691927
rect 497271 684314 501426 687895
rect 501727 685586 502104 685587
rect 501727 685552 501754 685586
rect 501788 685552 501826 685586
rect 501860 685552 501898 685586
rect 501932 685552 501970 685586
rect 502004 685552 502042 685586
rect 502076 685552 502104 685586
rect 495429 681011 495463 681041
rect 495429 680939 495463 680977
rect 495429 680867 495463 680905
rect 495429 680795 495463 680833
rect 495429 680723 495463 680761
rect 495429 680651 495463 680689
rect 495429 680579 495463 680617
rect 495429 680515 495463 680545
rect 496918 680454 497874 681038
rect 495092 678761 495257 678776
rect 495092 678727 495122 678761
rect 495158 678727 495192 678761
rect 495228 678727 495257 678761
rect 495092 678711 495257 678727
rect 513146 665566 513180 665598
rect 513146 665494 513180 665532
rect 513146 665422 513180 665460
rect 513146 665350 513180 665388
rect 513146 665278 513180 665316
rect 513146 665206 513180 665244
rect 513146 665134 513180 665172
rect 513146 665062 513180 665100
rect 513146 664990 513180 665028
rect 513146 664918 513180 664956
rect 513146 664846 513180 664884
rect 513146 664774 513180 664812
rect 513146 664702 513180 664740
rect 513146 664630 513180 664668
rect 513146 664558 513180 664596
rect 513146 664486 513180 664524
rect 513146 664414 513180 664452
rect 513146 664342 513180 664380
rect 513146 664270 513180 664308
rect 513146 664198 513180 664236
rect 513146 664126 513180 664164
rect 513146 664054 513180 664092
rect 513146 663982 513180 664020
rect 513146 663910 513180 663948
rect 513146 663838 513180 663876
rect 515592 664904 515626 664938
rect 515592 664832 515626 664870
rect 515592 664760 515626 664798
rect 515592 664688 515626 664726
rect 515592 664616 515626 664654
rect 515592 664544 515626 664582
rect 515592 664472 515626 664510
rect 515592 664400 515626 664438
rect 515592 664328 515626 664366
rect 515592 664256 515626 664294
rect 515592 664184 515626 664222
rect 515592 664112 515626 664150
rect 515592 664040 515626 664078
rect 515592 663968 515626 664006
rect 515592 663896 515626 663934
rect 515592 663828 515626 663862
rect 525120 664902 525154 664936
rect 525120 664830 525154 664868
rect 525120 664758 525154 664796
rect 525120 664686 525154 664724
rect 525120 664614 525154 664652
rect 525120 664542 525154 664580
rect 525120 664470 525154 664508
rect 525120 664398 525154 664436
rect 525120 664326 525154 664364
rect 525120 664254 525154 664292
rect 525120 664182 525154 664220
rect 525120 664110 525154 664148
rect 525120 664038 525154 664076
rect 525120 663966 525154 664004
rect 525120 663894 525154 663932
rect 525120 663826 525154 663860
rect 513146 663766 513180 663804
rect 513146 663694 513180 663732
rect 513146 663622 513180 663660
rect 513146 663557 513180 663588
rect 513854 663499 513861 663533
rect 513895 663499 513933 663533
rect 513967 663499 514005 663533
rect 514039 663499 514077 663533
rect 514111 663499 514149 663533
rect 514183 663499 514221 663533
rect 514255 663499 514293 663533
rect 514327 663499 514365 663533
rect 514399 663499 514437 663533
rect 514471 663499 514509 663533
rect 514543 663499 514581 663533
rect 514615 663499 514653 663533
rect 514687 663499 514725 663533
rect 514759 663499 514797 663533
rect 514831 663499 514838 663533
rect 525553 663081 525588 663115
rect 525622 663081 525660 663115
rect 525694 663081 525732 663115
rect 525766 663081 525804 663115
rect 525838 663081 525876 663115
rect 525910 663081 525948 663115
rect 525982 663081 526020 663115
rect 526054 663081 526092 663115
rect 526126 663081 526164 663115
rect 526198 663081 526236 663115
rect 526270 663081 526308 663115
rect 526342 663081 526380 663115
rect 526414 663081 526452 663115
rect 526486 663081 526524 663115
rect 526558 663081 526596 663115
rect 526630 663081 526668 663115
rect 526702 663081 526740 663115
rect 526774 663081 526810 663115
rect 388162 661263 388163 661297
rect 388197 661263 388235 661297
rect 388269 661263 388307 661297
rect 388341 661263 388379 661297
rect 388413 661263 388451 661297
rect 388485 661263 388523 661297
rect 388557 661263 388595 661297
rect 388629 661263 388667 661297
rect 388701 661263 388739 661297
rect 388773 661263 388811 661297
rect 388845 661263 388883 661297
rect 388917 661263 388955 661297
rect 388989 661263 388991 661297
rect 387303 660801 387337 660821
rect 387303 660729 387337 660767
rect 387303 660657 387337 660695
rect 387303 660585 387337 660623
rect 387303 660513 387337 660551
rect 387303 660441 387337 660479
rect 387303 660369 387337 660407
rect 387303 660297 387337 660335
rect 387303 660225 387337 660263
rect 387303 660153 387337 660191
rect 387303 660081 387337 660119
rect 387303 660009 387337 660047
rect 387303 659937 387337 659975
rect 387303 659865 387337 659903
rect 387303 659793 387337 659831
rect 387303 659721 387337 659759
rect 387303 659649 387337 659687
rect 468615 660203 468649 660227
rect 468615 660131 468649 660169
rect 468615 660059 468649 660097
rect 468615 659987 468649 660025
rect 468615 659915 468649 659953
rect 468615 659843 468649 659881
rect 468615 659771 468649 659809
rect 468615 659699 468649 659737
rect 468615 659642 468649 659665
rect 387303 659577 387337 659615
rect 387303 659505 387337 659543
rect 387303 659433 387337 659471
rect 387303 659361 387337 659399
rect 387303 659289 387337 659327
rect 387303 659217 387337 659255
rect 387303 659163 387337 659183
rect 497802 654106 497836 654131
rect 497802 654034 497836 654072
rect 497802 653962 497836 654000
rect 497802 653890 497836 653928
rect 497802 653818 497836 653856
rect 497802 653746 497836 653784
rect 497802 653674 497836 653712
rect 497802 653616 497836 653640
rect 496889 653382 496907 653416
rect 496941 653382 496979 653416
rect 497013 653382 497051 653416
rect 497085 653382 497123 653416
rect 497157 653382 497195 653416
rect 497229 653382 497267 653416
rect 497301 653382 497339 653416
rect 497373 653382 497411 653416
rect 497445 653382 497464 653416
rect 392043 652012 392059 652046
rect 392093 652012 392131 652046
rect 392165 652012 392203 652046
rect 392237 652012 392275 652046
rect 392309 652012 392347 652046
rect 392381 652012 392419 652046
rect 392453 652012 392491 652046
rect 392525 652012 392563 652046
rect 392597 652012 392635 652046
rect 392669 652012 392707 652046
rect 392741 652012 392779 652046
rect 392813 652012 392851 652046
rect 392885 652012 392923 652046
rect 392957 652012 392995 652046
rect 393029 652012 393067 652046
rect 393101 652012 393139 652046
rect 393173 652012 393211 652046
rect 393245 652012 393283 652046
rect 393317 652012 393355 652046
rect 393389 652012 393427 652046
rect 393461 652012 393499 652046
rect 393533 652012 393571 652046
rect 393605 652012 393622 652046
rect 391648 651451 391682 651478
rect 391648 651379 391682 651417
rect 391648 651307 391682 651345
rect 391648 651235 391682 651273
rect 391648 651163 391682 651201
rect 391648 651091 391682 651129
rect 391648 651019 391682 651057
rect 391648 650947 391682 650985
rect 391648 650875 391682 650913
rect 391648 650803 391682 650841
rect 391648 650731 391682 650769
rect 391648 650659 391682 650697
rect 391648 650587 391682 650625
rect 391648 650515 391682 650553
rect 391648 650443 391682 650481
rect 391648 650371 391682 650409
rect 391648 650299 391682 650337
rect 391648 650238 391682 650265
<< viali >>
rect 386438 693252 386472 693286
rect 386438 693180 386472 693214
rect 386438 693108 386472 693142
rect 386438 693036 386472 693070
rect 386438 692964 386472 692998
rect 386438 692892 386472 692926
rect 386438 692820 386472 692854
rect 386438 692748 386472 692782
rect 386438 692676 386472 692710
rect 386438 692604 386472 692638
rect 386438 692532 386472 692566
rect 386438 692460 386472 692494
rect 386918 691893 386952 691927
rect 386990 691893 387024 691927
rect 387062 691893 387096 691927
rect 387134 691893 387168 691927
rect 387206 691893 387240 691927
rect 387278 691893 387312 691927
rect 387350 691893 387384 691927
rect 387422 691893 387456 691927
rect 387494 691893 387528 691927
rect 387566 691893 387600 691927
rect 387638 691893 387672 691927
rect 387710 691893 387744 691927
rect 501754 685552 501788 685586
rect 501826 685552 501860 685586
rect 501898 685552 501932 685586
rect 501970 685552 502004 685586
rect 502042 685552 502076 685586
rect 495429 680977 495463 681011
rect 495429 680905 495463 680939
rect 495429 680833 495463 680867
rect 495429 680761 495463 680795
rect 495429 680689 495463 680723
rect 495429 680617 495463 680651
rect 495429 680545 495463 680579
rect 495122 678727 495124 678761
rect 495124 678727 495156 678761
rect 495194 678727 495226 678761
rect 495226 678727 495228 678761
rect 513146 665532 513180 665566
rect 513146 665460 513180 665494
rect 513146 665388 513180 665422
rect 513146 665316 513180 665350
rect 513146 665244 513180 665278
rect 513146 665172 513180 665206
rect 513146 665100 513180 665134
rect 513146 665028 513180 665062
rect 513146 664956 513180 664990
rect 513146 664884 513180 664918
rect 513146 664812 513180 664846
rect 513146 664740 513180 664774
rect 513146 664668 513180 664702
rect 513146 664596 513180 664630
rect 513146 664524 513180 664558
rect 513146 664452 513180 664486
rect 513146 664380 513180 664414
rect 513146 664308 513180 664342
rect 513146 664236 513180 664270
rect 513146 664164 513180 664198
rect 513146 664092 513180 664126
rect 513146 664020 513180 664054
rect 513146 663948 513180 663982
rect 513146 663876 513180 663910
rect 513146 663804 513180 663838
rect 515592 664870 515626 664904
rect 515592 664798 515626 664832
rect 515592 664726 515626 664760
rect 515592 664654 515626 664688
rect 515592 664582 515626 664616
rect 515592 664510 515626 664544
rect 515592 664438 515626 664472
rect 515592 664366 515626 664400
rect 515592 664294 515626 664328
rect 515592 664222 515626 664256
rect 515592 664150 515626 664184
rect 515592 664078 515626 664112
rect 515592 664006 515626 664040
rect 515592 663934 515626 663968
rect 515592 663862 515626 663896
rect 525120 664868 525154 664902
rect 525120 664796 525154 664830
rect 525120 664724 525154 664758
rect 525120 664652 525154 664686
rect 525120 664580 525154 664614
rect 525120 664508 525154 664542
rect 525120 664436 525154 664470
rect 525120 664364 525154 664398
rect 525120 664292 525154 664326
rect 525120 664220 525154 664254
rect 525120 664148 525154 664182
rect 525120 664076 525154 664110
rect 525120 664004 525154 664038
rect 525120 663932 525154 663966
rect 525120 663860 525154 663894
rect 513146 663732 513180 663766
rect 513146 663660 513180 663694
rect 513146 663588 513180 663622
rect 513861 663499 513895 663533
rect 513933 663499 513967 663533
rect 514005 663499 514039 663533
rect 514077 663499 514111 663533
rect 514149 663499 514183 663533
rect 514221 663499 514255 663533
rect 514293 663499 514327 663533
rect 514365 663499 514399 663533
rect 514437 663499 514471 663533
rect 514509 663499 514543 663533
rect 514581 663499 514615 663533
rect 514653 663499 514687 663533
rect 514725 663499 514759 663533
rect 514797 663499 514831 663533
rect 525588 663081 525622 663115
rect 525660 663081 525694 663115
rect 525732 663081 525766 663115
rect 525804 663081 525838 663115
rect 525876 663081 525910 663115
rect 525948 663081 525982 663115
rect 526020 663081 526054 663115
rect 526092 663081 526126 663115
rect 526164 663081 526198 663115
rect 526236 663081 526270 663115
rect 526308 663081 526342 663115
rect 526380 663081 526414 663115
rect 526452 663081 526486 663115
rect 526524 663081 526558 663115
rect 526596 663081 526630 663115
rect 526668 663081 526702 663115
rect 526740 663081 526774 663115
rect 388163 661263 388197 661297
rect 388235 661263 388269 661297
rect 388307 661263 388341 661297
rect 388379 661263 388413 661297
rect 388451 661263 388485 661297
rect 388523 661263 388557 661297
rect 388595 661263 388629 661297
rect 388667 661263 388701 661297
rect 388739 661263 388773 661297
rect 388811 661263 388845 661297
rect 388883 661263 388917 661297
rect 388955 661263 388989 661297
rect 387303 660767 387337 660801
rect 387303 660695 387337 660729
rect 387303 660623 387337 660657
rect 387303 660551 387337 660585
rect 387303 660479 387337 660513
rect 387303 660407 387337 660441
rect 387303 660335 387337 660369
rect 387303 660263 387337 660297
rect 387303 660191 387337 660225
rect 387303 660119 387337 660153
rect 387303 660047 387337 660081
rect 387303 659975 387337 660009
rect 387303 659903 387337 659937
rect 387303 659831 387337 659865
rect 387303 659759 387337 659793
rect 387303 659687 387337 659721
rect 387303 659615 387337 659649
rect 468615 660169 468649 660203
rect 468615 660097 468649 660131
rect 468615 660025 468649 660059
rect 468615 659953 468649 659987
rect 468615 659881 468649 659915
rect 468615 659809 468649 659843
rect 468615 659737 468649 659771
rect 468615 659665 468649 659699
rect 387303 659543 387337 659577
rect 387303 659471 387337 659505
rect 387303 659399 387337 659433
rect 387303 659327 387337 659361
rect 387303 659255 387337 659289
rect 387303 659183 387337 659217
rect 497802 654072 497836 654106
rect 497802 654000 497836 654034
rect 497802 653928 497836 653962
rect 497802 653856 497836 653890
rect 497802 653784 497836 653818
rect 497802 653712 497836 653746
rect 497802 653640 497836 653674
rect 496907 653382 496941 653416
rect 496979 653382 497013 653416
rect 497051 653382 497085 653416
rect 497123 653382 497157 653416
rect 497195 653382 497229 653416
rect 497267 653382 497301 653416
rect 497339 653382 497373 653416
rect 497411 653382 497445 653416
rect 392059 652012 392093 652046
rect 392131 652012 392165 652046
rect 392203 652012 392237 652046
rect 392275 652012 392309 652046
rect 392347 652012 392381 652046
rect 392419 652012 392453 652046
rect 392491 652012 392525 652046
rect 392563 652012 392597 652046
rect 392635 652012 392669 652046
rect 392707 652012 392741 652046
rect 392779 652012 392813 652046
rect 392851 652012 392885 652046
rect 392923 652012 392957 652046
rect 392995 652012 393029 652046
rect 393067 652012 393101 652046
rect 393139 652012 393173 652046
rect 393211 652012 393245 652046
rect 393283 652012 393317 652046
rect 393355 652012 393389 652046
rect 393427 652012 393461 652046
rect 393499 652012 393533 652046
rect 393571 652012 393605 652046
rect 391648 651417 391682 651451
rect 391648 651345 391682 651379
rect 391648 651273 391682 651307
rect 391648 651201 391682 651235
rect 391648 651129 391682 651163
rect 391648 651057 391682 651091
rect 391648 650985 391682 651019
rect 391648 650913 391682 650947
rect 391648 650841 391682 650875
rect 391648 650769 391682 650803
rect 391648 650697 391682 650731
rect 391648 650625 391682 650659
rect 391648 650553 391682 650587
rect 391648 650481 391682 650515
rect 391648 650409 391682 650443
rect 391648 650337 391682 650371
rect 391648 650265 391682 650299
<< metal1 >>
rect 386812 693765 388530 693796
rect 384496 693286 386501 693410
rect 384496 693252 386438 693286
rect 386472 693252 386501 693286
rect 384496 693214 386501 693252
rect 384496 693180 386438 693214
rect 386472 693180 386501 693214
rect 384496 693142 386501 693180
rect 384496 693108 386438 693142
rect 386472 693108 386501 693142
rect 384496 693070 386501 693108
rect 384496 693036 386438 693070
rect 386472 693036 386501 693070
rect 384496 692998 386501 693036
rect 384496 692964 386438 692998
rect 386472 692964 386501 692998
rect 384496 692926 386501 692964
rect 384496 692892 386438 692926
rect 386472 692892 386501 692926
rect 384496 692854 386501 692892
rect 384496 692820 386438 692854
rect 386472 692820 386501 692854
rect 384496 692782 386501 692820
rect 384496 692748 386438 692782
rect 386472 692748 386501 692782
rect 384496 692710 386501 692748
rect 384496 692676 386438 692710
rect 386472 692676 386501 692710
rect 384496 692638 386501 692676
rect 384496 692604 386438 692638
rect 386472 692604 386501 692638
rect 384496 692566 386501 692604
rect 384496 692532 386438 692566
rect 386472 692532 386501 692566
rect 384496 692494 386501 692532
rect 384496 692460 386438 692494
rect 386472 692460 386501 692494
rect 384496 692337 386501 692460
rect 384501 689979 386112 692337
rect 386812 692241 386813 693765
rect 388529 692241 388530 693765
rect 386812 692210 388530 692241
rect 386877 691927 387795 691941
rect 386877 691893 386918 691927
rect 386952 691893 386990 691927
rect 387024 691893 387062 691927
rect 387096 691893 387134 691927
rect 387168 691893 387206 691927
rect 387240 691893 387278 691927
rect 387312 691893 387350 691927
rect 387384 691893 387422 691927
rect 387456 691893 387494 691927
rect 387528 691893 387566 691927
rect 387600 691893 387638 691927
rect 387672 691893 387710 691927
rect 387744 691893 387795 691927
rect 386877 691147 387795 691893
rect 386877 690647 386992 691147
rect 387684 690647 387795 691147
rect 386877 690544 387795 690647
rect 83736 684024 479386 689979
rect 501821 687114 503448 687146
rect 501821 685846 501840 687114
rect 503428 685846 503448 687114
rect 501821 685815 503448 685846
rect 501704 685586 502133 685598
rect 501704 685552 501754 685586
rect 501788 685552 501826 685586
rect 501860 685552 501898 685586
rect 501932 685552 501970 685586
rect 502004 685552 502042 685586
rect 502076 685552 502133 685586
rect 501704 685157 502133 685552
rect 501704 684657 501807 685157
rect 502051 684657 502133 685157
rect 501704 684549 502133 684657
rect 380201 660899 384017 684024
rect 494064 681011 495475 681064
rect 494064 680977 495429 681011
rect 495463 680977 495475 681011
rect 494064 680954 495475 680977
rect 494064 680582 494238 680954
rect 494994 680939 495475 680954
rect 494994 680905 495429 680939
rect 495463 680905 495475 680939
rect 494994 680867 495475 680905
rect 494994 680833 495429 680867
rect 495463 680833 495475 680867
rect 494994 680795 495475 680833
rect 494994 680761 495429 680795
rect 495463 680761 495475 680795
rect 494994 680723 495475 680761
rect 494994 680689 495429 680723
rect 495463 680689 495475 680723
rect 494994 680651 495475 680689
rect 494994 680617 495429 680651
rect 495463 680617 495475 680651
rect 494994 680582 495475 680617
rect 494064 680579 495475 680582
rect 494064 680545 495429 680579
rect 495463 680545 495475 680579
rect 494064 680482 495475 680545
rect 495836 679090 496546 681114
rect 494993 678761 495260 678803
rect 494993 678727 495122 678761
rect 495156 678727 495194 678761
rect 495228 678727 495260 678761
rect 494993 678687 495260 678727
rect 466924 672500 467910 672501
rect 466924 672377 467917 672500
rect 466924 671109 467069 672377
rect 467761 671109 467917 672377
rect 466924 671001 467917 671109
rect 388119 667233 389052 667405
rect 388119 666413 388233 667233
rect 388925 666413 389052 667233
rect 388119 664360 389052 666413
rect 388119 662766 393657 664360
rect 388119 661297 389052 662766
rect 388119 661263 388163 661297
rect 388197 661263 388235 661297
rect 388269 661263 388307 661297
rect 388341 661263 388379 661297
rect 388413 661263 388451 661297
rect 388485 661263 388523 661297
rect 388557 661263 388595 661297
rect 388629 661263 388667 661297
rect 388701 661263 388739 661297
rect 388773 661263 388811 661297
rect 388845 661263 388883 661297
rect 388917 661263 388955 661297
rect 388989 661263 389052 661297
rect 388119 661245 389052 661263
rect 380201 660801 387356 660899
rect 380201 660767 387303 660801
rect 387337 660767 387356 660801
rect 380201 660729 387356 660767
rect 380201 660695 387303 660729
rect 387337 660695 387356 660729
rect 380201 660657 387356 660695
rect 380201 660623 387303 660657
rect 387337 660623 387356 660657
rect 380201 660585 387356 660623
rect 380201 660551 387303 660585
rect 387337 660551 387356 660585
rect 380201 660513 387356 660551
rect 380201 660479 387303 660513
rect 387337 660479 387356 660513
rect 380201 660441 387356 660479
rect 380201 660407 387303 660441
rect 387337 660407 387356 660441
rect 380201 660369 387356 660407
rect 380201 660335 387303 660369
rect 387337 660335 387356 660369
rect 380201 660297 387356 660335
rect 380201 660263 387303 660297
rect 387337 660263 387356 660297
rect 380201 660225 387356 660263
rect 380201 660191 387303 660225
rect 387337 660191 387356 660225
rect 380201 660153 387356 660191
rect 380201 660119 387303 660153
rect 387337 660119 387356 660153
rect 380201 660081 387356 660119
rect 380201 660047 387303 660081
rect 387337 660047 387356 660081
rect 380201 660009 387356 660047
rect 380201 659975 387303 660009
rect 387337 659975 387356 660009
rect 380201 659937 387356 659975
rect 380201 659903 387303 659937
rect 387337 659903 387356 659937
rect 380201 659865 387356 659903
rect 380201 659831 387303 659865
rect 387337 659831 387356 659865
rect 380201 659793 387356 659831
rect 380201 659759 387303 659793
rect 387337 659759 387356 659793
rect 387970 660742 389065 660764
rect 387970 659794 387979 660742
rect 389055 659794 389065 660742
rect 387970 659773 389065 659794
rect 380201 659721 387356 659759
rect 380201 659687 387303 659721
rect 387337 659687 387356 659721
rect 380201 659649 387356 659687
rect 380201 659615 387303 659649
rect 387337 659615 387356 659649
rect 380201 659577 387356 659615
rect 380201 659543 387303 659577
rect 387337 659543 387356 659577
rect 380201 659505 387356 659543
rect 380201 659471 387303 659505
rect 387337 659471 387356 659505
rect 380201 659433 387356 659471
rect 380201 659399 387303 659433
rect 387337 659399 387356 659433
rect 380201 659361 387356 659399
rect 380201 659327 387303 659361
rect 387337 659327 387356 659361
rect 380201 659289 387356 659327
rect 380201 659255 387303 659289
rect 387337 659255 387356 659289
rect 380201 659217 387356 659255
rect 380201 659183 387303 659217
rect 387337 659183 387356 659217
rect 380201 659141 387356 659183
rect 381359 651521 383362 659141
rect 392017 652046 393657 662766
rect 466927 661182 467917 671001
rect 513525 668328 515211 668609
rect 513525 666548 513698 668328
rect 515030 666548 515211 668328
rect 508085 665566 513201 665624
rect 508085 665532 513146 665566
rect 513180 665532 513201 665566
rect 508085 665494 513201 665532
rect 508085 665460 513146 665494
rect 513180 665460 513201 665494
rect 508085 665422 513201 665460
rect 508085 665388 513146 665422
rect 513180 665388 513201 665422
rect 508085 665350 513201 665388
rect 508085 665316 513146 665350
rect 513180 665316 513201 665350
rect 508085 665278 513201 665316
rect 508085 665244 513146 665278
rect 513180 665244 513201 665278
rect 508085 665206 513201 665244
rect 508085 665172 513146 665206
rect 513180 665172 513201 665206
rect 508085 665134 513201 665172
rect 508085 665100 513146 665134
rect 513180 665100 513201 665134
rect 508085 665062 513201 665100
rect 508085 665028 513146 665062
rect 513180 665028 513201 665062
rect 508085 664990 513201 665028
rect 508085 664956 513146 664990
rect 513180 664956 513201 664990
rect 508085 664918 513201 664956
rect 508085 664884 513146 664918
rect 513180 664884 513201 664918
rect 508085 664846 513201 664884
rect 508085 664812 513146 664846
rect 513180 664812 513201 664846
rect 508085 664774 513201 664812
rect 508085 664740 513146 664774
rect 513180 664740 513201 664774
rect 508085 664702 513201 664740
rect 508085 664668 513146 664702
rect 513180 664668 513201 664702
rect 508085 664630 513201 664668
rect 508085 664596 513146 664630
rect 513180 664596 513201 664630
rect 508085 664558 513201 664596
rect 508085 664524 513146 664558
rect 513180 664524 513201 664558
rect 508085 664486 513201 664524
rect 508085 664452 513146 664486
rect 513180 664452 513201 664486
rect 508085 664414 513201 664452
rect 508085 664380 513146 664414
rect 513180 664380 513201 664414
rect 508085 664342 513201 664380
rect 508085 664308 513146 664342
rect 513180 664308 513201 664342
rect 508085 664270 513201 664308
rect 508085 664236 513146 664270
rect 513180 664236 513201 664270
rect 508085 664198 513201 664236
rect 508085 664164 513146 664198
rect 513180 664164 513201 664198
rect 508085 664126 513201 664164
rect 508085 664092 513146 664126
rect 513180 664092 513201 664126
rect 508085 664054 513201 664092
rect 508085 664020 513146 664054
rect 513180 664020 513201 664054
rect 508085 663982 513201 664020
rect 508085 663948 513146 663982
rect 513180 663948 513201 663982
rect 508085 663910 513201 663948
rect 508085 663876 513146 663910
rect 513180 663876 513201 663910
rect 508085 663838 513201 663876
rect 508085 663804 513146 663838
rect 513180 663804 513201 663838
rect 508085 663766 513201 663804
rect 508085 663732 513146 663766
rect 513180 663732 513201 663766
rect 508085 663694 513201 663732
rect 508085 663660 513146 663694
rect 513180 663660 513201 663694
rect 508085 663622 513201 663660
rect 513525 663623 515211 666548
rect 515582 664904 525173 664959
rect 515582 664870 515592 664904
rect 515626 664902 525173 664904
rect 515626 664870 525120 664902
rect 515582 664868 525120 664870
rect 525154 664868 525173 664902
rect 515582 664832 525173 664868
rect 515582 664798 515592 664832
rect 515626 664830 525173 664832
rect 515626 664798 525120 664830
rect 515582 664796 525120 664798
rect 525154 664796 525173 664830
rect 515582 664760 525173 664796
rect 515582 664726 515592 664760
rect 515626 664758 525173 664760
rect 515626 664726 525120 664758
rect 515582 664724 525120 664726
rect 525154 664724 525173 664758
rect 515582 664688 525173 664724
rect 515582 664654 515592 664688
rect 515626 664686 525173 664688
rect 515626 664654 525120 664686
rect 515582 664652 525120 664654
rect 525154 664652 525173 664686
rect 515582 664616 525173 664652
rect 515582 664582 515592 664616
rect 515626 664614 525173 664616
rect 515626 664582 525120 664614
rect 515582 664580 525120 664582
rect 525154 664580 525173 664614
rect 515582 664544 525173 664580
rect 515582 664510 515592 664544
rect 515626 664542 525173 664544
rect 515626 664510 525120 664542
rect 515582 664508 525120 664510
rect 525154 664508 525173 664542
rect 515582 664472 525173 664508
rect 515582 664438 515592 664472
rect 515626 664470 525173 664472
rect 515626 664438 525120 664470
rect 515582 664436 525120 664438
rect 525154 664436 525173 664470
rect 515582 664400 525173 664436
rect 515582 664366 515592 664400
rect 515626 664398 525173 664400
rect 515626 664366 525120 664398
rect 515582 664364 525120 664366
rect 525154 664364 525173 664398
rect 515582 664328 525173 664364
rect 515582 664294 515592 664328
rect 515626 664326 525173 664328
rect 515626 664294 525120 664326
rect 515582 664292 525120 664294
rect 525154 664292 525173 664326
rect 515582 664256 525173 664292
rect 515582 664222 515592 664256
rect 515626 664254 525173 664256
rect 515626 664222 525120 664254
rect 515582 664220 525120 664222
rect 525154 664220 525173 664254
rect 515582 664184 525173 664220
rect 515582 664150 515592 664184
rect 515626 664182 525173 664184
rect 515626 664150 525120 664182
rect 515582 664148 525120 664150
rect 525154 664148 525173 664182
rect 515582 664112 525173 664148
rect 515582 664078 515592 664112
rect 515626 664110 525173 664112
rect 515626 664078 525120 664110
rect 515582 664076 525120 664078
rect 525154 664076 525173 664110
rect 515582 664040 525173 664076
rect 515582 664006 515592 664040
rect 515626 664038 525173 664040
rect 515626 664006 525120 664038
rect 515582 664004 525120 664006
rect 525154 664004 525173 664038
rect 515582 663968 525173 664004
rect 515582 663934 515592 663968
rect 515626 663966 525173 663968
rect 515626 663934 525120 663966
rect 515582 663932 525120 663934
rect 525154 663932 525173 663966
rect 515582 663896 525173 663932
rect 515582 663862 515592 663896
rect 515626 663894 525173 663896
rect 515626 663862 525120 663894
rect 515582 663860 525120 663862
rect 525154 663860 525173 663894
rect 515582 663801 525173 663860
rect 508085 663588 513146 663622
rect 513180 663588 513201 663622
rect 508085 663548 513201 663588
rect 513819 663533 514874 663551
rect 513819 663499 513861 663533
rect 513895 663499 513933 663533
rect 513967 663499 514005 663533
rect 514039 663499 514077 663533
rect 514111 663499 514149 663533
rect 514183 663499 514221 663533
rect 514255 663499 514293 663533
rect 514327 663499 514365 663533
rect 514399 663499 514437 663533
rect 514471 663499 514509 663533
rect 514543 663499 514581 663533
rect 514615 663499 514653 663533
rect 514687 663499 514725 663533
rect 514759 663499 514797 663533
rect 514831 663499 514874 663533
rect 525436 663513 534530 664820
rect 513819 660979 514874 663499
rect 525540 663115 526832 663133
rect 525540 663081 525588 663115
rect 525622 663081 525660 663115
rect 525694 663081 525732 663115
rect 525766 663081 525804 663115
rect 525838 663081 525876 663115
rect 525910 663081 525948 663115
rect 525982 663081 526020 663115
rect 526054 663081 526092 663115
rect 526126 663081 526164 663115
rect 526198 663081 526236 663115
rect 526270 663081 526308 663115
rect 526342 663081 526380 663115
rect 526414 663081 526452 663115
rect 526486 663081 526524 663115
rect 526558 663081 526596 663115
rect 526630 663081 526668 663115
rect 526702 663081 526740 663115
rect 526774 663081 526832 663115
rect 525540 662290 526832 663081
rect 466886 660600 467985 660626
rect 466886 659524 466897 660600
rect 467973 659524 467985 660600
rect 513819 660543 514002 660979
rect 514694 660543 514874 660979
rect 513819 660426 514874 660543
rect 519417 660880 526832 662290
rect 519417 660444 519721 660880
rect 520797 660444 526832 660880
rect 468606 660203 479200 660244
rect 519417 660237 526832 660444
rect 468606 660169 468615 660203
rect 468649 660169 479200 660203
rect 468606 660131 479200 660169
rect 468606 660097 468615 660131
rect 468649 660097 479200 660131
rect 468606 660059 479200 660097
rect 468606 660025 468615 660059
rect 468649 660025 479200 660059
rect 468606 659987 479200 660025
rect 468606 659953 468615 659987
rect 468649 659953 479200 659987
rect 468606 659915 479200 659953
rect 468606 659881 468615 659915
rect 468649 659881 479200 659915
rect 468606 659843 479200 659881
rect 468606 659809 468615 659843
rect 468649 659809 479200 659843
rect 468606 659771 479200 659809
rect 468606 659737 468615 659771
rect 468649 659737 479200 659771
rect 468606 659699 479200 659737
rect 468606 659665 468615 659699
rect 468649 659665 479200 659699
rect 468606 659623 479200 659665
rect 466886 659498 467985 659524
rect 496613 654614 497583 654641
rect 496613 653794 496624 654614
rect 497572 653794 497583 654614
rect 496613 653767 497583 653794
rect 497794 654106 502667 654162
rect 497794 654072 497802 654106
rect 497836 654094 502667 654106
rect 497836 654072 502430 654094
rect 497794 654034 502430 654072
rect 497794 654000 497802 654034
rect 497836 654000 502430 654034
rect 497794 653962 502430 654000
rect 497794 653928 497802 653962
rect 497836 653928 502430 653962
rect 497794 653890 502430 653928
rect 497794 653856 497802 653890
rect 497836 653856 502430 653890
rect 497794 653818 502430 653856
rect 497794 653784 497802 653818
rect 497836 653784 502430 653818
rect 497794 653746 502430 653784
rect 497794 653712 497802 653746
rect 497836 653712 502430 653746
rect 497794 653674 502430 653712
rect 497794 653640 497802 653674
rect 497836 653658 502430 653674
rect 502610 653658 502667 654094
rect 497836 653640 502667 653658
rect 497794 653601 502667 653640
rect 392017 652012 392059 652046
rect 392093 652012 392131 652046
rect 392165 652012 392203 652046
rect 392237 652012 392275 652046
rect 392309 652012 392347 652046
rect 392381 652012 392419 652046
rect 392453 652012 392491 652046
rect 392525 652012 392563 652046
rect 392597 652012 392635 652046
rect 392669 652012 392707 652046
rect 392741 652012 392779 652046
rect 392813 652012 392851 652046
rect 392885 652012 392923 652046
rect 392957 652012 392995 652046
rect 393029 652012 393067 652046
rect 393101 652012 393139 652046
rect 393173 652012 393211 652046
rect 393245 652012 393283 652046
rect 393317 652012 393355 652046
rect 393389 652012 393427 652046
rect 393461 652012 393499 652046
rect 393533 652012 393571 652046
rect 393605 652012 393657 652046
rect 392017 652006 393657 652012
rect 496862 653416 497517 653435
rect 496862 653382 496907 653416
rect 496941 653382 496979 653416
rect 497013 653382 497051 653416
rect 497085 653382 497123 653416
rect 497157 653382 497195 653416
rect 497229 653382 497267 653416
rect 497301 653382 497339 653416
rect 497373 653382 497411 653416
rect 497445 653382 497517 653416
rect 496862 652278 497517 653382
rect 391993 651847 393755 651866
rect 381359 651451 391700 651521
rect 381359 651417 391648 651451
rect 391682 651417 391700 651451
rect 381359 651379 391700 651417
rect 381359 651345 391648 651379
rect 391682 651345 391700 651379
rect 381359 651307 391700 651345
rect 381359 651273 391648 651307
rect 391682 651273 391700 651307
rect 381359 651235 391700 651273
rect 381359 651201 391648 651235
rect 391682 651201 391700 651235
rect 381359 651163 391700 651201
rect 381359 651129 391648 651163
rect 391682 651129 391700 651163
rect 381359 651091 391700 651129
rect 381359 651057 391648 651091
rect 391682 651057 391700 651091
rect 381359 651019 391700 651057
rect 381359 650985 391648 651019
rect 391682 650985 391700 651019
rect 381359 650947 391700 650985
rect 381359 650913 391648 650947
rect 391682 650913 391700 650947
rect 381359 650875 391700 650913
rect 381359 650841 391648 650875
rect 391682 650841 391700 650875
rect 381359 650803 391700 650841
rect 381359 650769 391648 650803
rect 391682 650769 391700 650803
rect 381359 650731 391700 650769
rect 381359 650697 391648 650731
rect 391682 650697 391700 650731
rect 381359 650659 391700 650697
rect 381359 650625 391648 650659
rect 391682 650625 391700 650659
rect 381359 650587 391700 650625
rect 381359 650553 391648 650587
rect 391682 650553 391700 650587
rect 381359 650515 391700 650553
rect 381359 650481 391648 650515
rect 391682 650481 391700 650515
rect 381359 650443 391700 650481
rect 381359 650409 391648 650443
rect 391682 650409 391700 650443
rect 381359 650371 391700 650409
rect 381359 650337 391648 650371
rect 391682 650337 391700 650371
rect 381359 650299 391700 650337
rect 381359 650265 391648 650299
rect 391682 650265 391700 650299
rect 381359 650198 391700 650265
rect 391993 650131 392016 651847
rect 393732 650131 393755 651847
rect 496862 651074 496976 652278
rect 497412 651074 497517 652278
rect 496862 650872 497517 651074
rect 391993 650112 393755 650131
<< via1 >>
rect 386813 692241 388529 693765
rect 386992 690647 387684 691147
rect 501840 685846 503428 687114
rect 501807 684657 502051 685157
rect 494238 680582 494994 680954
rect 467069 671109 467761 672377
rect 388233 666413 388925 667233
rect 387979 659794 389055 660742
rect 513698 666548 515030 668328
rect 466897 659524 467973 660600
rect 514002 660543 514694 660979
rect 519721 660444 520797 660880
rect 496624 653794 497572 654614
rect 502430 653658 502610 654094
rect 392016 650131 393732 651847
rect 496976 651074 497412 652278
<< metal2 >>
rect 499716 699818 525351 700436
rect 499716 696802 511635 699818
rect 514331 696802 521640 699818
rect 524336 696802 525351 699818
rect 499716 696313 525351 696802
rect 386691 693791 388631 693948
rect 386691 693765 386843 693791
rect 388499 693765 388631 693791
rect 386691 692241 386813 693765
rect 388529 692241 388631 693765
rect 386691 692215 386843 692241
rect 388499 692215 388631 692241
rect 386691 692048 388631 692215
rect 386877 691147 388253 691211
rect 386877 690647 386992 691147
rect 387684 690647 388253 691147
rect 386877 680424 388253 690647
rect 499716 687967 509125 696313
rect 501651 687114 503642 687376
rect 501651 685846 501840 687114
rect 503428 685846 503642 687114
rect 501651 685666 503642 685846
rect 494066 685157 502135 685259
rect 494066 684657 501807 685157
rect 502051 684657 502135 685157
rect 494066 684550 502135 684657
rect 494073 680954 495148 684550
rect 494073 680582 494238 680954
rect 494994 680582 495148 680954
rect 386877 679955 390668 680424
rect 386877 673553 387252 679955
rect 386899 671979 387252 673553
rect 390268 671979 390668 679955
rect 494073 679350 495148 680582
rect 386899 671303 390668 671979
rect 466924 672377 467910 672501
rect 466924 672371 467069 672377
rect 467761 672371 467910 672377
rect 387674 667233 389918 671303
rect 466924 671115 467067 672371
rect 467763 671115 467910 672371
rect 466924 671109 467069 671115
rect 467761 671109 467910 671115
rect 466924 671001 467910 671109
rect 387674 666413 388233 667233
rect 388925 666413 389918 667233
rect 387674 666033 389918 666413
rect 513525 668346 515211 668609
rect 513525 668328 513736 668346
rect 514992 668328 515211 668346
rect 513525 666548 513698 668328
rect 515030 666548 515211 668328
rect 513525 666530 513736 666548
rect 514992 666530 515211 666548
rect 513525 666352 515211 666530
rect 511501 660979 521142 661097
rect 387852 660742 389235 660906
rect 387852 659794 387979 660742
rect 389055 659794 389235 660742
rect 387852 659617 389235 659794
rect 466656 660610 468179 660817
rect 466656 659514 466887 660610
rect 467983 659514 468179 660610
rect 466656 659349 468179 659514
rect 511501 660543 514002 660979
rect 514694 660880 521142 660979
rect 514694 660543 519721 660880
rect 511501 660444 519721 660543
rect 520797 660444 521142 660880
rect 496545 654632 497667 654747
rect 496545 654614 496630 654632
rect 497566 654614 497667 654632
rect 496545 653794 496624 654614
rect 497572 653794 497667 654614
rect 511501 654506 521142 660444
rect 502950 654165 521142 654506
rect 496545 653776 496630 653794
rect 497566 653776 497667 653794
rect 496545 653687 497667 653776
rect 502371 654094 521142 654165
rect 502371 653658 502430 654094
rect 502610 653658 521142 654094
rect 502371 653601 521142 653658
rect 502950 653172 521142 653601
rect 496951 652278 497438 652305
rect 391947 651857 393810 651920
rect 391947 650121 392006 651857
rect 393742 650121 393810 651857
rect 496951 651074 496976 652278
rect 497412 651074 497438 652278
rect 496951 651048 497438 651074
rect 391947 649956 393810 650121
rect 511501 633907 521142 653172
rect 511501 628331 513582 633907
rect 520038 628331 521142 633907
rect 511501 626986 521142 628331
rect 5352 553952 9224 554786
rect 5352 549736 5828 553952
rect 8524 549736 9224 553952
rect 5352 528326 9224 549736
rect 5262 524863 190898 528326
rect 5262 518087 178927 524863
rect 187223 518087 190898 524863
rect 5262 516760 190898 518087
rect 175366 385504 176982 385578
rect 1202 385018 176982 385504
rect 1202 381762 1994 385018
rect 4130 381762 176982 385018
rect 1202 381490 176982 381762
rect 175366 337344 176982 381490
rect 174138 337300 176982 337344
rect 173622 336670 176982 337300
rect 173622 336644 175730 336670
rect 174138 336640 175730 336644
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 511635 696802 514331 699818
rect 521640 696802 524336 699818
rect 386843 693765 388499 693791
rect 386843 692241 388499 693765
rect 386843 692215 388499 692241
rect 501846 685852 503422 687108
rect 387252 671979 390268 679955
rect 467067 671115 467069 672371
rect 467069 671115 467761 672371
rect 467761 671115 467763 672371
rect 513736 668328 514992 668346
rect 513736 666548 514992 668328
rect 513736 666530 514992 666548
rect 388009 659800 389025 660736
rect 466887 660600 467983 660610
rect 466887 659524 466897 660600
rect 466897 659524 467973 660600
rect 467973 659524 467983 660600
rect 466887 659514 467983 659524
rect 496630 654614 497566 654632
rect 496630 653794 497566 654614
rect 496630 653776 497566 653794
rect 392006 651847 393742 651857
rect 392006 650131 392016 651847
rect 392016 650131 393732 651847
rect 393732 650131 393742 651847
rect 392006 650121 393742 650131
rect 513582 628331 520038 633907
rect 5828 549736 8524 553952
rect 178927 518087 187223 524863
rect 1994 381762 4130 385018
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 16194 702283 21448 702300
rect 16028 694401 21448 702283
rect 68194 702217 73846 702300
rect 120194 702298 125382 702300
rect 165594 702298 170580 702300
rect 16028 691457 16476 694401
rect 20940 691457 21448 694401
rect 16028 691092 21448 691457
rect 1709 685242 59742 685252
rect 0 684489 59742 685242
rect 0 681065 54399 684489
rect 59343 681065 59742 684489
rect 0 680368 59742 681065
rect 0 680242 1700 680368
rect 67682 658160 73846 702217
rect 120078 689243 125382 702298
rect 67760 656983 73846 658160
rect 67760 654359 68696 656983
rect 72920 654359 73846 656983
rect 67760 653506 73846 654359
rect 0 643842 1660 648642
rect 116940 640785 127975 689243
rect 0 633842 1660 638642
rect 116940 633921 119075 640785
rect 126259 633921 127975 640785
rect 116940 632804 127975 633921
rect 165284 621462 170580 702298
rect 14132 612258 170822 621462
rect 0 562844 1660 564242
rect 0 562025 4628 562844
rect 0 559442 1660 562025
rect 2853 554860 4603 562025
rect 2853 554242 9298 554860
rect 0 553952 9298 554242
rect 0 549736 5828 553952
rect 8524 549736 9298 553952
rect 14602 553900 25988 612258
rect 165284 612044 170580 612258
rect 217648 603536 221632 702300
rect 318942 632280 323910 702300
rect 413394 702299 418405 702300
rect 465394 702299 470394 704800
rect 413374 701955 418405 702299
rect 413374 700451 414079 701955
rect 417743 700451 418405 701955
rect 413374 700212 418405 700451
rect 465303 701799 470414 702299
rect 465303 695495 466102 701799
rect 469766 695495 470414 701799
rect 510594 699818 515394 704800
rect 510594 696802 511635 699818
rect 514331 696802 515394 699818
rect 510594 696313 515394 696802
rect 520594 699818 525394 704800
rect 566594 702300 571594 704800
rect 566594 702296 571462 702300
rect 520594 696802 521640 699818
rect 524336 696802 525394 699818
rect 520594 696313 525394 696802
rect 465303 694826 470414 695495
rect 472532 694612 496804 694656
rect 405424 694323 496804 694612
rect 405424 694010 495102 694323
rect 386691 693795 388631 693948
rect 386691 692211 386839 693795
rect 388503 692211 388631 693795
rect 386691 692048 388631 692211
rect 405424 691626 406211 694010
rect 411635 691699 495102 694010
rect 496446 691699 496804 694323
rect 411635 691626 496804 691699
rect 405424 691458 496804 691626
rect 405424 691262 478494 691458
rect 501651 687112 503642 687376
rect 501651 685848 501842 687112
rect 503426 685848 503642 687112
rect 501651 685666 503642 685848
rect 386899 679959 390668 680424
rect 386899 671975 387248 679959
rect 390272 671975 390668 679959
rect 386899 671303 390668 671975
rect 440756 679130 472683 680412
rect 440756 672666 443027 679130
rect 452611 672666 472683 679130
rect 440756 672371 472683 672666
rect 440756 671115 467067 672371
rect 467763 671388 472683 672371
rect 509653 674517 518248 674844
rect 509653 672053 515807 674517
rect 517951 672053 518248 674517
rect 509653 671772 518248 672053
rect 509653 671771 518242 671772
rect 467763 671115 479676 671388
rect 440756 670996 479676 671115
rect 387852 660740 389235 660906
rect 387852 659796 388005 660740
rect 389029 659796 389235 660740
rect 387852 659617 389235 659796
rect 391947 651861 393810 651920
rect 391947 650117 392002 651861
rect 393746 650117 393810 651861
rect 391947 649956 393810 650117
rect 440756 634756 454681 670996
rect 460702 667842 464759 668464
rect 468400 668314 479676 670996
rect 566522 670616 571462 702296
rect 574676 682984 582300 682991
rect 574676 682293 584800 682984
rect 574676 678469 575284 682293
rect 577988 678469 584800 682293
rect 574676 677984 584800 678469
rect 574676 677978 582300 677984
rect 510812 669564 571462 670616
rect 468400 668264 476816 668314
rect 468400 668240 472648 668264
rect 478486 668084 479676 668314
rect 503876 668346 534529 668575
rect 460702 663138 461606 667842
rect 464230 666065 464759 667842
rect 471704 666710 481406 666878
rect 471704 666406 472068 666710
rect 476212 666406 481406 666710
rect 471704 666258 481406 666406
rect 503876 666530 513736 668346
rect 514992 668160 534529 668346
rect 514992 666816 531160 668160
rect 533864 666816 534529 668160
rect 514992 666530 534529 666816
rect 503876 666352 534529 666530
rect 464230 664995 479143 666065
rect 464230 663138 464759 664995
rect 460702 662421 464759 663138
rect 466656 660614 468179 660817
rect 466656 660610 466923 660614
rect 467947 660610 468179 660614
rect 466656 659514 466887 660610
rect 467983 659514 468179 660610
rect 466656 659510 466923 659514
rect 467947 659510 468179 659514
rect 466656 659349 468179 659510
rect 510461 659393 519321 659775
rect 510461 656689 515436 659393
rect 518940 656689 519321 659393
rect 510461 656346 519321 656689
rect 496545 654636 497667 654747
rect 496545 653772 496626 654636
rect 497570 653772 497667 654636
rect 496545 653687 497667 653772
rect 573550 644584 582340 644618
rect 573550 639784 584800 644584
rect 573550 634756 582340 639784
rect 440756 634584 582340 634756
rect 440756 633907 584800 634584
rect 318942 629780 323636 632280
rect 317558 629626 323636 629780
rect 245352 626867 323636 629626
rect 440756 628331 513582 633907
rect 520038 629784 584800 633907
rect 520038 628331 582027 629784
rect 440756 626915 582027 628331
rect 245352 624706 246463 626867
rect 244934 619683 246463 624706
rect 252767 619683 323636 626867
rect 244934 618958 323636 619683
rect 217648 596032 218304 603536
rect 221088 596032 221632 603536
rect 217648 595400 221632 596032
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 580997 584182 583475 584190
rect 515013 583674 583475 584182
rect 515013 583562 584800 583674
rect 515013 583499 583475 583562
rect 515013 575115 515430 583499
rect 518774 583163 583475 583499
rect 518774 575115 581000 583163
rect 515013 574808 581000 575115
rect 582420 555362 584274 555374
rect 0 549498 9298 549736
rect 14408 553184 25988 553900
rect 0 549442 1668 549498
rect 14408 549474 25928 553184
rect 582340 550562 584800 555362
rect 14408 549076 25988 549474
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 1292 385018 4602 385526
rect 1292 383512 1994 385018
rect 910 381976 1994 383512
rect -800 381864 1994 381976
rect 910 381762 1994 381864
rect 4130 381762 4602 385018
rect 910 381546 4602 381762
rect 910 381491 2080 381546
rect 1065 381490 2080 381491
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 14602 234506 25988 549076
rect 582340 540562 584800 545362
rect 177162 524863 188990 526546
rect 177162 518087 178927 524863
rect 187223 518087 188990 524863
rect 177162 423452 188990 518087
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 530221 496519 580953 497230
rect 530221 493015 530852 496519
rect 533956 494540 580953 496519
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 533956 494252 583330 494540
rect 533956 494140 584800 494252
rect 533956 493663 583330 494140
rect 533956 493015 580953 493663
rect 530221 492473 580953 493015
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 16476 691457 20940 694401
rect 54399 681065 59343 684489
rect 68696 654359 72920 656983
rect 119075 633921 126259 640785
rect 414079 700451 417743 701955
rect 466102 695495 469766 701799
rect 386839 693791 388503 693795
rect 386839 692215 386843 693791
rect 386843 692215 388499 693791
rect 388499 692215 388503 693791
rect 386839 692211 388503 692215
rect 406211 691626 411635 694010
rect 495102 691699 496446 694323
rect 501842 687108 503426 687112
rect 501842 685852 501846 687108
rect 501846 685852 503422 687108
rect 503422 685852 503426 687108
rect 501842 685848 503426 685852
rect 387248 679955 390272 679959
rect 387248 671979 387252 679955
rect 387252 671979 390268 679955
rect 390268 671979 390272 679955
rect 387248 671975 390272 671979
rect 443027 672666 452611 679130
rect 515807 672053 517951 674517
rect 388005 660736 389029 660740
rect 388005 659800 388009 660736
rect 388009 659800 389025 660736
rect 389025 659800 389029 660736
rect 388005 659796 389029 659800
rect 392002 651857 393746 651861
rect 392002 650121 392006 651857
rect 392006 650121 393742 651857
rect 393742 650121 393746 651857
rect 392002 650117 393746 650121
rect 575284 678469 577988 682293
rect 461606 663138 464230 667842
rect 472068 666406 476212 666710
rect 531160 666816 533864 668160
rect 466923 660610 467947 660614
rect 466923 659514 467947 660610
rect 466923 659510 467947 659514
rect 515436 656689 518940 659393
rect 496626 654632 497570 654636
rect 496626 653776 496630 654632
rect 496630 653776 497566 654632
rect 497566 653776 497570 654632
rect 496626 653772 497570 653776
rect 246463 619683 252767 626867
rect 218304 596032 221088 603536
rect 515430 575115 518774 583499
rect 530852 493015 533956 496519
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 465394 702299 470394 702300
rect 413368 701961 418404 702299
rect 413368 701955 414193 701961
rect 417629 701955 418404 701961
rect 413368 700451 414079 701955
rect 417743 700451 418404 701955
rect 413368 700445 414193 700451
rect 417629 700445 418404 700451
rect 413368 700215 418404 700445
rect 465303 701799 486932 702299
rect 465303 695495 466102 701799
rect 469766 695495 486932 701799
rect 397560 695124 412594 695352
rect 15908 694401 412594 695124
rect 465303 694840 486932 695495
rect 465303 694826 470414 694840
rect 15908 691457 16476 694401
rect 20940 694010 412594 694401
rect 20940 693795 406211 694010
rect 20940 692211 386839 693795
rect 388503 692211 406211 693795
rect 20940 691626 406211 692211
rect 411635 691626 412594 694010
rect 20940 691457 412594 691626
rect 15908 690804 412594 691457
rect 397560 690628 412594 690804
rect 53538 684489 59808 685318
rect 53538 681065 54399 684489
rect 59343 681065 59808 684489
rect 53538 648101 59808 681065
rect 81882 679959 455140 680411
rect 81882 671975 387248 679959
rect 390272 679130 455140 679959
rect 483624 679283 486932 694840
rect 494816 694323 496732 694654
rect 494816 693530 495102 694323
rect 494804 691699 495102 693530
rect 496446 691699 496732 694323
rect 494804 691490 496732 691699
rect 494804 687554 496680 691490
rect 494834 687378 496680 687554
rect 494834 687262 504530 687378
rect 494834 687112 504560 687262
rect 494834 685848 501842 687112
rect 503426 685848 504560 687112
rect 494834 685474 504560 685848
rect 494834 685386 504530 685474
rect 494834 685356 496680 685386
rect 574676 682293 578731 682938
rect 390272 672666 443027 679130
rect 452611 672666 455140 679130
rect 574676 678469 575284 682293
rect 577988 678469 578731 682293
rect 574676 677978 578731 678469
rect 390272 671975 455140 672666
rect 81882 671370 455140 671975
rect 515442 674523 518248 674844
rect 515442 672047 515801 674523
rect 517957 672047 518248 674523
rect 515442 671772 518248 672047
rect 460702 667848 464759 668464
rect 460702 667842 461680 667848
rect 464156 667842 464759 667848
rect 460702 663138 461606 667842
rect 464230 663138 464759 667842
rect 530221 668160 534529 668575
rect 460702 663132 461680 663138
rect 464156 663132 464759 663138
rect 460702 662421 464759 663132
rect 471786 666710 476352 666868
rect 471786 666406 472068 666710
rect 476212 666406 476352 666710
rect 387851 660740 389235 660906
rect 387851 659796 388005 660740
rect 389029 659796 389235 660740
rect 387851 657590 389235 659796
rect 466656 660614 468174 660820
rect 466656 659510 466923 660614
rect 467947 659510 468174 660614
rect 466656 657728 468174 659510
rect 471786 657728 476352 666406
rect 530221 666816 531160 668160
rect 533864 666816 534529 668160
rect 466286 657590 476352 657728
rect 67760 656983 476352 657590
rect 67760 654359 68696 656983
rect 72920 655060 476352 656983
rect 515013 659393 519321 659775
rect 515013 656689 515436 659393
rect 518940 656689 519321 659393
rect 72920 654359 476406 655060
rect 67760 652424 476406 654359
rect 494784 654636 497667 654747
rect 494784 653772 496626 654636
rect 497570 653772 497667 654636
rect 494784 653686 497667 653772
rect 391947 651861 393810 651920
rect 391947 650117 392002 651861
rect 393746 650117 393810 651861
rect 391947 649956 393810 650117
rect 497501 650170 501446 650191
rect 491326 650042 496078 650084
rect 490858 648740 496078 650042
rect 53538 644985 54348 648101
rect 59064 644985 59808 648101
rect 53538 644332 59808 644985
rect 490670 648726 496078 648740
rect 490670 647975 493914 648726
rect 490670 644859 491042 647975
rect 493198 645560 493914 647975
rect 497501 645560 501468 650170
rect 493198 644859 493868 645560
rect 490670 644432 493868 644859
rect 116934 640785 127975 642210
rect 116934 633921 119075 640785
rect 126259 633921 127975 640785
rect 116934 632792 127975 633921
rect 497501 641619 501446 645560
rect 497501 638503 497693 641619
rect 501129 638503 501446 641619
rect 497501 637430 501446 638503
rect 497501 633994 497971 637430
rect 500767 633994 501446 637430
rect 497501 632828 501446 633994
rect 245344 626867 253976 627902
rect 245344 619683 246463 626867
rect 252767 619683 253976 626867
rect 84806 604254 208762 604378
rect 84806 604132 221660 604254
rect 63698 603536 221660 604132
rect 63698 596032 218304 603536
rect 221088 596032 221660 603536
rect 63698 595214 221660 596032
rect 63698 595050 208762 595214
rect 63698 554306 74252 595050
rect 245344 428990 253976 619683
rect 515013 583499 519321 656689
rect 515013 575115 515430 583499
rect 518774 575115 519321 583499
rect 515013 574609 519321 575115
rect 530221 496519 534529 666816
rect 530221 493015 530852 496519
rect 533956 493015 534529 496519
rect 530221 492473 534529 493015
<< via4 >>
rect 414193 701955 417629 701961
rect 414193 700451 417629 701955
rect 414193 700445 417629 700451
rect 575398 678503 577874 682259
rect 515801 674517 517957 674523
rect 515801 672053 515807 674517
rect 515807 672053 517951 674517
rect 517951 672053 517957 674517
rect 515801 672047 517957 672053
rect 461680 667842 464156 667848
rect 461680 663138 464156 667842
rect 461680 663132 464156 663138
rect 392116 650231 393632 651747
rect 54348 644985 59064 648101
rect 491042 644859 493198 647975
rect 119189 634035 126145 640671
rect 497693 638503 501129 641619
rect 497971 633994 500767 637430
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 167655 700990 169333 702300
rect 177453 700990 179131 702300
rect 219319 701674 220665 702300
rect 229375 701674 230398 702300
rect 167655 700532 179165 700990
rect 219319 700638 230411 701674
rect 320552 700638 322040 702300
rect 331030 700638 332518 702300
rect 413394 701961 418396 702299
rect 167666 700204 179165 700532
rect 320433 698996 332746 700638
rect 413394 700445 414193 701961
rect 417629 700445 418396 701961
rect 413394 668441 418396 700445
rect 515442 682259 578716 682935
rect 515442 678503 575398 682259
rect 577874 678503 578716 682259
rect 515442 674523 578716 678503
rect 515442 672047 515801 674523
rect 517957 672047 578716 674523
rect 515442 671771 578716 672047
rect 413394 667848 464766 668441
rect 413394 663132 461680 667848
rect 464156 663132 464766 667848
rect 413394 662413 464766 663132
rect 391947 651747 393810 651920
rect 391947 650231 392116 651747
rect 393632 650231 393810 651747
rect 391947 648544 393810 650231
rect 53770 648101 493804 648544
rect 53770 644985 54348 648101
rect 59064 647975 493804 648101
rect 59064 644985 491042 647975
rect 53770 644859 491042 644985
rect 493198 644859 493804 647975
rect 53770 644498 493804 644859
rect 116940 641619 501378 642210
rect 116940 640671 497693 641619
rect 116940 634035 119189 640671
rect 126145 638503 497693 640671
rect 501129 638503 501378 641619
rect 126145 637430 501378 638503
rect 126145 634035 497971 637430
rect 116940 633994 497971 634035
rect 500767 633994 501378 637430
rect 116940 632850 501378 633994
use sky130_fd_pr__diode_pd2nw_05v5_D66R4S  sky130_fd_pr__diode_pd2nw_05v5_D66R4S_4
timestamp 1636132012
transform 1 0 467409 0 1 660132
box -1266 -1266 1266 1266
use sky130_fd_pr__diode_pd2nw_05v5_D66R4S  sky130_fd_pr__diode_pd2nw_05v5_D66R4S_5
timestamp 1636132012
transform 1 0 388543 0 1 660195
box -1266 -1266 1266 1266
use sky130_fd_pr__diode_pd2nw_05v5_D66R4S  sky130_fd_pr__diode_pd2nw_05v5_D66R4S_6
timestamp 1636132012
transform 1 0 392888 0 1 650944
box -1266 -1266 1266 1266
use TopModule_VSW  TopModule_VSW_0
timestamp 1636132012
transform 0 -1 507832 -1 0 682696
box -7310 -3837 33458 29402
use sky130_fd_pr__diode_pd2nw_05v5_3DATV4  sky130_fd_pr__diode_pd2nw_05v5_3DATV4_0
timestamp 1636132012
transform 1 0 496131 0 1 680637
box -866 -866 866 866
use sky130_fd_pr__diode_pd2nw_05v5_D66R4S  sky130_fd_pr__diode_pd2nw_05v5_D66R4S_1
timestamp 1636132012
transform 1 0 526360 0 1 664183
box -1266 -1266 1266 1266
use sky130_fd_pr__diode_pd2nw_05v5_D66R4S  sky130_fd_pr__diode_pd2nw_05v5_D66R4S_2
timestamp 1636132012
transform 1 0 514386 0 1 664601
box -1266 -1266 1266 1266
use sky130_fd_pr__diode_pd2nw_05v5_D66R4S  sky130_fd_pr__diode_pd2nw_05v5_D66R4S_3
timestamp 1636132012
transform 1 0 502641 0 1 686655
box -1266 -1266 1266 1266
use sky130_fd_pr__diode_pd2nw_05v5_3DATV4  sky130_fd_pr__diode_pd2nw_05v5_3DATV4_1
timestamp 1636132012
transform 1 0 497134 0 1 654222
box -866 -866 866 866
use sky130_fd_pr__diode_pd2nw_05v5_D66R4S  sky130_fd_pr__diode_pd2nw_05v5_D66R4S_0
timestamp 1636132012
transform 1 0 387678 0 1 692995
box -1266 -1266 1266 1266
use FINAL_2nov  FINAL_2nov_0
timestamp 1636132012
transform 1 0 129572 0 1 331748
box -114970 -97242 441030 280758
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 2733 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 2733 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 2733 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 2733 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 2733 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 2733 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 2733 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 2733 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 2733 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 2733 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 2733 0 0 0 gpio_analog[2]
port 11 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 2733 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 2733 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 2733 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 2733 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 2733 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 2733 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 2733 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 2733 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 2733 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 2733 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 2733 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 2733 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 2733 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 2733 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 2733 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 2733 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 2733 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 2733 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 2733 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 2733 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 2733 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 2733 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 2733 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 2733 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 2733 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 2733 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 2733 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 4687 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 4687 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 4687 180 0 0 io_analog[3]
port 41 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 4687 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 4687 180 0 0 io_analog[4]
port 42 nsew
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 4687 180 0 0 io_analog[4]
port 42 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 4687 180 0 0 io_analog[4]
port 42 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 4687 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 4687 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 4687 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 4687 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 4687 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 4687 180 0 0 io_analog[5]
port 43 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 4687 180 0 0 io_analog[5]
port 43 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 4687 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 4687 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 4687 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 4687 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 4687 180 0 0 io_analog[6]
port 44 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 4687 180 0 0 io_analog[6]
port 44 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 4687 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 4687 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 4687 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 4687 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 4687 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 4687 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 4687 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 4687 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 4687 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 4687 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 2733 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 2733 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 2733 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 2733 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 2733 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 2733 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 2733 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 2733 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 2733 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 2733 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 2733 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 2733 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 2733 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 2733 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 2733 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 2733 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 2733 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 2733 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 2733 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 2733 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 2733 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 2733 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 2733 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 2733 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 2733 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 2733 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 2733 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 2733 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 2733 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 2733 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 2733 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 2733 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 2733 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 2733 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 2733 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 2733 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 2733 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 2733 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 2733 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 2733 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 2733 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 2733 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 2733 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 2733 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 2733 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 2733 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 2733 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 2733 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 2733 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 2733 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 2733 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 2733 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 2733 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 2733 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 2733 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 2733 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 2733 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 2733 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 2733 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 2733 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 2733 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 2733 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 2733 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 2733 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 2733 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 2733 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 2733 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 2733 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 2733 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 2733 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 2733 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 2733 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 2733 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 2733 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 2733 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 2733 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 2733 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 2733 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 2733 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 2733 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 2733 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 2733 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 2733 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 2733 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 2733 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 2733 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 2733 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 2733 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 2733 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 2733 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 2733 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 2733 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 2733 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 2733 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 2733 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 2733 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 2733 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 2733 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 2733 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 2733 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 2733 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 2733 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 2733 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 2733 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 2733 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 2733 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 2733 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 2733 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 2733 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 2733 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 2733 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 2733 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 2733 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 2733 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 2733 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 2733 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 2733 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 2733 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 2733 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 2733 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 2733 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 2733 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 2733 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 2733 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 2733 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 2733 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 2733 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 2733 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 2733 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 2733 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 2733 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 2733 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 2733 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 2733 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 2733 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 2733 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 2733 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 2733 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 2733 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 2733 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 2733 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 2733 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 2733 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 2733 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 2733 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 2733 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 2733 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 2733 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 2733 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 2733 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 2733 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 2733 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 2733 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 2733 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 2733 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 2733 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 2733 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 2733 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 2733 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 2733 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 2733 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 2733 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 2733 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 2733 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 2733 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 2733 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 2733 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 2733 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 2733 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 2733 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 2733 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 2733 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 2733 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 2733 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 2733 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 2733 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 2733 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 2733 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 2733 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 2733 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 2733 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 2733 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 2733 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 2733 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 2733 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 2733 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 2733 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 2733 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 2733 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 2733 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 2733 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 2733 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 2733 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 2733 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 2733 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 2733 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 2733 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 2733 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 2733 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 2733 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 2733 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 2733 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 2733 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 2733 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 2733 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 2733 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 2733 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 2733 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 2733 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 2733 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 2733 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 2733 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 2733 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 2733 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 2733 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 2733 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 2733 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 2733 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 2733 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 2733 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 2733 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 2733 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 2733 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 2733 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 2733 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 2733 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 2733 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 2733 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 2733 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 2733 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 2733 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 2733 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 2733 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 2733 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 2733 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 2733 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 2733 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 2733 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 2733 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 2733 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 2733 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 2733 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 2733 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 2733 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 2733 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 2733 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 2733 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 2733 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 2733 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 2733 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 2733 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 2733 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 2733 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 2733 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 2733 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 2733 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 2733 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 2733 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 2733 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 2733 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 2733 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 2733 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 2733 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 2733 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 2733 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 2733 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 2733 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 2733 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 2733 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 2733 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 2733 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 2733 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 2733 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 2733 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 2733 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 2733 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 2733 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 2733 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 2733 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 2733 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 2733 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 2733 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 2733 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 2733 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 2733 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 2733 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 2733 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 2733 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 2733 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 2733 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 2733 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 2733 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 2733 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 2733 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 2733 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 2733 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 2733 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 2733 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 2733 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 2733 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 2733 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 2733 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 2733 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 2733 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 2733 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 2733 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 2733 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 2733 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 2733 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 2733 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 2733 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 2733 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 2733 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 2733 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 2733 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 2733 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 2733 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 2733 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 2733 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 2733 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 2733 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 2733 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 2733 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 2733 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 2733 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 2733 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 2733 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 2733 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 2733 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 2733 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 2733 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 2733 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 2733 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 2733 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 2733 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 2733 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 2733 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 2733 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 2733 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 2733 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 2733 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 2733 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 2733 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 2733 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 2733 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 2733 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 2733 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 2733 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 2733 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 2733 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 2733 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 2733 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 2733 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 2733 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 2733 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 2733 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 2733 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 2733 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 2733 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 2733 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 2733 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 2733 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 2733 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 2733 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 2733 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 2733 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 2733 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 2733 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 2733 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 2733 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 2733 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 2733 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 2733 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 2733 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 2733 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 2733 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 2733 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 2733 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 2733 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 2733 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 2733 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 2733 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 2733 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 2733 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 2733 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 2733 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 2733 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 2733 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 2733 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 2733 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 2733 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 2733 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 2733 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 2733 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 2733 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 2733 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 2733 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 2733 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 2733 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 2733 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 2733 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 2733 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 2733 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 2733 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 2733 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 2733 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 2733 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 2733 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 2733 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 2733 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 2733 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 2733 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 2733 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 2733 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 2733 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 2733 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 2733 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 2733 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 2733 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 2733 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 2733 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 2733 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 2733 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 2733 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 2733 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 2733 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 2733 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 2733 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 2733 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 2733 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 2733 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 2733 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 2733 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 2733 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 2733 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 2733 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 2733 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 2733 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 2733 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 2733 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 2733 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 2733 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 2733 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 2733 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 2733 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 2733 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 2733 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 2733 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 2733 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 2733 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 2733 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 2733 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 2733 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 2733 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 2733 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 2733 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 2733 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 2733 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 2733 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 2733 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 2733 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 2733 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 2733 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 2733 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 2733 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 2733 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 2733 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 2733 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 2733 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 2733 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 2733 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 2733 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 2733 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 2733 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 2733 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 2733 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 2733 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 2733 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 2733 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 2733 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 2733 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 2733 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 2733 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 2733 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 2733 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 2733 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 2733 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 2733 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 2733 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 2733 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 2733 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 2733 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 2733 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 2733 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 2733 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 2733 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 2733 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 2733 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 2733 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 2733 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 2733 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 2733 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 2733 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 2733 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 2733 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 2733 0 0 0 vdda2
port 553 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 4687 180 0 0 vssa1
port 554 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 4687 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 2733 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 2733 0 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 2733 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 2733 0 0 0 vssa2
port 555 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 2733 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 2733 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 2733 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 2733 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 2733 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 2733 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 2733 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 2733 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 2733 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 2733 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 2733 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 2733 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 2733 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 2733 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 2733 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 2733 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 2733 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 2733 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 2733 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 2733 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 2733 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 2733 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 2733 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 2733 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 2733 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 2733 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 2733 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 2733 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 2733 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 2733 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 2733 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 2733 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 2733 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 2733 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 2733 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 2733 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 2733 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 2733 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 2733 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 2733 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 2733 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 2733 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 2733 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 2733 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 2733 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 2733 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 2733 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 2733 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 2733 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 2733 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 2733 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 2733 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 2733 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 2733 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 2733 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 2733 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 2733 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 2733 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 2733 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 2733 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 2733 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 2733 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 2733 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 2733 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 2733 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 2733 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 2733 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 2733 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 2733 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 2733 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 2733 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 2733 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 2733 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 2733 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 2733 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 2733 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 2733 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 2733 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 2733 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 2733 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 2733 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 2733 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 2733 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 2733 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 2733 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 2733 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 2733 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 2733 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 2733 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 2733 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 2733 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 2733 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 2733 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 2733 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 2733 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 2733 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 2733 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 2733 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 2733 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 2733 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 2733 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 2733 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 2733 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 2733 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 2733 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 2733 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 2733 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 2733 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 2733 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 2733 90 0 0 wbs_we_i
port 663 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
