magic
tech sky130A
magscale 1 2
timestamp 1635855079
<< pwell >>
rect -191 552 191 638
rect -191 -552 -105 552
rect 105 -552 191 552
rect -191 -638 191 -552
<< psubdiff >>
rect -165 578 -51 612
rect -17 578 17 612
rect 51 578 165 612
rect -165 493 -131 578
rect 131 493 165 578
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect -165 -578 -131 -493
rect 131 -578 165 -493
rect -165 -612 -51 -578
rect -17 -612 17 -578
rect 51 -612 165 -578
<< psubdiffcont >>
rect -51 578 -17 612
rect 17 578 51 612
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect -51 -612 -17 -578
rect 17 -612 51 -578
<< xpolycontact >>
rect -35 50 35 482
rect -35 -482 35 -50
<< ppolyres >>
rect -35 -50 35 50
<< locali >>
rect -165 578 -51 612
rect -17 578 17 612
rect 51 578 165 612
rect -165 493 -131 578
rect 131 493 165 578
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect -165 -51 -131 -17
rect 131 17 165 51
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect -165 -578 -131 -493
rect 131 -578 165 -493
rect -165 -612 -51 -578
rect -17 -612 17 -578
rect 51 -612 165 -578
<< viali >>
rect -17 428 17 462
rect -17 356 17 390
rect -17 284 17 318
rect -17 212 17 246
rect -17 140 17 174
rect -17 68 17 102
rect -17 -103 17 -69
rect -17 -175 17 -141
rect -17 -247 17 -213
rect -17 -319 17 -285
rect -17 -391 17 -357
rect -17 -463 17 -429
<< metal1 >>
rect -25 462 25 476
rect -25 428 -17 462
rect 17 428 25 462
rect -25 390 25 428
rect -25 356 -17 390
rect 17 356 25 390
rect -25 318 25 356
rect -25 284 -17 318
rect 17 284 25 318
rect -25 246 25 284
rect -25 212 -17 246
rect 17 212 25 246
rect -25 174 25 212
rect -25 140 -17 174
rect 17 140 25 174
rect -25 102 25 140
rect -25 68 -17 102
rect 17 68 25 102
rect -25 55 25 68
rect -25 -69 25 -55
rect -25 -103 -17 -69
rect 17 -103 25 -69
rect -25 -141 25 -103
rect -25 -175 -17 -141
rect 17 -175 25 -141
rect -25 -213 25 -175
rect -25 -247 -17 -213
rect 17 -247 25 -213
rect -25 -285 25 -247
rect -25 -319 -17 -285
rect 17 -319 25 -285
rect -25 -357 25 -319
rect -25 -391 -17 -357
rect 17 -391 25 -357
rect -25 -429 25 -391
rect -25 -463 -17 -429
rect 17 -463 25 -429
rect -25 -476 25 -463
<< properties >>
string FIXED_BBOX -148 -595 148 595
<< end >>
