magic
tech sky130A
magscale 1 2
timestamp 1635855079
<< poly >>
rect 1010 110 1042 136
rect 2412 118 2442 134
rect 2506 118 2540 136
rect 898 70 1042 110
rect 2406 68 2540 118
<< locali >>
rect -127 262 1 1117
rect 1170 358 1322 546
rect 1177 300 1317 358
rect 1177 286 1326 300
rect -140 -18 18 262
rect 1177 252 1291 286
rect 1325 252 1326 286
rect 1177 238 1326 252
rect 1177 74 1317 238
rect 1177 14 1319 74
rect 316 -121 1319 14
rect 882 -339 916 -330
rect 882 -411 916 -373
rect 882 -483 916 -445
rect 1027 -481 1319 -121
rect 882 -555 916 -517
rect 882 -627 916 -589
rect 882 -699 916 -661
rect 882 -742 916 -733
rect 1025 -936 1319 -481
<< viali >>
rect 1291 252 1325 286
rect 882 -373 916 -339
rect 882 -445 916 -411
rect 882 -517 916 -483
rect 882 -589 916 -555
rect 882 -661 916 -627
rect 882 -733 916 -699
<< metal1 >>
rect -312 986 -238 1242
rect 2106 1046 2172 1256
rect 222 1036 290 1042
rect 222 986 1060 1036
rect 1526 1034 2562 1046
rect 1432 988 2562 1034
rect 1526 986 2562 988
rect 88 791 152 804
rect 88 739 97 791
rect 149 739 152 791
rect 88 724 152 739
rect 274 791 338 806
rect 274 739 284 791
rect 336 739 338 791
rect 274 726 338 739
rect 474 791 538 806
rect 474 739 478 791
rect 530 739 538 791
rect 474 726 538 739
rect 656 791 720 804
rect 656 739 666 791
rect 718 739 720 791
rect 656 724 720 739
rect 850 791 914 804
rect 850 739 858 791
rect 910 739 914 791
rect 850 724 914 739
rect 1044 791 1108 804
rect 1044 739 1050 791
rect 1102 739 1108 791
rect 1044 724 1108 739
rect 1388 790 1462 804
rect 1388 738 1396 790
rect 1448 738 1462 790
rect 1388 726 1462 738
rect 1578 790 1652 802
rect 1578 738 1588 790
rect 1640 738 1652 790
rect 1578 724 1652 738
rect 1770 790 1844 804
rect 1770 738 1778 790
rect 1830 738 1844 790
rect 1770 726 1844 738
rect 1960 790 2034 802
rect 1960 738 1970 790
rect 2022 738 2034 790
rect 1960 724 2034 738
rect 2152 790 2226 802
rect 2152 738 2162 790
rect 2214 738 2226 790
rect 2152 724 2226 738
rect 2350 790 2424 804
rect 2350 738 2360 790
rect 2412 738 2424 790
rect 2350 726 2424 738
rect 2538 790 2612 802
rect 2538 738 2550 790
rect 2602 738 2612 790
rect 2538 724 2612 738
rect -310 582 -240 592
rect -310 548 -140 582
rect -310 496 -286 548
rect -234 496 -222 548
rect -170 496 -140 548
rect -310 460 -140 496
rect 180 296 248 310
rect 180 244 187 296
rect 239 244 248 296
rect 180 230 248 244
rect 370 296 438 310
rect 370 244 377 296
rect 429 244 438 296
rect 370 230 438 244
rect 562 296 630 310
rect 562 244 571 296
rect 623 244 630 296
rect 562 230 630 244
rect 754 296 822 310
rect 754 244 761 296
rect 813 244 822 296
rect 754 230 822 244
rect 946 296 1014 310
rect 946 244 955 296
rect 1007 244 1014 296
rect 946 230 1014 244
rect 1274 308 1328 312
rect 1274 296 1360 308
rect 1274 286 1296 296
rect 1274 252 1291 286
rect 1274 244 1296 252
rect 1348 244 1360 296
rect 1274 232 1360 244
rect 1484 297 1558 314
rect 1484 245 1492 297
rect 1544 245 1558 297
rect 1274 226 1328 232
rect 1484 226 1558 245
rect 1674 297 1748 316
rect 1674 245 1684 297
rect 1736 245 1748 297
rect 1674 228 1748 245
rect 1862 297 1936 314
rect 1862 245 1874 297
rect 1926 245 1936 297
rect 1862 226 1936 245
rect 2052 297 2126 314
rect 2052 245 2062 297
rect 2114 245 2126 297
rect 2052 226 2126 245
rect 2250 297 2322 316
rect 2446 314 2510 316
rect 2250 245 2260 297
rect 2312 245 2322 297
rect 2250 228 2322 245
rect 2440 296 2510 314
rect 2440 244 2448 296
rect 2500 244 2510 296
rect 2440 234 2510 244
rect 2440 226 2508 234
rect 527 128 753 129
rect 128 110 964 128
rect 128 58 170 110
rect 222 78 964 110
rect 1522 126 2554 128
rect 222 58 260 78
rect 128 46 260 58
rect 527 -547 753 78
rect 1522 74 2556 126
rect 1522 66 2554 74
rect 847 -339 951 -283
rect 847 -348 882 -339
rect 916 -348 951 -339
rect 847 -400 877 -348
rect 929 -400 951 -348
rect 847 -411 951 -400
rect 847 -412 882 -411
rect 916 -412 951 -411
rect 847 -464 877 -412
rect 929 -464 951 -412
rect 847 -476 951 -464
rect 847 -528 877 -476
rect 929 -528 951 -476
rect 847 -540 951 -528
rect 847 -592 877 -540
rect 929 -592 951 -540
rect 847 -604 951 -592
rect 847 -656 877 -604
rect 929 -656 951 -604
rect 847 -661 882 -656
rect 916 -661 951 -656
rect 847 -668 951 -661
rect 847 -720 877 -668
rect 929 -720 951 -668
rect 847 -733 882 -720
rect 916 -733 951 -720
rect 847 -777 951 -733
rect -42 -2424 260 -2422
rect -310 -2491 434 -2424
rect -310 -2863 -13 -2491
rect 231 -2863 434 -2491
rect -310 -2870 434 -2863
rect -42 -2872 260 -2870
<< via1 >>
rect 97 739 149 791
rect 284 739 336 791
rect 478 739 530 791
rect 666 739 718 791
rect 858 739 910 791
rect 1050 739 1102 791
rect 1396 738 1448 790
rect 1588 738 1640 790
rect 1778 738 1830 790
rect 1970 738 2022 790
rect 2162 738 2214 790
rect 2360 738 2412 790
rect 2550 738 2602 790
rect -286 496 -234 548
rect -222 496 -170 548
rect 187 244 239 296
rect 377 244 429 296
rect 571 244 623 296
rect 761 244 813 296
rect 955 244 1007 296
rect 1296 286 1348 296
rect 1296 252 1325 286
rect 1325 252 1348 286
rect 1296 244 1348 252
rect 1492 245 1544 297
rect 1684 245 1736 297
rect 1874 245 1926 297
rect 2062 245 2114 297
rect 2260 245 2312 297
rect 2448 244 2500 296
rect 170 58 222 110
rect 877 -373 882 -348
rect 882 -373 916 -348
rect 916 -373 929 -348
rect 877 -400 929 -373
rect 877 -445 882 -412
rect 882 -445 916 -412
rect 916 -445 929 -412
rect 877 -464 929 -445
rect 877 -483 929 -476
rect 877 -517 882 -483
rect 882 -517 916 -483
rect 916 -517 929 -483
rect 877 -528 929 -517
rect 877 -555 929 -540
rect 877 -589 882 -555
rect 882 -589 916 -555
rect 916 -589 929 -555
rect 877 -592 929 -589
rect 877 -627 929 -604
rect 877 -656 882 -627
rect 882 -656 916 -627
rect 916 -656 929 -627
rect 877 -699 929 -668
rect 877 -720 882 -699
rect 882 -720 916 -699
rect 916 -720 929 -699
rect -13 -2863 231 -2491
<< metal2 >>
rect 1174 798 1320 1400
rect 2538 798 2612 802
rect 90 791 2612 798
rect 90 739 97 791
rect 149 739 284 791
rect 336 739 478 791
rect 530 739 666 791
rect 718 739 858 791
rect 910 739 1050 791
rect 1102 790 2612 791
rect 1102 739 1396 790
rect 90 738 1396 739
rect 1448 738 1588 790
rect 1640 738 1778 790
rect 1830 738 1970 790
rect 2022 738 2162 790
rect 2214 738 2360 790
rect 2412 738 2550 790
rect 2602 738 2612 790
rect 90 732 2612 738
rect 2538 724 2612 732
rect -310 548 324 592
rect -310 496 -286 548
rect -234 496 -222 548
rect -170 496 324 548
rect -310 460 324 496
rect 180 304 322 460
rect 847 304 1014 311
rect 180 296 1014 304
rect 180 244 187 296
rect 239 244 377 296
rect 429 244 571 296
rect 623 244 761 296
rect 813 244 955 296
rect 1007 244 1014 296
rect 180 236 1014 244
rect 128 110 260 120
rect 128 58 170 110
rect 222 58 260 110
rect 128 -2420 260 58
rect 847 -348 1014 236
rect 1282 297 2508 308
rect 1282 296 1492 297
rect 1282 244 1296 296
rect 1348 245 1492 296
rect 1544 245 1684 297
rect 1736 245 1874 297
rect 1926 245 2062 297
rect 2114 245 2260 297
rect 2312 296 2508 297
rect 2312 245 2448 296
rect 1348 244 2448 245
rect 2500 244 2508 296
rect 1282 234 2508 244
rect 1282 232 1356 234
rect 847 -400 877 -348
rect 929 -400 1014 -348
rect 847 -412 1014 -400
rect 847 -464 877 -412
rect 929 -464 1014 -412
rect 847 -476 1014 -464
rect 847 -528 877 -476
rect 929 -528 1014 -476
rect 847 -540 1014 -528
rect 847 -592 877 -540
rect 929 -592 1014 -540
rect 847 -604 1014 -592
rect 847 -656 877 -604
rect 929 -656 1014 -604
rect 847 -668 1014 -656
rect 847 -720 877 -668
rect 929 -720 1014 -668
rect 847 -863 1014 -720
rect 6028 -2420 6668 -2418
rect 128 -2422 6668 -2420
rect -42 -2491 6668 -2422
rect -42 -2863 -13 -2491
rect 231 -2506 6668 -2491
rect 231 -2802 5972 -2506
rect 6588 -2802 6668 -2506
rect 231 -2863 6668 -2802
rect -42 -2872 6668 -2863
<< via2 >>
rect 5972 -2802 6588 -2506
<< metal3 >>
rect 4976 -2418 6654 -2414
rect 4976 -2461 6974 -2418
rect 4976 -2506 6676 -2461
rect 4976 -2802 5972 -2506
rect 6588 -2802 6676 -2506
rect 4976 -2845 6676 -2802
rect 6900 -2845 6974 -2461
rect 4976 -2878 6974 -2845
<< via3 >>
rect 6676 -2845 6900 -2461
<< metal4 >>
rect 6608 -2461 6978 -2116
rect 6608 -2845 6676 -2461
rect 6900 -2845 6978 -2461
rect 6608 -3128 6978 -2845
<< metal5 >>
rect 3922 582 4548 1638
use sky130_fd_pr__nfet_01v8_lvt_KVAFL2  sky130_fd_pr__nfet_01v8_lvt_KVAFL2_0
timestamp 1635855079
transform 1 0 594 0 1 557
box -637 -600 637 600
use sky130_fd_pr__nfet_01v8_lvt_BKUEL6  sky130_fd_pr__nfet_01v8_lvt_BKUEL6_0
timestamp 1635855079
transform -1 0 1995 0 1 556
box -733 -600 733 600
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1635855079
transform 1 0 3295 0 1 -1933
box -3351 -3101 3373 3101
use sky130_fd_pr__res_high_po_0p35_MGFMH8  sky130_fd_pr__res_high_po_0p35_MGFMH8_0
timestamp 1635855079
transform 1 0 -275 0 1 -932
box -191 -2088 191 2088
use sky130_fd_pr__diode_pd2nw_05v5_WW7YB9  sky130_fd_pr__diode_pd2nw_05v5_WW7YB9_0
timestamp 1635855079
transform 1 0 614 0 1 -536
box -466 -466 466 466
<< labels >>
rlabel metal1 s 2136 1230 2136 1230 4 BIAS1
port 1 nsew
rlabel metal5 s 4166 1500 4166 1500 4 RFIN
port 2 nsew
rlabel metal2 s 1224 1388 1224 1388 4 RFOUT_C7T
port 3 nsew
rlabel metal1 s -280 1230 -280 1230 4 VDD
port 4 nsew
rlabel locali s -68 -18 -68 -18 4 VSS
port 5 nsew
<< end >>
