magic
tech sky130A
magscale 1 2
timestamp 1635855079
<< error_p >>
rect -41144 41000 -41084 47200
rect -41064 41000 -41004 47200
rect -34825 41000 -34765 47200
rect -34745 41000 -34685 47200
rect -28506 41000 -28446 47200
rect -28426 41000 -28366 47200
rect -22187 41000 -22127 47200
rect -22107 41000 -22047 47200
rect -15868 41000 -15808 47200
rect -15788 41000 -15728 47200
rect -9549 41000 -9489 47200
rect -9469 41000 -9409 47200
rect -3230 41000 -3170 47200
rect -3150 41000 -3090 47200
rect 3089 41000 3149 47200
rect 3169 41000 3229 47200
rect 9408 41000 9468 47200
rect 9488 41000 9548 47200
rect 15727 41000 15787 47200
rect 15807 41000 15867 47200
rect 22046 41000 22106 47200
rect 22126 41000 22186 47200
rect 28365 41000 28425 47200
rect 28445 41000 28505 47200
rect 34684 41000 34744 47200
rect 34764 41000 34824 47200
rect 41003 41000 41063 47200
rect 41083 41000 41143 47200
rect -41144 34700 -41084 40900
rect -41064 34700 -41004 40900
rect -34825 34700 -34765 40900
rect -34745 34700 -34685 40900
rect -28506 34700 -28446 40900
rect -28426 34700 -28366 40900
rect -22187 34700 -22127 40900
rect -22107 34700 -22047 40900
rect -15868 34700 -15808 40900
rect -15788 34700 -15728 40900
rect -9549 34700 -9489 40900
rect -9469 34700 -9409 40900
rect -3230 34700 -3170 40900
rect -3150 34700 -3090 40900
rect 3089 34700 3149 40900
rect 3169 34700 3229 40900
rect 9408 34700 9468 40900
rect 9488 34700 9548 40900
rect 15727 34700 15787 40900
rect 15807 34700 15867 40900
rect 22046 34700 22106 40900
rect 22126 34700 22186 40900
rect 28365 34700 28425 40900
rect 28445 34700 28505 40900
rect 34684 34700 34744 40900
rect 34764 34700 34824 40900
rect 41003 34700 41063 40900
rect 41083 34700 41143 40900
rect -41144 28400 -41084 34600
rect -41064 28400 -41004 34600
rect -34825 28400 -34765 34600
rect -34745 28400 -34685 34600
rect -28506 28400 -28446 34600
rect -28426 28400 -28366 34600
rect -22187 28400 -22127 34600
rect -22107 28400 -22047 34600
rect -15868 28400 -15808 34600
rect -15788 28400 -15728 34600
rect -9549 28400 -9489 34600
rect -9469 28400 -9409 34600
rect -3230 28400 -3170 34600
rect -3150 28400 -3090 34600
rect 3089 28400 3149 34600
rect 3169 28400 3229 34600
rect 9408 28400 9468 34600
rect 9488 28400 9548 34600
rect 15727 28400 15787 34600
rect 15807 28400 15867 34600
rect 22046 28400 22106 34600
rect 22126 28400 22186 34600
rect 28365 28400 28425 34600
rect 28445 28400 28505 34600
rect 34684 28400 34744 34600
rect 34764 28400 34824 34600
rect 41003 28400 41063 34600
rect 41083 28400 41143 34600
rect -41144 22100 -41084 28300
rect -41064 22100 -41004 28300
rect -34825 22100 -34765 28300
rect -34745 22100 -34685 28300
rect -28506 22100 -28446 28300
rect -28426 22100 -28366 28300
rect -22187 22100 -22127 28300
rect -22107 22100 -22047 28300
rect -15868 22100 -15808 28300
rect -15788 22100 -15728 28300
rect -9549 22100 -9489 28300
rect -9469 22100 -9409 28300
rect -3230 22100 -3170 28300
rect -3150 22100 -3090 28300
rect 3089 22100 3149 28300
rect 3169 22100 3229 28300
rect 9408 22100 9468 28300
rect 9488 22100 9548 28300
rect 15727 22100 15787 28300
rect 15807 22100 15867 28300
rect 22046 22100 22106 28300
rect 22126 22100 22186 28300
rect 28365 22100 28425 28300
rect 28445 22100 28505 28300
rect 34684 22100 34744 28300
rect 34764 22100 34824 28300
rect 41003 22100 41063 28300
rect 41083 22100 41143 28300
rect -41144 15800 -41084 22000
rect -41064 15800 -41004 22000
rect -34825 15800 -34765 22000
rect -34745 15800 -34685 22000
rect -28506 15800 -28446 22000
rect -28426 15800 -28366 22000
rect -22187 15800 -22127 22000
rect -22107 15800 -22047 22000
rect -15868 15800 -15808 22000
rect -15788 15800 -15728 22000
rect -9549 15800 -9489 22000
rect -9469 15800 -9409 22000
rect -3230 15800 -3170 22000
rect -3150 15800 -3090 22000
rect 3089 15800 3149 22000
rect 3169 15800 3229 22000
rect 9408 15800 9468 22000
rect 9488 15800 9548 22000
rect 15727 15800 15787 22000
rect 15807 15800 15867 22000
rect 22046 15800 22106 22000
rect 22126 15800 22186 22000
rect 28365 15800 28425 22000
rect 28445 15800 28505 22000
rect 34684 15800 34744 22000
rect 34764 15800 34824 22000
rect 41003 15800 41063 22000
rect 41083 15800 41143 22000
rect -41144 9500 -41084 15700
rect -41064 9500 -41004 15700
rect -34825 9500 -34765 15700
rect -34745 9500 -34685 15700
rect -28506 9500 -28446 15700
rect -28426 9500 -28366 15700
rect -22187 9500 -22127 15700
rect -22107 9500 -22047 15700
rect -15868 9500 -15808 15700
rect -15788 9500 -15728 15700
rect -9549 9500 -9489 15700
rect -9469 9500 -9409 15700
rect -3230 9500 -3170 15700
rect -3150 9500 -3090 15700
rect 3089 9500 3149 15700
rect 3169 9500 3229 15700
rect 9408 9500 9468 15700
rect 9488 9500 9548 15700
rect 15727 9500 15787 15700
rect 15807 9500 15867 15700
rect 22046 9500 22106 15700
rect 22126 9500 22186 15700
rect 28365 9500 28425 15700
rect 28445 9500 28505 15700
rect 34684 9500 34744 15700
rect 34764 9500 34824 15700
rect 41003 9500 41063 15700
rect 41083 9500 41143 15700
rect -41144 3200 -41084 9400
rect -41064 3200 -41004 9400
rect -34825 3200 -34765 9400
rect -34745 3200 -34685 9400
rect -28506 3200 -28446 9400
rect -28426 3200 -28366 9400
rect -22187 3200 -22127 9400
rect -22107 3200 -22047 9400
rect -15868 3200 -15808 9400
rect -15788 3200 -15728 9400
rect -9549 3200 -9489 9400
rect -9469 3200 -9409 9400
rect -3230 3200 -3170 9400
rect -3150 3200 -3090 9400
rect 3089 3200 3149 9400
rect 3169 3200 3229 9400
rect 9408 3200 9468 9400
rect 9488 3200 9548 9400
rect 15727 3200 15787 9400
rect 15807 3200 15867 9400
rect 22046 3200 22106 9400
rect 22126 3200 22186 9400
rect 28365 3200 28425 9400
rect 28445 3200 28505 9400
rect 34684 3200 34744 9400
rect 34764 3200 34824 9400
rect 41003 3200 41063 9400
rect 41083 3200 41143 9400
rect -41144 -3100 -41084 3100
rect -41064 -3100 -41004 3100
rect -34825 -3100 -34765 3100
rect -34745 -3100 -34685 3100
rect -28506 -3100 -28446 3100
rect -28426 -3100 -28366 3100
rect -22187 -3100 -22127 3100
rect -22107 -3100 -22047 3100
rect -15868 -3100 -15808 3100
rect -15788 -3100 -15728 3100
rect -9549 -3100 -9489 3100
rect -9469 -3100 -9409 3100
rect -3230 -3100 -3170 3100
rect -3150 -3100 -3090 3100
rect 3089 -3100 3149 3100
rect 3169 -3100 3229 3100
rect 9408 -3100 9468 3100
rect 9488 -3100 9548 3100
rect 15727 -3100 15787 3100
rect 15807 -3100 15867 3100
rect 22046 -3100 22106 3100
rect 22126 -3100 22186 3100
rect 28365 -3100 28425 3100
rect 28445 -3100 28505 3100
rect 34684 -3100 34744 3100
rect 34764 -3100 34824 3100
rect 41003 -3100 41063 3100
rect 41083 -3100 41143 3100
rect -41144 -9400 -41084 -3200
rect -41064 -9400 -41004 -3200
rect -34825 -9400 -34765 -3200
rect -34745 -9400 -34685 -3200
rect -28506 -9400 -28446 -3200
rect -28426 -9400 -28366 -3200
rect -22187 -9400 -22127 -3200
rect -22107 -9400 -22047 -3200
rect -15868 -9400 -15808 -3200
rect -15788 -9400 -15728 -3200
rect -9549 -9400 -9489 -3200
rect -9469 -9400 -9409 -3200
rect -3230 -9400 -3170 -3200
rect -3150 -9400 -3090 -3200
rect 3089 -9400 3149 -3200
rect 3169 -9400 3229 -3200
rect 9408 -9400 9468 -3200
rect 9488 -9400 9548 -3200
rect 15727 -9400 15787 -3200
rect 15807 -9400 15867 -3200
rect 22046 -9400 22106 -3200
rect 22126 -9400 22186 -3200
rect 28365 -9400 28425 -3200
rect 28445 -9400 28505 -3200
rect 34684 -9400 34744 -3200
rect 34764 -9400 34824 -3200
rect 41003 -9400 41063 -3200
rect 41083 -9400 41143 -3200
rect -41144 -15700 -41084 -9500
rect -41064 -15700 -41004 -9500
rect -34825 -15700 -34765 -9500
rect -34745 -15700 -34685 -9500
rect -28506 -15700 -28446 -9500
rect -28426 -15700 -28366 -9500
rect -22187 -15700 -22127 -9500
rect -22107 -15700 -22047 -9500
rect -15868 -15700 -15808 -9500
rect -15788 -15700 -15728 -9500
rect -9549 -15700 -9489 -9500
rect -9469 -15700 -9409 -9500
rect -3230 -15700 -3170 -9500
rect -3150 -15700 -3090 -9500
rect 3089 -15700 3149 -9500
rect 3169 -15700 3229 -9500
rect 9408 -15700 9468 -9500
rect 9488 -15700 9548 -9500
rect 15727 -15700 15787 -9500
rect 15807 -15700 15867 -9500
rect 22046 -15700 22106 -9500
rect 22126 -15700 22186 -9500
rect 28365 -15700 28425 -9500
rect 28445 -15700 28505 -9500
rect 34684 -15700 34744 -9500
rect 34764 -15700 34824 -9500
rect 41003 -15700 41063 -9500
rect 41083 -15700 41143 -9500
rect -41144 -22000 -41084 -15800
rect -41064 -22000 -41004 -15800
rect -34825 -22000 -34765 -15800
rect -34745 -22000 -34685 -15800
rect -28506 -22000 -28446 -15800
rect -28426 -22000 -28366 -15800
rect -22187 -22000 -22127 -15800
rect -22107 -22000 -22047 -15800
rect -15868 -22000 -15808 -15800
rect -15788 -22000 -15728 -15800
rect -9549 -22000 -9489 -15800
rect -9469 -22000 -9409 -15800
rect -3230 -22000 -3170 -15800
rect -3150 -22000 -3090 -15800
rect 3089 -22000 3149 -15800
rect 3169 -22000 3229 -15800
rect 9408 -22000 9468 -15800
rect 9488 -22000 9548 -15800
rect 15727 -22000 15787 -15800
rect 15807 -22000 15867 -15800
rect 22046 -22000 22106 -15800
rect 22126 -22000 22186 -15800
rect 28365 -22000 28425 -15800
rect 28445 -22000 28505 -15800
rect 34684 -22000 34744 -15800
rect 34764 -22000 34824 -15800
rect 41003 -22000 41063 -15800
rect 41083 -22000 41143 -15800
rect -41144 -28300 -41084 -22100
rect -41064 -28300 -41004 -22100
rect -34825 -28300 -34765 -22100
rect -34745 -28300 -34685 -22100
rect -28506 -28300 -28446 -22100
rect -28426 -28300 -28366 -22100
rect -22187 -28300 -22127 -22100
rect -22107 -28300 -22047 -22100
rect -15868 -28300 -15808 -22100
rect -15788 -28300 -15728 -22100
rect -9549 -28300 -9489 -22100
rect -9469 -28300 -9409 -22100
rect -3230 -28300 -3170 -22100
rect -3150 -28300 -3090 -22100
rect 3089 -28300 3149 -22100
rect 3169 -28300 3229 -22100
rect 9408 -28300 9468 -22100
rect 9488 -28300 9548 -22100
rect 15727 -28300 15787 -22100
rect 15807 -28300 15867 -22100
rect 22046 -28300 22106 -22100
rect 22126 -28300 22186 -22100
rect 28365 -28300 28425 -22100
rect 28445 -28300 28505 -22100
rect 34684 -28300 34744 -22100
rect 34764 -28300 34824 -22100
rect 41003 -28300 41063 -22100
rect 41083 -28300 41143 -22100
rect -41144 -34600 -41084 -28400
rect -41064 -34600 -41004 -28400
rect -34825 -34600 -34765 -28400
rect -34745 -34600 -34685 -28400
rect -28506 -34600 -28446 -28400
rect -28426 -34600 -28366 -28400
rect -22187 -34600 -22127 -28400
rect -22107 -34600 -22047 -28400
rect -15868 -34600 -15808 -28400
rect -15788 -34600 -15728 -28400
rect -9549 -34600 -9489 -28400
rect -9469 -34600 -9409 -28400
rect -3230 -34600 -3170 -28400
rect -3150 -34600 -3090 -28400
rect 3089 -34600 3149 -28400
rect 3169 -34600 3229 -28400
rect 9408 -34600 9468 -28400
rect 9488 -34600 9548 -28400
rect 15727 -34600 15787 -28400
rect 15807 -34600 15867 -28400
rect 22046 -34600 22106 -28400
rect 22126 -34600 22186 -28400
rect 28365 -34600 28425 -28400
rect 28445 -34600 28505 -28400
rect 34684 -34600 34744 -28400
rect 34764 -34600 34824 -28400
rect 41003 -34600 41063 -28400
rect 41083 -34600 41143 -28400
rect -41144 -40900 -41084 -34700
rect -41064 -40900 -41004 -34700
rect -34825 -40900 -34765 -34700
rect -34745 -40900 -34685 -34700
rect -28506 -40900 -28446 -34700
rect -28426 -40900 -28366 -34700
rect -22187 -40900 -22127 -34700
rect -22107 -40900 -22047 -34700
rect -15868 -40900 -15808 -34700
rect -15788 -40900 -15728 -34700
rect -9549 -40900 -9489 -34700
rect -9469 -40900 -9409 -34700
rect -3230 -40900 -3170 -34700
rect -3150 -40900 -3090 -34700
rect 3089 -40900 3149 -34700
rect 3169 -40900 3229 -34700
rect 9408 -40900 9468 -34700
rect 9488 -40900 9548 -34700
rect 15727 -40900 15787 -34700
rect 15807 -40900 15867 -34700
rect 22046 -40900 22106 -34700
rect 22126 -40900 22186 -34700
rect 28365 -40900 28425 -34700
rect 28445 -40900 28505 -34700
rect 34684 -40900 34744 -34700
rect 34764 -40900 34824 -34700
rect 41003 -40900 41063 -34700
rect 41083 -40900 41143 -34700
rect -41144 -47200 -41084 -41000
rect -41064 -47200 -41004 -41000
rect -34825 -47200 -34765 -41000
rect -34745 -47200 -34685 -41000
rect -28506 -47200 -28446 -41000
rect -28426 -47200 -28366 -41000
rect -22187 -47200 -22127 -41000
rect -22107 -47200 -22047 -41000
rect -15868 -47200 -15808 -41000
rect -15788 -47200 -15728 -41000
rect -9549 -47200 -9489 -41000
rect -9469 -47200 -9409 -41000
rect -3230 -47200 -3170 -41000
rect -3150 -47200 -3090 -41000
rect 3089 -47200 3149 -41000
rect 3169 -47200 3229 -41000
rect 9408 -47200 9468 -41000
rect 9488 -47200 9548 -41000
rect 15727 -47200 15787 -41000
rect 15807 -47200 15867 -41000
rect 22046 -47200 22106 -41000
rect 22126 -47200 22186 -41000
rect 28365 -47200 28425 -41000
rect 28445 -47200 28505 -41000
rect 34684 -47200 34744 -41000
rect 34764 -47200 34824 -41000
rect 41003 -47200 41063 -41000
rect 41083 -47200 41143 -41000
<< metal3 >>
rect -47383 47172 -41084 47200
rect -47383 47108 -41168 47172
rect -41104 47108 -41084 47172
rect -47383 47092 -41084 47108
rect -47383 47028 -41168 47092
rect -41104 47028 -41084 47092
rect -47383 47012 -41084 47028
rect -47383 46948 -41168 47012
rect -41104 46948 -41084 47012
rect -47383 46932 -41084 46948
rect -47383 46868 -41168 46932
rect -41104 46868 -41084 46932
rect -47383 46852 -41084 46868
rect -47383 46788 -41168 46852
rect -41104 46788 -41084 46852
rect -47383 46772 -41084 46788
rect -47383 46708 -41168 46772
rect -41104 46708 -41084 46772
rect -47383 46692 -41084 46708
rect -47383 46628 -41168 46692
rect -41104 46628 -41084 46692
rect -47383 46612 -41084 46628
rect -47383 46548 -41168 46612
rect -41104 46548 -41084 46612
rect -47383 46532 -41084 46548
rect -47383 46468 -41168 46532
rect -41104 46468 -41084 46532
rect -47383 46452 -41084 46468
rect -47383 46388 -41168 46452
rect -41104 46388 -41084 46452
rect -47383 46372 -41084 46388
rect -47383 46308 -41168 46372
rect -41104 46308 -41084 46372
rect -47383 46292 -41084 46308
rect -47383 46228 -41168 46292
rect -41104 46228 -41084 46292
rect -47383 46212 -41084 46228
rect -47383 46148 -41168 46212
rect -41104 46148 -41084 46212
rect -47383 46132 -41084 46148
rect -47383 46068 -41168 46132
rect -41104 46068 -41084 46132
rect -47383 46052 -41084 46068
rect -47383 45988 -41168 46052
rect -41104 45988 -41084 46052
rect -47383 45972 -41084 45988
rect -47383 45908 -41168 45972
rect -41104 45908 -41084 45972
rect -47383 45892 -41084 45908
rect -47383 45828 -41168 45892
rect -41104 45828 -41084 45892
rect -47383 45812 -41084 45828
rect -47383 45748 -41168 45812
rect -41104 45748 -41084 45812
rect -47383 45732 -41084 45748
rect -47383 45668 -41168 45732
rect -41104 45668 -41084 45732
rect -47383 45652 -41084 45668
rect -47383 45588 -41168 45652
rect -41104 45588 -41084 45652
rect -47383 45572 -41084 45588
rect -47383 45508 -41168 45572
rect -41104 45508 -41084 45572
rect -47383 45492 -41084 45508
rect -47383 45428 -41168 45492
rect -41104 45428 -41084 45492
rect -47383 45412 -41084 45428
rect -47383 45348 -41168 45412
rect -41104 45348 -41084 45412
rect -47383 45332 -41084 45348
rect -47383 45268 -41168 45332
rect -41104 45268 -41084 45332
rect -47383 45252 -41084 45268
rect -47383 45188 -41168 45252
rect -41104 45188 -41084 45252
rect -47383 45172 -41084 45188
rect -47383 45108 -41168 45172
rect -41104 45108 -41084 45172
rect -47383 45092 -41084 45108
rect -47383 45028 -41168 45092
rect -41104 45028 -41084 45092
rect -47383 45012 -41084 45028
rect -47383 44948 -41168 45012
rect -41104 44948 -41084 45012
rect -47383 44932 -41084 44948
rect -47383 44868 -41168 44932
rect -41104 44868 -41084 44932
rect -47383 44852 -41084 44868
rect -47383 44788 -41168 44852
rect -41104 44788 -41084 44852
rect -47383 44772 -41084 44788
rect -47383 44708 -41168 44772
rect -41104 44708 -41084 44772
rect -47383 44692 -41084 44708
rect -47383 44628 -41168 44692
rect -41104 44628 -41084 44692
rect -47383 44612 -41084 44628
rect -47383 44548 -41168 44612
rect -41104 44548 -41084 44612
rect -47383 44532 -41084 44548
rect -47383 44468 -41168 44532
rect -41104 44468 -41084 44532
rect -47383 44452 -41084 44468
rect -47383 44388 -41168 44452
rect -41104 44388 -41084 44452
rect -47383 44372 -41084 44388
rect -47383 44308 -41168 44372
rect -41104 44308 -41084 44372
rect -47383 44292 -41084 44308
rect -47383 44228 -41168 44292
rect -41104 44228 -41084 44292
rect -47383 44212 -41084 44228
rect -47383 44148 -41168 44212
rect -41104 44148 -41084 44212
rect -47383 44132 -41084 44148
rect -47383 44068 -41168 44132
rect -41104 44068 -41084 44132
rect -47383 44052 -41084 44068
rect -47383 43988 -41168 44052
rect -41104 43988 -41084 44052
rect -47383 43972 -41084 43988
rect -47383 43908 -41168 43972
rect -41104 43908 -41084 43972
rect -47383 43892 -41084 43908
rect -47383 43828 -41168 43892
rect -41104 43828 -41084 43892
rect -47383 43812 -41084 43828
rect -47383 43748 -41168 43812
rect -41104 43748 -41084 43812
rect -47383 43732 -41084 43748
rect -47383 43668 -41168 43732
rect -41104 43668 -41084 43732
rect -47383 43652 -41084 43668
rect -47383 43588 -41168 43652
rect -41104 43588 -41084 43652
rect -47383 43572 -41084 43588
rect -47383 43508 -41168 43572
rect -41104 43508 -41084 43572
rect -47383 43492 -41084 43508
rect -47383 43428 -41168 43492
rect -41104 43428 -41084 43492
rect -47383 43412 -41084 43428
rect -47383 43348 -41168 43412
rect -41104 43348 -41084 43412
rect -47383 43332 -41084 43348
rect -47383 43268 -41168 43332
rect -41104 43268 -41084 43332
rect -47383 43252 -41084 43268
rect -47383 43188 -41168 43252
rect -41104 43188 -41084 43252
rect -47383 43172 -41084 43188
rect -47383 43108 -41168 43172
rect -41104 43108 -41084 43172
rect -47383 43092 -41084 43108
rect -47383 43028 -41168 43092
rect -41104 43028 -41084 43092
rect -47383 43012 -41084 43028
rect -47383 42948 -41168 43012
rect -41104 42948 -41084 43012
rect -47383 42932 -41084 42948
rect -47383 42868 -41168 42932
rect -41104 42868 -41084 42932
rect -47383 42852 -41084 42868
rect -47383 42788 -41168 42852
rect -41104 42788 -41084 42852
rect -47383 42772 -41084 42788
rect -47383 42708 -41168 42772
rect -41104 42708 -41084 42772
rect -47383 42692 -41084 42708
rect -47383 42628 -41168 42692
rect -41104 42628 -41084 42692
rect -47383 42612 -41084 42628
rect -47383 42548 -41168 42612
rect -41104 42548 -41084 42612
rect -47383 42532 -41084 42548
rect -47383 42468 -41168 42532
rect -41104 42468 -41084 42532
rect -47383 42452 -41084 42468
rect -47383 42388 -41168 42452
rect -41104 42388 -41084 42452
rect -47383 42372 -41084 42388
rect -47383 42308 -41168 42372
rect -41104 42308 -41084 42372
rect -47383 42292 -41084 42308
rect -47383 42228 -41168 42292
rect -41104 42228 -41084 42292
rect -47383 42212 -41084 42228
rect -47383 42148 -41168 42212
rect -41104 42148 -41084 42212
rect -47383 42132 -41084 42148
rect -47383 42068 -41168 42132
rect -41104 42068 -41084 42132
rect -47383 42052 -41084 42068
rect -47383 41988 -41168 42052
rect -41104 41988 -41084 42052
rect -47383 41972 -41084 41988
rect -47383 41908 -41168 41972
rect -41104 41908 -41084 41972
rect -47383 41892 -41084 41908
rect -47383 41828 -41168 41892
rect -41104 41828 -41084 41892
rect -47383 41812 -41084 41828
rect -47383 41748 -41168 41812
rect -41104 41748 -41084 41812
rect -47383 41732 -41084 41748
rect -47383 41668 -41168 41732
rect -41104 41668 -41084 41732
rect -47383 41652 -41084 41668
rect -47383 41588 -41168 41652
rect -41104 41588 -41084 41652
rect -47383 41572 -41084 41588
rect -47383 41508 -41168 41572
rect -41104 41508 -41084 41572
rect -47383 41492 -41084 41508
rect -47383 41428 -41168 41492
rect -41104 41428 -41084 41492
rect -47383 41412 -41084 41428
rect -47383 41348 -41168 41412
rect -41104 41348 -41084 41412
rect -47383 41332 -41084 41348
rect -47383 41268 -41168 41332
rect -41104 41268 -41084 41332
rect -47383 41252 -41084 41268
rect -47383 41188 -41168 41252
rect -41104 41188 -41084 41252
rect -47383 41172 -41084 41188
rect -47383 41108 -41168 41172
rect -41104 41108 -41084 41172
rect -47383 41092 -41084 41108
rect -47383 41028 -41168 41092
rect -41104 41028 -41084 41092
rect -47383 41000 -41084 41028
rect -41064 47172 -34765 47200
rect -41064 47108 -34849 47172
rect -34785 47108 -34765 47172
rect -41064 47092 -34765 47108
rect -41064 47028 -34849 47092
rect -34785 47028 -34765 47092
rect -41064 47012 -34765 47028
rect -41064 46948 -34849 47012
rect -34785 46948 -34765 47012
rect -41064 46932 -34765 46948
rect -41064 46868 -34849 46932
rect -34785 46868 -34765 46932
rect -41064 46852 -34765 46868
rect -41064 46788 -34849 46852
rect -34785 46788 -34765 46852
rect -41064 46772 -34765 46788
rect -41064 46708 -34849 46772
rect -34785 46708 -34765 46772
rect -41064 46692 -34765 46708
rect -41064 46628 -34849 46692
rect -34785 46628 -34765 46692
rect -41064 46612 -34765 46628
rect -41064 46548 -34849 46612
rect -34785 46548 -34765 46612
rect -41064 46532 -34765 46548
rect -41064 46468 -34849 46532
rect -34785 46468 -34765 46532
rect -41064 46452 -34765 46468
rect -41064 46388 -34849 46452
rect -34785 46388 -34765 46452
rect -41064 46372 -34765 46388
rect -41064 46308 -34849 46372
rect -34785 46308 -34765 46372
rect -41064 46292 -34765 46308
rect -41064 46228 -34849 46292
rect -34785 46228 -34765 46292
rect -41064 46212 -34765 46228
rect -41064 46148 -34849 46212
rect -34785 46148 -34765 46212
rect -41064 46132 -34765 46148
rect -41064 46068 -34849 46132
rect -34785 46068 -34765 46132
rect -41064 46052 -34765 46068
rect -41064 45988 -34849 46052
rect -34785 45988 -34765 46052
rect -41064 45972 -34765 45988
rect -41064 45908 -34849 45972
rect -34785 45908 -34765 45972
rect -41064 45892 -34765 45908
rect -41064 45828 -34849 45892
rect -34785 45828 -34765 45892
rect -41064 45812 -34765 45828
rect -41064 45748 -34849 45812
rect -34785 45748 -34765 45812
rect -41064 45732 -34765 45748
rect -41064 45668 -34849 45732
rect -34785 45668 -34765 45732
rect -41064 45652 -34765 45668
rect -41064 45588 -34849 45652
rect -34785 45588 -34765 45652
rect -41064 45572 -34765 45588
rect -41064 45508 -34849 45572
rect -34785 45508 -34765 45572
rect -41064 45492 -34765 45508
rect -41064 45428 -34849 45492
rect -34785 45428 -34765 45492
rect -41064 45412 -34765 45428
rect -41064 45348 -34849 45412
rect -34785 45348 -34765 45412
rect -41064 45332 -34765 45348
rect -41064 45268 -34849 45332
rect -34785 45268 -34765 45332
rect -41064 45252 -34765 45268
rect -41064 45188 -34849 45252
rect -34785 45188 -34765 45252
rect -41064 45172 -34765 45188
rect -41064 45108 -34849 45172
rect -34785 45108 -34765 45172
rect -41064 45092 -34765 45108
rect -41064 45028 -34849 45092
rect -34785 45028 -34765 45092
rect -41064 45012 -34765 45028
rect -41064 44948 -34849 45012
rect -34785 44948 -34765 45012
rect -41064 44932 -34765 44948
rect -41064 44868 -34849 44932
rect -34785 44868 -34765 44932
rect -41064 44852 -34765 44868
rect -41064 44788 -34849 44852
rect -34785 44788 -34765 44852
rect -41064 44772 -34765 44788
rect -41064 44708 -34849 44772
rect -34785 44708 -34765 44772
rect -41064 44692 -34765 44708
rect -41064 44628 -34849 44692
rect -34785 44628 -34765 44692
rect -41064 44612 -34765 44628
rect -41064 44548 -34849 44612
rect -34785 44548 -34765 44612
rect -41064 44532 -34765 44548
rect -41064 44468 -34849 44532
rect -34785 44468 -34765 44532
rect -41064 44452 -34765 44468
rect -41064 44388 -34849 44452
rect -34785 44388 -34765 44452
rect -41064 44372 -34765 44388
rect -41064 44308 -34849 44372
rect -34785 44308 -34765 44372
rect -41064 44292 -34765 44308
rect -41064 44228 -34849 44292
rect -34785 44228 -34765 44292
rect -41064 44212 -34765 44228
rect -41064 44148 -34849 44212
rect -34785 44148 -34765 44212
rect -41064 44132 -34765 44148
rect -41064 44068 -34849 44132
rect -34785 44068 -34765 44132
rect -41064 44052 -34765 44068
rect -41064 43988 -34849 44052
rect -34785 43988 -34765 44052
rect -41064 43972 -34765 43988
rect -41064 43908 -34849 43972
rect -34785 43908 -34765 43972
rect -41064 43892 -34765 43908
rect -41064 43828 -34849 43892
rect -34785 43828 -34765 43892
rect -41064 43812 -34765 43828
rect -41064 43748 -34849 43812
rect -34785 43748 -34765 43812
rect -41064 43732 -34765 43748
rect -41064 43668 -34849 43732
rect -34785 43668 -34765 43732
rect -41064 43652 -34765 43668
rect -41064 43588 -34849 43652
rect -34785 43588 -34765 43652
rect -41064 43572 -34765 43588
rect -41064 43508 -34849 43572
rect -34785 43508 -34765 43572
rect -41064 43492 -34765 43508
rect -41064 43428 -34849 43492
rect -34785 43428 -34765 43492
rect -41064 43412 -34765 43428
rect -41064 43348 -34849 43412
rect -34785 43348 -34765 43412
rect -41064 43332 -34765 43348
rect -41064 43268 -34849 43332
rect -34785 43268 -34765 43332
rect -41064 43252 -34765 43268
rect -41064 43188 -34849 43252
rect -34785 43188 -34765 43252
rect -41064 43172 -34765 43188
rect -41064 43108 -34849 43172
rect -34785 43108 -34765 43172
rect -41064 43092 -34765 43108
rect -41064 43028 -34849 43092
rect -34785 43028 -34765 43092
rect -41064 43012 -34765 43028
rect -41064 42948 -34849 43012
rect -34785 42948 -34765 43012
rect -41064 42932 -34765 42948
rect -41064 42868 -34849 42932
rect -34785 42868 -34765 42932
rect -41064 42852 -34765 42868
rect -41064 42788 -34849 42852
rect -34785 42788 -34765 42852
rect -41064 42772 -34765 42788
rect -41064 42708 -34849 42772
rect -34785 42708 -34765 42772
rect -41064 42692 -34765 42708
rect -41064 42628 -34849 42692
rect -34785 42628 -34765 42692
rect -41064 42612 -34765 42628
rect -41064 42548 -34849 42612
rect -34785 42548 -34765 42612
rect -41064 42532 -34765 42548
rect -41064 42468 -34849 42532
rect -34785 42468 -34765 42532
rect -41064 42452 -34765 42468
rect -41064 42388 -34849 42452
rect -34785 42388 -34765 42452
rect -41064 42372 -34765 42388
rect -41064 42308 -34849 42372
rect -34785 42308 -34765 42372
rect -41064 42292 -34765 42308
rect -41064 42228 -34849 42292
rect -34785 42228 -34765 42292
rect -41064 42212 -34765 42228
rect -41064 42148 -34849 42212
rect -34785 42148 -34765 42212
rect -41064 42132 -34765 42148
rect -41064 42068 -34849 42132
rect -34785 42068 -34765 42132
rect -41064 42052 -34765 42068
rect -41064 41988 -34849 42052
rect -34785 41988 -34765 42052
rect -41064 41972 -34765 41988
rect -41064 41908 -34849 41972
rect -34785 41908 -34765 41972
rect -41064 41892 -34765 41908
rect -41064 41828 -34849 41892
rect -34785 41828 -34765 41892
rect -41064 41812 -34765 41828
rect -41064 41748 -34849 41812
rect -34785 41748 -34765 41812
rect -41064 41732 -34765 41748
rect -41064 41668 -34849 41732
rect -34785 41668 -34765 41732
rect -41064 41652 -34765 41668
rect -41064 41588 -34849 41652
rect -34785 41588 -34765 41652
rect -41064 41572 -34765 41588
rect -41064 41508 -34849 41572
rect -34785 41508 -34765 41572
rect -41064 41492 -34765 41508
rect -41064 41428 -34849 41492
rect -34785 41428 -34765 41492
rect -41064 41412 -34765 41428
rect -41064 41348 -34849 41412
rect -34785 41348 -34765 41412
rect -41064 41332 -34765 41348
rect -41064 41268 -34849 41332
rect -34785 41268 -34765 41332
rect -41064 41252 -34765 41268
rect -41064 41188 -34849 41252
rect -34785 41188 -34765 41252
rect -41064 41172 -34765 41188
rect -41064 41108 -34849 41172
rect -34785 41108 -34765 41172
rect -41064 41092 -34765 41108
rect -41064 41028 -34849 41092
rect -34785 41028 -34765 41092
rect -41064 41000 -34765 41028
rect -34745 47172 -28446 47200
rect -34745 47108 -28530 47172
rect -28466 47108 -28446 47172
rect -34745 47092 -28446 47108
rect -34745 47028 -28530 47092
rect -28466 47028 -28446 47092
rect -34745 47012 -28446 47028
rect -34745 46948 -28530 47012
rect -28466 46948 -28446 47012
rect -34745 46932 -28446 46948
rect -34745 46868 -28530 46932
rect -28466 46868 -28446 46932
rect -34745 46852 -28446 46868
rect -34745 46788 -28530 46852
rect -28466 46788 -28446 46852
rect -34745 46772 -28446 46788
rect -34745 46708 -28530 46772
rect -28466 46708 -28446 46772
rect -34745 46692 -28446 46708
rect -34745 46628 -28530 46692
rect -28466 46628 -28446 46692
rect -34745 46612 -28446 46628
rect -34745 46548 -28530 46612
rect -28466 46548 -28446 46612
rect -34745 46532 -28446 46548
rect -34745 46468 -28530 46532
rect -28466 46468 -28446 46532
rect -34745 46452 -28446 46468
rect -34745 46388 -28530 46452
rect -28466 46388 -28446 46452
rect -34745 46372 -28446 46388
rect -34745 46308 -28530 46372
rect -28466 46308 -28446 46372
rect -34745 46292 -28446 46308
rect -34745 46228 -28530 46292
rect -28466 46228 -28446 46292
rect -34745 46212 -28446 46228
rect -34745 46148 -28530 46212
rect -28466 46148 -28446 46212
rect -34745 46132 -28446 46148
rect -34745 46068 -28530 46132
rect -28466 46068 -28446 46132
rect -34745 46052 -28446 46068
rect -34745 45988 -28530 46052
rect -28466 45988 -28446 46052
rect -34745 45972 -28446 45988
rect -34745 45908 -28530 45972
rect -28466 45908 -28446 45972
rect -34745 45892 -28446 45908
rect -34745 45828 -28530 45892
rect -28466 45828 -28446 45892
rect -34745 45812 -28446 45828
rect -34745 45748 -28530 45812
rect -28466 45748 -28446 45812
rect -34745 45732 -28446 45748
rect -34745 45668 -28530 45732
rect -28466 45668 -28446 45732
rect -34745 45652 -28446 45668
rect -34745 45588 -28530 45652
rect -28466 45588 -28446 45652
rect -34745 45572 -28446 45588
rect -34745 45508 -28530 45572
rect -28466 45508 -28446 45572
rect -34745 45492 -28446 45508
rect -34745 45428 -28530 45492
rect -28466 45428 -28446 45492
rect -34745 45412 -28446 45428
rect -34745 45348 -28530 45412
rect -28466 45348 -28446 45412
rect -34745 45332 -28446 45348
rect -34745 45268 -28530 45332
rect -28466 45268 -28446 45332
rect -34745 45252 -28446 45268
rect -34745 45188 -28530 45252
rect -28466 45188 -28446 45252
rect -34745 45172 -28446 45188
rect -34745 45108 -28530 45172
rect -28466 45108 -28446 45172
rect -34745 45092 -28446 45108
rect -34745 45028 -28530 45092
rect -28466 45028 -28446 45092
rect -34745 45012 -28446 45028
rect -34745 44948 -28530 45012
rect -28466 44948 -28446 45012
rect -34745 44932 -28446 44948
rect -34745 44868 -28530 44932
rect -28466 44868 -28446 44932
rect -34745 44852 -28446 44868
rect -34745 44788 -28530 44852
rect -28466 44788 -28446 44852
rect -34745 44772 -28446 44788
rect -34745 44708 -28530 44772
rect -28466 44708 -28446 44772
rect -34745 44692 -28446 44708
rect -34745 44628 -28530 44692
rect -28466 44628 -28446 44692
rect -34745 44612 -28446 44628
rect -34745 44548 -28530 44612
rect -28466 44548 -28446 44612
rect -34745 44532 -28446 44548
rect -34745 44468 -28530 44532
rect -28466 44468 -28446 44532
rect -34745 44452 -28446 44468
rect -34745 44388 -28530 44452
rect -28466 44388 -28446 44452
rect -34745 44372 -28446 44388
rect -34745 44308 -28530 44372
rect -28466 44308 -28446 44372
rect -34745 44292 -28446 44308
rect -34745 44228 -28530 44292
rect -28466 44228 -28446 44292
rect -34745 44212 -28446 44228
rect -34745 44148 -28530 44212
rect -28466 44148 -28446 44212
rect -34745 44132 -28446 44148
rect -34745 44068 -28530 44132
rect -28466 44068 -28446 44132
rect -34745 44052 -28446 44068
rect -34745 43988 -28530 44052
rect -28466 43988 -28446 44052
rect -34745 43972 -28446 43988
rect -34745 43908 -28530 43972
rect -28466 43908 -28446 43972
rect -34745 43892 -28446 43908
rect -34745 43828 -28530 43892
rect -28466 43828 -28446 43892
rect -34745 43812 -28446 43828
rect -34745 43748 -28530 43812
rect -28466 43748 -28446 43812
rect -34745 43732 -28446 43748
rect -34745 43668 -28530 43732
rect -28466 43668 -28446 43732
rect -34745 43652 -28446 43668
rect -34745 43588 -28530 43652
rect -28466 43588 -28446 43652
rect -34745 43572 -28446 43588
rect -34745 43508 -28530 43572
rect -28466 43508 -28446 43572
rect -34745 43492 -28446 43508
rect -34745 43428 -28530 43492
rect -28466 43428 -28446 43492
rect -34745 43412 -28446 43428
rect -34745 43348 -28530 43412
rect -28466 43348 -28446 43412
rect -34745 43332 -28446 43348
rect -34745 43268 -28530 43332
rect -28466 43268 -28446 43332
rect -34745 43252 -28446 43268
rect -34745 43188 -28530 43252
rect -28466 43188 -28446 43252
rect -34745 43172 -28446 43188
rect -34745 43108 -28530 43172
rect -28466 43108 -28446 43172
rect -34745 43092 -28446 43108
rect -34745 43028 -28530 43092
rect -28466 43028 -28446 43092
rect -34745 43012 -28446 43028
rect -34745 42948 -28530 43012
rect -28466 42948 -28446 43012
rect -34745 42932 -28446 42948
rect -34745 42868 -28530 42932
rect -28466 42868 -28446 42932
rect -34745 42852 -28446 42868
rect -34745 42788 -28530 42852
rect -28466 42788 -28446 42852
rect -34745 42772 -28446 42788
rect -34745 42708 -28530 42772
rect -28466 42708 -28446 42772
rect -34745 42692 -28446 42708
rect -34745 42628 -28530 42692
rect -28466 42628 -28446 42692
rect -34745 42612 -28446 42628
rect -34745 42548 -28530 42612
rect -28466 42548 -28446 42612
rect -34745 42532 -28446 42548
rect -34745 42468 -28530 42532
rect -28466 42468 -28446 42532
rect -34745 42452 -28446 42468
rect -34745 42388 -28530 42452
rect -28466 42388 -28446 42452
rect -34745 42372 -28446 42388
rect -34745 42308 -28530 42372
rect -28466 42308 -28446 42372
rect -34745 42292 -28446 42308
rect -34745 42228 -28530 42292
rect -28466 42228 -28446 42292
rect -34745 42212 -28446 42228
rect -34745 42148 -28530 42212
rect -28466 42148 -28446 42212
rect -34745 42132 -28446 42148
rect -34745 42068 -28530 42132
rect -28466 42068 -28446 42132
rect -34745 42052 -28446 42068
rect -34745 41988 -28530 42052
rect -28466 41988 -28446 42052
rect -34745 41972 -28446 41988
rect -34745 41908 -28530 41972
rect -28466 41908 -28446 41972
rect -34745 41892 -28446 41908
rect -34745 41828 -28530 41892
rect -28466 41828 -28446 41892
rect -34745 41812 -28446 41828
rect -34745 41748 -28530 41812
rect -28466 41748 -28446 41812
rect -34745 41732 -28446 41748
rect -34745 41668 -28530 41732
rect -28466 41668 -28446 41732
rect -34745 41652 -28446 41668
rect -34745 41588 -28530 41652
rect -28466 41588 -28446 41652
rect -34745 41572 -28446 41588
rect -34745 41508 -28530 41572
rect -28466 41508 -28446 41572
rect -34745 41492 -28446 41508
rect -34745 41428 -28530 41492
rect -28466 41428 -28446 41492
rect -34745 41412 -28446 41428
rect -34745 41348 -28530 41412
rect -28466 41348 -28446 41412
rect -34745 41332 -28446 41348
rect -34745 41268 -28530 41332
rect -28466 41268 -28446 41332
rect -34745 41252 -28446 41268
rect -34745 41188 -28530 41252
rect -28466 41188 -28446 41252
rect -34745 41172 -28446 41188
rect -34745 41108 -28530 41172
rect -28466 41108 -28446 41172
rect -34745 41092 -28446 41108
rect -34745 41028 -28530 41092
rect -28466 41028 -28446 41092
rect -34745 41000 -28446 41028
rect -28426 47172 -22127 47200
rect -28426 47108 -22211 47172
rect -22147 47108 -22127 47172
rect -28426 47092 -22127 47108
rect -28426 47028 -22211 47092
rect -22147 47028 -22127 47092
rect -28426 47012 -22127 47028
rect -28426 46948 -22211 47012
rect -22147 46948 -22127 47012
rect -28426 46932 -22127 46948
rect -28426 46868 -22211 46932
rect -22147 46868 -22127 46932
rect -28426 46852 -22127 46868
rect -28426 46788 -22211 46852
rect -22147 46788 -22127 46852
rect -28426 46772 -22127 46788
rect -28426 46708 -22211 46772
rect -22147 46708 -22127 46772
rect -28426 46692 -22127 46708
rect -28426 46628 -22211 46692
rect -22147 46628 -22127 46692
rect -28426 46612 -22127 46628
rect -28426 46548 -22211 46612
rect -22147 46548 -22127 46612
rect -28426 46532 -22127 46548
rect -28426 46468 -22211 46532
rect -22147 46468 -22127 46532
rect -28426 46452 -22127 46468
rect -28426 46388 -22211 46452
rect -22147 46388 -22127 46452
rect -28426 46372 -22127 46388
rect -28426 46308 -22211 46372
rect -22147 46308 -22127 46372
rect -28426 46292 -22127 46308
rect -28426 46228 -22211 46292
rect -22147 46228 -22127 46292
rect -28426 46212 -22127 46228
rect -28426 46148 -22211 46212
rect -22147 46148 -22127 46212
rect -28426 46132 -22127 46148
rect -28426 46068 -22211 46132
rect -22147 46068 -22127 46132
rect -28426 46052 -22127 46068
rect -28426 45988 -22211 46052
rect -22147 45988 -22127 46052
rect -28426 45972 -22127 45988
rect -28426 45908 -22211 45972
rect -22147 45908 -22127 45972
rect -28426 45892 -22127 45908
rect -28426 45828 -22211 45892
rect -22147 45828 -22127 45892
rect -28426 45812 -22127 45828
rect -28426 45748 -22211 45812
rect -22147 45748 -22127 45812
rect -28426 45732 -22127 45748
rect -28426 45668 -22211 45732
rect -22147 45668 -22127 45732
rect -28426 45652 -22127 45668
rect -28426 45588 -22211 45652
rect -22147 45588 -22127 45652
rect -28426 45572 -22127 45588
rect -28426 45508 -22211 45572
rect -22147 45508 -22127 45572
rect -28426 45492 -22127 45508
rect -28426 45428 -22211 45492
rect -22147 45428 -22127 45492
rect -28426 45412 -22127 45428
rect -28426 45348 -22211 45412
rect -22147 45348 -22127 45412
rect -28426 45332 -22127 45348
rect -28426 45268 -22211 45332
rect -22147 45268 -22127 45332
rect -28426 45252 -22127 45268
rect -28426 45188 -22211 45252
rect -22147 45188 -22127 45252
rect -28426 45172 -22127 45188
rect -28426 45108 -22211 45172
rect -22147 45108 -22127 45172
rect -28426 45092 -22127 45108
rect -28426 45028 -22211 45092
rect -22147 45028 -22127 45092
rect -28426 45012 -22127 45028
rect -28426 44948 -22211 45012
rect -22147 44948 -22127 45012
rect -28426 44932 -22127 44948
rect -28426 44868 -22211 44932
rect -22147 44868 -22127 44932
rect -28426 44852 -22127 44868
rect -28426 44788 -22211 44852
rect -22147 44788 -22127 44852
rect -28426 44772 -22127 44788
rect -28426 44708 -22211 44772
rect -22147 44708 -22127 44772
rect -28426 44692 -22127 44708
rect -28426 44628 -22211 44692
rect -22147 44628 -22127 44692
rect -28426 44612 -22127 44628
rect -28426 44548 -22211 44612
rect -22147 44548 -22127 44612
rect -28426 44532 -22127 44548
rect -28426 44468 -22211 44532
rect -22147 44468 -22127 44532
rect -28426 44452 -22127 44468
rect -28426 44388 -22211 44452
rect -22147 44388 -22127 44452
rect -28426 44372 -22127 44388
rect -28426 44308 -22211 44372
rect -22147 44308 -22127 44372
rect -28426 44292 -22127 44308
rect -28426 44228 -22211 44292
rect -22147 44228 -22127 44292
rect -28426 44212 -22127 44228
rect -28426 44148 -22211 44212
rect -22147 44148 -22127 44212
rect -28426 44132 -22127 44148
rect -28426 44068 -22211 44132
rect -22147 44068 -22127 44132
rect -28426 44052 -22127 44068
rect -28426 43988 -22211 44052
rect -22147 43988 -22127 44052
rect -28426 43972 -22127 43988
rect -28426 43908 -22211 43972
rect -22147 43908 -22127 43972
rect -28426 43892 -22127 43908
rect -28426 43828 -22211 43892
rect -22147 43828 -22127 43892
rect -28426 43812 -22127 43828
rect -28426 43748 -22211 43812
rect -22147 43748 -22127 43812
rect -28426 43732 -22127 43748
rect -28426 43668 -22211 43732
rect -22147 43668 -22127 43732
rect -28426 43652 -22127 43668
rect -28426 43588 -22211 43652
rect -22147 43588 -22127 43652
rect -28426 43572 -22127 43588
rect -28426 43508 -22211 43572
rect -22147 43508 -22127 43572
rect -28426 43492 -22127 43508
rect -28426 43428 -22211 43492
rect -22147 43428 -22127 43492
rect -28426 43412 -22127 43428
rect -28426 43348 -22211 43412
rect -22147 43348 -22127 43412
rect -28426 43332 -22127 43348
rect -28426 43268 -22211 43332
rect -22147 43268 -22127 43332
rect -28426 43252 -22127 43268
rect -28426 43188 -22211 43252
rect -22147 43188 -22127 43252
rect -28426 43172 -22127 43188
rect -28426 43108 -22211 43172
rect -22147 43108 -22127 43172
rect -28426 43092 -22127 43108
rect -28426 43028 -22211 43092
rect -22147 43028 -22127 43092
rect -28426 43012 -22127 43028
rect -28426 42948 -22211 43012
rect -22147 42948 -22127 43012
rect -28426 42932 -22127 42948
rect -28426 42868 -22211 42932
rect -22147 42868 -22127 42932
rect -28426 42852 -22127 42868
rect -28426 42788 -22211 42852
rect -22147 42788 -22127 42852
rect -28426 42772 -22127 42788
rect -28426 42708 -22211 42772
rect -22147 42708 -22127 42772
rect -28426 42692 -22127 42708
rect -28426 42628 -22211 42692
rect -22147 42628 -22127 42692
rect -28426 42612 -22127 42628
rect -28426 42548 -22211 42612
rect -22147 42548 -22127 42612
rect -28426 42532 -22127 42548
rect -28426 42468 -22211 42532
rect -22147 42468 -22127 42532
rect -28426 42452 -22127 42468
rect -28426 42388 -22211 42452
rect -22147 42388 -22127 42452
rect -28426 42372 -22127 42388
rect -28426 42308 -22211 42372
rect -22147 42308 -22127 42372
rect -28426 42292 -22127 42308
rect -28426 42228 -22211 42292
rect -22147 42228 -22127 42292
rect -28426 42212 -22127 42228
rect -28426 42148 -22211 42212
rect -22147 42148 -22127 42212
rect -28426 42132 -22127 42148
rect -28426 42068 -22211 42132
rect -22147 42068 -22127 42132
rect -28426 42052 -22127 42068
rect -28426 41988 -22211 42052
rect -22147 41988 -22127 42052
rect -28426 41972 -22127 41988
rect -28426 41908 -22211 41972
rect -22147 41908 -22127 41972
rect -28426 41892 -22127 41908
rect -28426 41828 -22211 41892
rect -22147 41828 -22127 41892
rect -28426 41812 -22127 41828
rect -28426 41748 -22211 41812
rect -22147 41748 -22127 41812
rect -28426 41732 -22127 41748
rect -28426 41668 -22211 41732
rect -22147 41668 -22127 41732
rect -28426 41652 -22127 41668
rect -28426 41588 -22211 41652
rect -22147 41588 -22127 41652
rect -28426 41572 -22127 41588
rect -28426 41508 -22211 41572
rect -22147 41508 -22127 41572
rect -28426 41492 -22127 41508
rect -28426 41428 -22211 41492
rect -22147 41428 -22127 41492
rect -28426 41412 -22127 41428
rect -28426 41348 -22211 41412
rect -22147 41348 -22127 41412
rect -28426 41332 -22127 41348
rect -28426 41268 -22211 41332
rect -22147 41268 -22127 41332
rect -28426 41252 -22127 41268
rect -28426 41188 -22211 41252
rect -22147 41188 -22127 41252
rect -28426 41172 -22127 41188
rect -28426 41108 -22211 41172
rect -22147 41108 -22127 41172
rect -28426 41092 -22127 41108
rect -28426 41028 -22211 41092
rect -22147 41028 -22127 41092
rect -28426 41000 -22127 41028
rect -22107 47172 -15808 47200
rect -22107 47108 -15892 47172
rect -15828 47108 -15808 47172
rect -22107 47092 -15808 47108
rect -22107 47028 -15892 47092
rect -15828 47028 -15808 47092
rect -22107 47012 -15808 47028
rect -22107 46948 -15892 47012
rect -15828 46948 -15808 47012
rect -22107 46932 -15808 46948
rect -22107 46868 -15892 46932
rect -15828 46868 -15808 46932
rect -22107 46852 -15808 46868
rect -22107 46788 -15892 46852
rect -15828 46788 -15808 46852
rect -22107 46772 -15808 46788
rect -22107 46708 -15892 46772
rect -15828 46708 -15808 46772
rect -22107 46692 -15808 46708
rect -22107 46628 -15892 46692
rect -15828 46628 -15808 46692
rect -22107 46612 -15808 46628
rect -22107 46548 -15892 46612
rect -15828 46548 -15808 46612
rect -22107 46532 -15808 46548
rect -22107 46468 -15892 46532
rect -15828 46468 -15808 46532
rect -22107 46452 -15808 46468
rect -22107 46388 -15892 46452
rect -15828 46388 -15808 46452
rect -22107 46372 -15808 46388
rect -22107 46308 -15892 46372
rect -15828 46308 -15808 46372
rect -22107 46292 -15808 46308
rect -22107 46228 -15892 46292
rect -15828 46228 -15808 46292
rect -22107 46212 -15808 46228
rect -22107 46148 -15892 46212
rect -15828 46148 -15808 46212
rect -22107 46132 -15808 46148
rect -22107 46068 -15892 46132
rect -15828 46068 -15808 46132
rect -22107 46052 -15808 46068
rect -22107 45988 -15892 46052
rect -15828 45988 -15808 46052
rect -22107 45972 -15808 45988
rect -22107 45908 -15892 45972
rect -15828 45908 -15808 45972
rect -22107 45892 -15808 45908
rect -22107 45828 -15892 45892
rect -15828 45828 -15808 45892
rect -22107 45812 -15808 45828
rect -22107 45748 -15892 45812
rect -15828 45748 -15808 45812
rect -22107 45732 -15808 45748
rect -22107 45668 -15892 45732
rect -15828 45668 -15808 45732
rect -22107 45652 -15808 45668
rect -22107 45588 -15892 45652
rect -15828 45588 -15808 45652
rect -22107 45572 -15808 45588
rect -22107 45508 -15892 45572
rect -15828 45508 -15808 45572
rect -22107 45492 -15808 45508
rect -22107 45428 -15892 45492
rect -15828 45428 -15808 45492
rect -22107 45412 -15808 45428
rect -22107 45348 -15892 45412
rect -15828 45348 -15808 45412
rect -22107 45332 -15808 45348
rect -22107 45268 -15892 45332
rect -15828 45268 -15808 45332
rect -22107 45252 -15808 45268
rect -22107 45188 -15892 45252
rect -15828 45188 -15808 45252
rect -22107 45172 -15808 45188
rect -22107 45108 -15892 45172
rect -15828 45108 -15808 45172
rect -22107 45092 -15808 45108
rect -22107 45028 -15892 45092
rect -15828 45028 -15808 45092
rect -22107 45012 -15808 45028
rect -22107 44948 -15892 45012
rect -15828 44948 -15808 45012
rect -22107 44932 -15808 44948
rect -22107 44868 -15892 44932
rect -15828 44868 -15808 44932
rect -22107 44852 -15808 44868
rect -22107 44788 -15892 44852
rect -15828 44788 -15808 44852
rect -22107 44772 -15808 44788
rect -22107 44708 -15892 44772
rect -15828 44708 -15808 44772
rect -22107 44692 -15808 44708
rect -22107 44628 -15892 44692
rect -15828 44628 -15808 44692
rect -22107 44612 -15808 44628
rect -22107 44548 -15892 44612
rect -15828 44548 -15808 44612
rect -22107 44532 -15808 44548
rect -22107 44468 -15892 44532
rect -15828 44468 -15808 44532
rect -22107 44452 -15808 44468
rect -22107 44388 -15892 44452
rect -15828 44388 -15808 44452
rect -22107 44372 -15808 44388
rect -22107 44308 -15892 44372
rect -15828 44308 -15808 44372
rect -22107 44292 -15808 44308
rect -22107 44228 -15892 44292
rect -15828 44228 -15808 44292
rect -22107 44212 -15808 44228
rect -22107 44148 -15892 44212
rect -15828 44148 -15808 44212
rect -22107 44132 -15808 44148
rect -22107 44068 -15892 44132
rect -15828 44068 -15808 44132
rect -22107 44052 -15808 44068
rect -22107 43988 -15892 44052
rect -15828 43988 -15808 44052
rect -22107 43972 -15808 43988
rect -22107 43908 -15892 43972
rect -15828 43908 -15808 43972
rect -22107 43892 -15808 43908
rect -22107 43828 -15892 43892
rect -15828 43828 -15808 43892
rect -22107 43812 -15808 43828
rect -22107 43748 -15892 43812
rect -15828 43748 -15808 43812
rect -22107 43732 -15808 43748
rect -22107 43668 -15892 43732
rect -15828 43668 -15808 43732
rect -22107 43652 -15808 43668
rect -22107 43588 -15892 43652
rect -15828 43588 -15808 43652
rect -22107 43572 -15808 43588
rect -22107 43508 -15892 43572
rect -15828 43508 -15808 43572
rect -22107 43492 -15808 43508
rect -22107 43428 -15892 43492
rect -15828 43428 -15808 43492
rect -22107 43412 -15808 43428
rect -22107 43348 -15892 43412
rect -15828 43348 -15808 43412
rect -22107 43332 -15808 43348
rect -22107 43268 -15892 43332
rect -15828 43268 -15808 43332
rect -22107 43252 -15808 43268
rect -22107 43188 -15892 43252
rect -15828 43188 -15808 43252
rect -22107 43172 -15808 43188
rect -22107 43108 -15892 43172
rect -15828 43108 -15808 43172
rect -22107 43092 -15808 43108
rect -22107 43028 -15892 43092
rect -15828 43028 -15808 43092
rect -22107 43012 -15808 43028
rect -22107 42948 -15892 43012
rect -15828 42948 -15808 43012
rect -22107 42932 -15808 42948
rect -22107 42868 -15892 42932
rect -15828 42868 -15808 42932
rect -22107 42852 -15808 42868
rect -22107 42788 -15892 42852
rect -15828 42788 -15808 42852
rect -22107 42772 -15808 42788
rect -22107 42708 -15892 42772
rect -15828 42708 -15808 42772
rect -22107 42692 -15808 42708
rect -22107 42628 -15892 42692
rect -15828 42628 -15808 42692
rect -22107 42612 -15808 42628
rect -22107 42548 -15892 42612
rect -15828 42548 -15808 42612
rect -22107 42532 -15808 42548
rect -22107 42468 -15892 42532
rect -15828 42468 -15808 42532
rect -22107 42452 -15808 42468
rect -22107 42388 -15892 42452
rect -15828 42388 -15808 42452
rect -22107 42372 -15808 42388
rect -22107 42308 -15892 42372
rect -15828 42308 -15808 42372
rect -22107 42292 -15808 42308
rect -22107 42228 -15892 42292
rect -15828 42228 -15808 42292
rect -22107 42212 -15808 42228
rect -22107 42148 -15892 42212
rect -15828 42148 -15808 42212
rect -22107 42132 -15808 42148
rect -22107 42068 -15892 42132
rect -15828 42068 -15808 42132
rect -22107 42052 -15808 42068
rect -22107 41988 -15892 42052
rect -15828 41988 -15808 42052
rect -22107 41972 -15808 41988
rect -22107 41908 -15892 41972
rect -15828 41908 -15808 41972
rect -22107 41892 -15808 41908
rect -22107 41828 -15892 41892
rect -15828 41828 -15808 41892
rect -22107 41812 -15808 41828
rect -22107 41748 -15892 41812
rect -15828 41748 -15808 41812
rect -22107 41732 -15808 41748
rect -22107 41668 -15892 41732
rect -15828 41668 -15808 41732
rect -22107 41652 -15808 41668
rect -22107 41588 -15892 41652
rect -15828 41588 -15808 41652
rect -22107 41572 -15808 41588
rect -22107 41508 -15892 41572
rect -15828 41508 -15808 41572
rect -22107 41492 -15808 41508
rect -22107 41428 -15892 41492
rect -15828 41428 -15808 41492
rect -22107 41412 -15808 41428
rect -22107 41348 -15892 41412
rect -15828 41348 -15808 41412
rect -22107 41332 -15808 41348
rect -22107 41268 -15892 41332
rect -15828 41268 -15808 41332
rect -22107 41252 -15808 41268
rect -22107 41188 -15892 41252
rect -15828 41188 -15808 41252
rect -22107 41172 -15808 41188
rect -22107 41108 -15892 41172
rect -15828 41108 -15808 41172
rect -22107 41092 -15808 41108
rect -22107 41028 -15892 41092
rect -15828 41028 -15808 41092
rect -22107 41000 -15808 41028
rect -15788 47172 -9489 47200
rect -15788 47108 -9573 47172
rect -9509 47108 -9489 47172
rect -15788 47092 -9489 47108
rect -15788 47028 -9573 47092
rect -9509 47028 -9489 47092
rect -15788 47012 -9489 47028
rect -15788 46948 -9573 47012
rect -9509 46948 -9489 47012
rect -15788 46932 -9489 46948
rect -15788 46868 -9573 46932
rect -9509 46868 -9489 46932
rect -15788 46852 -9489 46868
rect -15788 46788 -9573 46852
rect -9509 46788 -9489 46852
rect -15788 46772 -9489 46788
rect -15788 46708 -9573 46772
rect -9509 46708 -9489 46772
rect -15788 46692 -9489 46708
rect -15788 46628 -9573 46692
rect -9509 46628 -9489 46692
rect -15788 46612 -9489 46628
rect -15788 46548 -9573 46612
rect -9509 46548 -9489 46612
rect -15788 46532 -9489 46548
rect -15788 46468 -9573 46532
rect -9509 46468 -9489 46532
rect -15788 46452 -9489 46468
rect -15788 46388 -9573 46452
rect -9509 46388 -9489 46452
rect -15788 46372 -9489 46388
rect -15788 46308 -9573 46372
rect -9509 46308 -9489 46372
rect -15788 46292 -9489 46308
rect -15788 46228 -9573 46292
rect -9509 46228 -9489 46292
rect -15788 46212 -9489 46228
rect -15788 46148 -9573 46212
rect -9509 46148 -9489 46212
rect -15788 46132 -9489 46148
rect -15788 46068 -9573 46132
rect -9509 46068 -9489 46132
rect -15788 46052 -9489 46068
rect -15788 45988 -9573 46052
rect -9509 45988 -9489 46052
rect -15788 45972 -9489 45988
rect -15788 45908 -9573 45972
rect -9509 45908 -9489 45972
rect -15788 45892 -9489 45908
rect -15788 45828 -9573 45892
rect -9509 45828 -9489 45892
rect -15788 45812 -9489 45828
rect -15788 45748 -9573 45812
rect -9509 45748 -9489 45812
rect -15788 45732 -9489 45748
rect -15788 45668 -9573 45732
rect -9509 45668 -9489 45732
rect -15788 45652 -9489 45668
rect -15788 45588 -9573 45652
rect -9509 45588 -9489 45652
rect -15788 45572 -9489 45588
rect -15788 45508 -9573 45572
rect -9509 45508 -9489 45572
rect -15788 45492 -9489 45508
rect -15788 45428 -9573 45492
rect -9509 45428 -9489 45492
rect -15788 45412 -9489 45428
rect -15788 45348 -9573 45412
rect -9509 45348 -9489 45412
rect -15788 45332 -9489 45348
rect -15788 45268 -9573 45332
rect -9509 45268 -9489 45332
rect -15788 45252 -9489 45268
rect -15788 45188 -9573 45252
rect -9509 45188 -9489 45252
rect -15788 45172 -9489 45188
rect -15788 45108 -9573 45172
rect -9509 45108 -9489 45172
rect -15788 45092 -9489 45108
rect -15788 45028 -9573 45092
rect -9509 45028 -9489 45092
rect -15788 45012 -9489 45028
rect -15788 44948 -9573 45012
rect -9509 44948 -9489 45012
rect -15788 44932 -9489 44948
rect -15788 44868 -9573 44932
rect -9509 44868 -9489 44932
rect -15788 44852 -9489 44868
rect -15788 44788 -9573 44852
rect -9509 44788 -9489 44852
rect -15788 44772 -9489 44788
rect -15788 44708 -9573 44772
rect -9509 44708 -9489 44772
rect -15788 44692 -9489 44708
rect -15788 44628 -9573 44692
rect -9509 44628 -9489 44692
rect -15788 44612 -9489 44628
rect -15788 44548 -9573 44612
rect -9509 44548 -9489 44612
rect -15788 44532 -9489 44548
rect -15788 44468 -9573 44532
rect -9509 44468 -9489 44532
rect -15788 44452 -9489 44468
rect -15788 44388 -9573 44452
rect -9509 44388 -9489 44452
rect -15788 44372 -9489 44388
rect -15788 44308 -9573 44372
rect -9509 44308 -9489 44372
rect -15788 44292 -9489 44308
rect -15788 44228 -9573 44292
rect -9509 44228 -9489 44292
rect -15788 44212 -9489 44228
rect -15788 44148 -9573 44212
rect -9509 44148 -9489 44212
rect -15788 44132 -9489 44148
rect -15788 44068 -9573 44132
rect -9509 44068 -9489 44132
rect -15788 44052 -9489 44068
rect -15788 43988 -9573 44052
rect -9509 43988 -9489 44052
rect -15788 43972 -9489 43988
rect -15788 43908 -9573 43972
rect -9509 43908 -9489 43972
rect -15788 43892 -9489 43908
rect -15788 43828 -9573 43892
rect -9509 43828 -9489 43892
rect -15788 43812 -9489 43828
rect -15788 43748 -9573 43812
rect -9509 43748 -9489 43812
rect -15788 43732 -9489 43748
rect -15788 43668 -9573 43732
rect -9509 43668 -9489 43732
rect -15788 43652 -9489 43668
rect -15788 43588 -9573 43652
rect -9509 43588 -9489 43652
rect -15788 43572 -9489 43588
rect -15788 43508 -9573 43572
rect -9509 43508 -9489 43572
rect -15788 43492 -9489 43508
rect -15788 43428 -9573 43492
rect -9509 43428 -9489 43492
rect -15788 43412 -9489 43428
rect -15788 43348 -9573 43412
rect -9509 43348 -9489 43412
rect -15788 43332 -9489 43348
rect -15788 43268 -9573 43332
rect -9509 43268 -9489 43332
rect -15788 43252 -9489 43268
rect -15788 43188 -9573 43252
rect -9509 43188 -9489 43252
rect -15788 43172 -9489 43188
rect -15788 43108 -9573 43172
rect -9509 43108 -9489 43172
rect -15788 43092 -9489 43108
rect -15788 43028 -9573 43092
rect -9509 43028 -9489 43092
rect -15788 43012 -9489 43028
rect -15788 42948 -9573 43012
rect -9509 42948 -9489 43012
rect -15788 42932 -9489 42948
rect -15788 42868 -9573 42932
rect -9509 42868 -9489 42932
rect -15788 42852 -9489 42868
rect -15788 42788 -9573 42852
rect -9509 42788 -9489 42852
rect -15788 42772 -9489 42788
rect -15788 42708 -9573 42772
rect -9509 42708 -9489 42772
rect -15788 42692 -9489 42708
rect -15788 42628 -9573 42692
rect -9509 42628 -9489 42692
rect -15788 42612 -9489 42628
rect -15788 42548 -9573 42612
rect -9509 42548 -9489 42612
rect -15788 42532 -9489 42548
rect -15788 42468 -9573 42532
rect -9509 42468 -9489 42532
rect -15788 42452 -9489 42468
rect -15788 42388 -9573 42452
rect -9509 42388 -9489 42452
rect -15788 42372 -9489 42388
rect -15788 42308 -9573 42372
rect -9509 42308 -9489 42372
rect -15788 42292 -9489 42308
rect -15788 42228 -9573 42292
rect -9509 42228 -9489 42292
rect -15788 42212 -9489 42228
rect -15788 42148 -9573 42212
rect -9509 42148 -9489 42212
rect -15788 42132 -9489 42148
rect -15788 42068 -9573 42132
rect -9509 42068 -9489 42132
rect -15788 42052 -9489 42068
rect -15788 41988 -9573 42052
rect -9509 41988 -9489 42052
rect -15788 41972 -9489 41988
rect -15788 41908 -9573 41972
rect -9509 41908 -9489 41972
rect -15788 41892 -9489 41908
rect -15788 41828 -9573 41892
rect -9509 41828 -9489 41892
rect -15788 41812 -9489 41828
rect -15788 41748 -9573 41812
rect -9509 41748 -9489 41812
rect -15788 41732 -9489 41748
rect -15788 41668 -9573 41732
rect -9509 41668 -9489 41732
rect -15788 41652 -9489 41668
rect -15788 41588 -9573 41652
rect -9509 41588 -9489 41652
rect -15788 41572 -9489 41588
rect -15788 41508 -9573 41572
rect -9509 41508 -9489 41572
rect -15788 41492 -9489 41508
rect -15788 41428 -9573 41492
rect -9509 41428 -9489 41492
rect -15788 41412 -9489 41428
rect -15788 41348 -9573 41412
rect -9509 41348 -9489 41412
rect -15788 41332 -9489 41348
rect -15788 41268 -9573 41332
rect -9509 41268 -9489 41332
rect -15788 41252 -9489 41268
rect -15788 41188 -9573 41252
rect -9509 41188 -9489 41252
rect -15788 41172 -9489 41188
rect -15788 41108 -9573 41172
rect -9509 41108 -9489 41172
rect -15788 41092 -9489 41108
rect -15788 41028 -9573 41092
rect -9509 41028 -9489 41092
rect -15788 41000 -9489 41028
rect -9469 47172 -3170 47200
rect -9469 47108 -3254 47172
rect -3190 47108 -3170 47172
rect -9469 47092 -3170 47108
rect -9469 47028 -3254 47092
rect -3190 47028 -3170 47092
rect -9469 47012 -3170 47028
rect -9469 46948 -3254 47012
rect -3190 46948 -3170 47012
rect -9469 46932 -3170 46948
rect -9469 46868 -3254 46932
rect -3190 46868 -3170 46932
rect -9469 46852 -3170 46868
rect -9469 46788 -3254 46852
rect -3190 46788 -3170 46852
rect -9469 46772 -3170 46788
rect -9469 46708 -3254 46772
rect -3190 46708 -3170 46772
rect -9469 46692 -3170 46708
rect -9469 46628 -3254 46692
rect -3190 46628 -3170 46692
rect -9469 46612 -3170 46628
rect -9469 46548 -3254 46612
rect -3190 46548 -3170 46612
rect -9469 46532 -3170 46548
rect -9469 46468 -3254 46532
rect -3190 46468 -3170 46532
rect -9469 46452 -3170 46468
rect -9469 46388 -3254 46452
rect -3190 46388 -3170 46452
rect -9469 46372 -3170 46388
rect -9469 46308 -3254 46372
rect -3190 46308 -3170 46372
rect -9469 46292 -3170 46308
rect -9469 46228 -3254 46292
rect -3190 46228 -3170 46292
rect -9469 46212 -3170 46228
rect -9469 46148 -3254 46212
rect -3190 46148 -3170 46212
rect -9469 46132 -3170 46148
rect -9469 46068 -3254 46132
rect -3190 46068 -3170 46132
rect -9469 46052 -3170 46068
rect -9469 45988 -3254 46052
rect -3190 45988 -3170 46052
rect -9469 45972 -3170 45988
rect -9469 45908 -3254 45972
rect -3190 45908 -3170 45972
rect -9469 45892 -3170 45908
rect -9469 45828 -3254 45892
rect -3190 45828 -3170 45892
rect -9469 45812 -3170 45828
rect -9469 45748 -3254 45812
rect -3190 45748 -3170 45812
rect -9469 45732 -3170 45748
rect -9469 45668 -3254 45732
rect -3190 45668 -3170 45732
rect -9469 45652 -3170 45668
rect -9469 45588 -3254 45652
rect -3190 45588 -3170 45652
rect -9469 45572 -3170 45588
rect -9469 45508 -3254 45572
rect -3190 45508 -3170 45572
rect -9469 45492 -3170 45508
rect -9469 45428 -3254 45492
rect -3190 45428 -3170 45492
rect -9469 45412 -3170 45428
rect -9469 45348 -3254 45412
rect -3190 45348 -3170 45412
rect -9469 45332 -3170 45348
rect -9469 45268 -3254 45332
rect -3190 45268 -3170 45332
rect -9469 45252 -3170 45268
rect -9469 45188 -3254 45252
rect -3190 45188 -3170 45252
rect -9469 45172 -3170 45188
rect -9469 45108 -3254 45172
rect -3190 45108 -3170 45172
rect -9469 45092 -3170 45108
rect -9469 45028 -3254 45092
rect -3190 45028 -3170 45092
rect -9469 45012 -3170 45028
rect -9469 44948 -3254 45012
rect -3190 44948 -3170 45012
rect -9469 44932 -3170 44948
rect -9469 44868 -3254 44932
rect -3190 44868 -3170 44932
rect -9469 44852 -3170 44868
rect -9469 44788 -3254 44852
rect -3190 44788 -3170 44852
rect -9469 44772 -3170 44788
rect -9469 44708 -3254 44772
rect -3190 44708 -3170 44772
rect -9469 44692 -3170 44708
rect -9469 44628 -3254 44692
rect -3190 44628 -3170 44692
rect -9469 44612 -3170 44628
rect -9469 44548 -3254 44612
rect -3190 44548 -3170 44612
rect -9469 44532 -3170 44548
rect -9469 44468 -3254 44532
rect -3190 44468 -3170 44532
rect -9469 44452 -3170 44468
rect -9469 44388 -3254 44452
rect -3190 44388 -3170 44452
rect -9469 44372 -3170 44388
rect -9469 44308 -3254 44372
rect -3190 44308 -3170 44372
rect -9469 44292 -3170 44308
rect -9469 44228 -3254 44292
rect -3190 44228 -3170 44292
rect -9469 44212 -3170 44228
rect -9469 44148 -3254 44212
rect -3190 44148 -3170 44212
rect -9469 44132 -3170 44148
rect -9469 44068 -3254 44132
rect -3190 44068 -3170 44132
rect -9469 44052 -3170 44068
rect -9469 43988 -3254 44052
rect -3190 43988 -3170 44052
rect -9469 43972 -3170 43988
rect -9469 43908 -3254 43972
rect -3190 43908 -3170 43972
rect -9469 43892 -3170 43908
rect -9469 43828 -3254 43892
rect -3190 43828 -3170 43892
rect -9469 43812 -3170 43828
rect -9469 43748 -3254 43812
rect -3190 43748 -3170 43812
rect -9469 43732 -3170 43748
rect -9469 43668 -3254 43732
rect -3190 43668 -3170 43732
rect -9469 43652 -3170 43668
rect -9469 43588 -3254 43652
rect -3190 43588 -3170 43652
rect -9469 43572 -3170 43588
rect -9469 43508 -3254 43572
rect -3190 43508 -3170 43572
rect -9469 43492 -3170 43508
rect -9469 43428 -3254 43492
rect -3190 43428 -3170 43492
rect -9469 43412 -3170 43428
rect -9469 43348 -3254 43412
rect -3190 43348 -3170 43412
rect -9469 43332 -3170 43348
rect -9469 43268 -3254 43332
rect -3190 43268 -3170 43332
rect -9469 43252 -3170 43268
rect -9469 43188 -3254 43252
rect -3190 43188 -3170 43252
rect -9469 43172 -3170 43188
rect -9469 43108 -3254 43172
rect -3190 43108 -3170 43172
rect -9469 43092 -3170 43108
rect -9469 43028 -3254 43092
rect -3190 43028 -3170 43092
rect -9469 43012 -3170 43028
rect -9469 42948 -3254 43012
rect -3190 42948 -3170 43012
rect -9469 42932 -3170 42948
rect -9469 42868 -3254 42932
rect -3190 42868 -3170 42932
rect -9469 42852 -3170 42868
rect -9469 42788 -3254 42852
rect -3190 42788 -3170 42852
rect -9469 42772 -3170 42788
rect -9469 42708 -3254 42772
rect -3190 42708 -3170 42772
rect -9469 42692 -3170 42708
rect -9469 42628 -3254 42692
rect -3190 42628 -3170 42692
rect -9469 42612 -3170 42628
rect -9469 42548 -3254 42612
rect -3190 42548 -3170 42612
rect -9469 42532 -3170 42548
rect -9469 42468 -3254 42532
rect -3190 42468 -3170 42532
rect -9469 42452 -3170 42468
rect -9469 42388 -3254 42452
rect -3190 42388 -3170 42452
rect -9469 42372 -3170 42388
rect -9469 42308 -3254 42372
rect -3190 42308 -3170 42372
rect -9469 42292 -3170 42308
rect -9469 42228 -3254 42292
rect -3190 42228 -3170 42292
rect -9469 42212 -3170 42228
rect -9469 42148 -3254 42212
rect -3190 42148 -3170 42212
rect -9469 42132 -3170 42148
rect -9469 42068 -3254 42132
rect -3190 42068 -3170 42132
rect -9469 42052 -3170 42068
rect -9469 41988 -3254 42052
rect -3190 41988 -3170 42052
rect -9469 41972 -3170 41988
rect -9469 41908 -3254 41972
rect -3190 41908 -3170 41972
rect -9469 41892 -3170 41908
rect -9469 41828 -3254 41892
rect -3190 41828 -3170 41892
rect -9469 41812 -3170 41828
rect -9469 41748 -3254 41812
rect -3190 41748 -3170 41812
rect -9469 41732 -3170 41748
rect -9469 41668 -3254 41732
rect -3190 41668 -3170 41732
rect -9469 41652 -3170 41668
rect -9469 41588 -3254 41652
rect -3190 41588 -3170 41652
rect -9469 41572 -3170 41588
rect -9469 41508 -3254 41572
rect -3190 41508 -3170 41572
rect -9469 41492 -3170 41508
rect -9469 41428 -3254 41492
rect -3190 41428 -3170 41492
rect -9469 41412 -3170 41428
rect -9469 41348 -3254 41412
rect -3190 41348 -3170 41412
rect -9469 41332 -3170 41348
rect -9469 41268 -3254 41332
rect -3190 41268 -3170 41332
rect -9469 41252 -3170 41268
rect -9469 41188 -3254 41252
rect -3190 41188 -3170 41252
rect -9469 41172 -3170 41188
rect -9469 41108 -3254 41172
rect -3190 41108 -3170 41172
rect -9469 41092 -3170 41108
rect -9469 41028 -3254 41092
rect -3190 41028 -3170 41092
rect -9469 41000 -3170 41028
rect -3150 47172 3149 47200
rect -3150 47108 3065 47172
rect 3129 47108 3149 47172
rect -3150 47092 3149 47108
rect -3150 47028 3065 47092
rect 3129 47028 3149 47092
rect -3150 47012 3149 47028
rect -3150 46948 3065 47012
rect 3129 46948 3149 47012
rect -3150 46932 3149 46948
rect -3150 46868 3065 46932
rect 3129 46868 3149 46932
rect -3150 46852 3149 46868
rect -3150 46788 3065 46852
rect 3129 46788 3149 46852
rect -3150 46772 3149 46788
rect -3150 46708 3065 46772
rect 3129 46708 3149 46772
rect -3150 46692 3149 46708
rect -3150 46628 3065 46692
rect 3129 46628 3149 46692
rect -3150 46612 3149 46628
rect -3150 46548 3065 46612
rect 3129 46548 3149 46612
rect -3150 46532 3149 46548
rect -3150 46468 3065 46532
rect 3129 46468 3149 46532
rect -3150 46452 3149 46468
rect -3150 46388 3065 46452
rect 3129 46388 3149 46452
rect -3150 46372 3149 46388
rect -3150 46308 3065 46372
rect 3129 46308 3149 46372
rect -3150 46292 3149 46308
rect -3150 46228 3065 46292
rect 3129 46228 3149 46292
rect -3150 46212 3149 46228
rect -3150 46148 3065 46212
rect 3129 46148 3149 46212
rect -3150 46132 3149 46148
rect -3150 46068 3065 46132
rect 3129 46068 3149 46132
rect -3150 46052 3149 46068
rect -3150 45988 3065 46052
rect 3129 45988 3149 46052
rect -3150 45972 3149 45988
rect -3150 45908 3065 45972
rect 3129 45908 3149 45972
rect -3150 45892 3149 45908
rect -3150 45828 3065 45892
rect 3129 45828 3149 45892
rect -3150 45812 3149 45828
rect -3150 45748 3065 45812
rect 3129 45748 3149 45812
rect -3150 45732 3149 45748
rect -3150 45668 3065 45732
rect 3129 45668 3149 45732
rect -3150 45652 3149 45668
rect -3150 45588 3065 45652
rect 3129 45588 3149 45652
rect -3150 45572 3149 45588
rect -3150 45508 3065 45572
rect 3129 45508 3149 45572
rect -3150 45492 3149 45508
rect -3150 45428 3065 45492
rect 3129 45428 3149 45492
rect -3150 45412 3149 45428
rect -3150 45348 3065 45412
rect 3129 45348 3149 45412
rect -3150 45332 3149 45348
rect -3150 45268 3065 45332
rect 3129 45268 3149 45332
rect -3150 45252 3149 45268
rect -3150 45188 3065 45252
rect 3129 45188 3149 45252
rect -3150 45172 3149 45188
rect -3150 45108 3065 45172
rect 3129 45108 3149 45172
rect -3150 45092 3149 45108
rect -3150 45028 3065 45092
rect 3129 45028 3149 45092
rect -3150 45012 3149 45028
rect -3150 44948 3065 45012
rect 3129 44948 3149 45012
rect -3150 44932 3149 44948
rect -3150 44868 3065 44932
rect 3129 44868 3149 44932
rect -3150 44852 3149 44868
rect -3150 44788 3065 44852
rect 3129 44788 3149 44852
rect -3150 44772 3149 44788
rect -3150 44708 3065 44772
rect 3129 44708 3149 44772
rect -3150 44692 3149 44708
rect -3150 44628 3065 44692
rect 3129 44628 3149 44692
rect -3150 44612 3149 44628
rect -3150 44548 3065 44612
rect 3129 44548 3149 44612
rect -3150 44532 3149 44548
rect -3150 44468 3065 44532
rect 3129 44468 3149 44532
rect -3150 44452 3149 44468
rect -3150 44388 3065 44452
rect 3129 44388 3149 44452
rect -3150 44372 3149 44388
rect -3150 44308 3065 44372
rect 3129 44308 3149 44372
rect -3150 44292 3149 44308
rect -3150 44228 3065 44292
rect 3129 44228 3149 44292
rect -3150 44212 3149 44228
rect -3150 44148 3065 44212
rect 3129 44148 3149 44212
rect -3150 44132 3149 44148
rect -3150 44068 3065 44132
rect 3129 44068 3149 44132
rect -3150 44052 3149 44068
rect -3150 43988 3065 44052
rect 3129 43988 3149 44052
rect -3150 43972 3149 43988
rect -3150 43908 3065 43972
rect 3129 43908 3149 43972
rect -3150 43892 3149 43908
rect -3150 43828 3065 43892
rect 3129 43828 3149 43892
rect -3150 43812 3149 43828
rect -3150 43748 3065 43812
rect 3129 43748 3149 43812
rect -3150 43732 3149 43748
rect -3150 43668 3065 43732
rect 3129 43668 3149 43732
rect -3150 43652 3149 43668
rect -3150 43588 3065 43652
rect 3129 43588 3149 43652
rect -3150 43572 3149 43588
rect -3150 43508 3065 43572
rect 3129 43508 3149 43572
rect -3150 43492 3149 43508
rect -3150 43428 3065 43492
rect 3129 43428 3149 43492
rect -3150 43412 3149 43428
rect -3150 43348 3065 43412
rect 3129 43348 3149 43412
rect -3150 43332 3149 43348
rect -3150 43268 3065 43332
rect 3129 43268 3149 43332
rect -3150 43252 3149 43268
rect -3150 43188 3065 43252
rect 3129 43188 3149 43252
rect -3150 43172 3149 43188
rect -3150 43108 3065 43172
rect 3129 43108 3149 43172
rect -3150 43092 3149 43108
rect -3150 43028 3065 43092
rect 3129 43028 3149 43092
rect -3150 43012 3149 43028
rect -3150 42948 3065 43012
rect 3129 42948 3149 43012
rect -3150 42932 3149 42948
rect -3150 42868 3065 42932
rect 3129 42868 3149 42932
rect -3150 42852 3149 42868
rect -3150 42788 3065 42852
rect 3129 42788 3149 42852
rect -3150 42772 3149 42788
rect -3150 42708 3065 42772
rect 3129 42708 3149 42772
rect -3150 42692 3149 42708
rect -3150 42628 3065 42692
rect 3129 42628 3149 42692
rect -3150 42612 3149 42628
rect -3150 42548 3065 42612
rect 3129 42548 3149 42612
rect -3150 42532 3149 42548
rect -3150 42468 3065 42532
rect 3129 42468 3149 42532
rect -3150 42452 3149 42468
rect -3150 42388 3065 42452
rect 3129 42388 3149 42452
rect -3150 42372 3149 42388
rect -3150 42308 3065 42372
rect 3129 42308 3149 42372
rect -3150 42292 3149 42308
rect -3150 42228 3065 42292
rect 3129 42228 3149 42292
rect -3150 42212 3149 42228
rect -3150 42148 3065 42212
rect 3129 42148 3149 42212
rect -3150 42132 3149 42148
rect -3150 42068 3065 42132
rect 3129 42068 3149 42132
rect -3150 42052 3149 42068
rect -3150 41988 3065 42052
rect 3129 41988 3149 42052
rect -3150 41972 3149 41988
rect -3150 41908 3065 41972
rect 3129 41908 3149 41972
rect -3150 41892 3149 41908
rect -3150 41828 3065 41892
rect 3129 41828 3149 41892
rect -3150 41812 3149 41828
rect -3150 41748 3065 41812
rect 3129 41748 3149 41812
rect -3150 41732 3149 41748
rect -3150 41668 3065 41732
rect 3129 41668 3149 41732
rect -3150 41652 3149 41668
rect -3150 41588 3065 41652
rect 3129 41588 3149 41652
rect -3150 41572 3149 41588
rect -3150 41508 3065 41572
rect 3129 41508 3149 41572
rect -3150 41492 3149 41508
rect -3150 41428 3065 41492
rect 3129 41428 3149 41492
rect -3150 41412 3149 41428
rect -3150 41348 3065 41412
rect 3129 41348 3149 41412
rect -3150 41332 3149 41348
rect -3150 41268 3065 41332
rect 3129 41268 3149 41332
rect -3150 41252 3149 41268
rect -3150 41188 3065 41252
rect 3129 41188 3149 41252
rect -3150 41172 3149 41188
rect -3150 41108 3065 41172
rect 3129 41108 3149 41172
rect -3150 41092 3149 41108
rect -3150 41028 3065 41092
rect 3129 41028 3149 41092
rect -3150 41000 3149 41028
rect 3169 47172 9468 47200
rect 3169 47108 9384 47172
rect 9448 47108 9468 47172
rect 3169 47092 9468 47108
rect 3169 47028 9384 47092
rect 9448 47028 9468 47092
rect 3169 47012 9468 47028
rect 3169 46948 9384 47012
rect 9448 46948 9468 47012
rect 3169 46932 9468 46948
rect 3169 46868 9384 46932
rect 9448 46868 9468 46932
rect 3169 46852 9468 46868
rect 3169 46788 9384 46852
rect 9448 46788 9468 46852
rect 3169 46772 9468 46788
rect 3169 46708 9384 46772
rect 9448 46708 9468 46772
rect 3169 46692 9468 46708
rect 3169 46628 9384 46692
rect 9448 46628 9468 46692
rect 3169 46612 9468 46628
rect 3169 46548 9384 46612
rect 9448 46548 9468 46612
rect 3169 46532 9468 46548
rect 3169 46468 9384 46532
rect 9448 46468 9468 46532
rect 3169 46452 9468 46468
rect 3169 46388 9384 46452
rect 9448 46388 9468 46452
rect 3169 46372 9468 46388
rect 3169 46308 9384 46372
rect 9448 46308 9468 46372
rect 3169 46292 9468 46308
rect 3169 46228 9384 46292
rect 9448 46228 9468 46292
rect 3169 46212 9468 46228
rect 3169 46148 9384 46212
rect 9448 46148 9468 46212
rect 3169 46132 9468 46148
rect 3169 46068 9384 46132
rect 9448 46068 9468 46132
rect 3169 46052 9468 46068
rect 3169 45988 9384 46052
rect 9448 45988 9468 46052
rect 3169 45972 9468 45988
rect 3169 45908 9384 45972
rect 9448 45908 9468 45972
rect 3169 45892 9468 45908
rect 3169 45828 9384 45892
rect 9448 45828 9468 45892
rect 3169 45812 9468 45828
rect 3169 45748 9384 45812
rect 9448 45748 9468 45812
rect 3169 45732 9468 45748
rect 3169 45668 9384 45732
rect 9448 45668 9468 45732
rect 3169 45652 9468 45668
rect 3169 45588 9384 45652
rect 9448 45588 9468 45652
rect 3169 45572 9468 45588
rect 3169 45508 9384 45572
rect 9448 45508 9468 45572
rect 3169 45492 9468 45508
rect 3169 45428 9384 45492
rect 9448 45428 9468 45492
rect 3169 45412 9468 45428
rect 3169 45348 9384 45412
rect 9448 45348 9468 45412
rect 3169 45332 9468 45348
rect 3169 45268 9384 45332
rect 9448 45268 9468 45332
rect 3169 45252 9468 45268
rect 3169 45188 9384 45252
rect 9448 45188 9468 45252
rect 3169 45172 9468 45188
rect 3169 45108 9384 45172
rect 9448 45108 9468 45172
rect 3169 45092 9468 45108
rect 3169 45028 9384 45092
rect 9448 45028 9468 45092
rect 3169 45012 9468 45028
rect 3169 44948 9384 45012
rect 9448 44948 9468 45012
rect 3169 44932 9468 44948
rect 3169 44868 9384 44932
rect 9448 44868 9468 44932
rect 3169 44852 9468 44868
rect 3169 44788 9384 44852
rect 9448 44788 9468 44852
rect 3169 44772 9468 44788
rect 3169 44708 9384 44772
rect 9448 44708 9468 44772
rect 3169 44692 9468 44708
rect 3169 44628 9384 44692
rect 9448 44628 9468 44692
rect 3169 44612 9468 44628
rect 3169 44548 9384 44612
rect 9448 44548 9468 44612
rect 3169 44532 9468 44548
rect 3169 44468 9384 44532
rect 9448 44468 9468 44532
rect 3169 44452 9468 44468
rect 3169 44388 9384 44452
rect 9448 44388 9468 44452
rect 3169 44372 9468 44388
rect 3169 44308 9384 44372
rect 9448 44308 9468 44372
rect 3169 44292 9468 44308
rect 3169 44228 9384 44292
rect 9448 44228 9468 44292
rect 3169 44212 9468 44228
rect 3169 44148 9384 44212
rect 9448 44148 9468 44212
rect 3169 44132 9468 44148
rect 3169 44068 9384 44132
rect 9448 44068 9468 44132
rect 3169 44052 9468 44068
rect 3169 43988 9384 44052
rect 9448 43988 9468 44052
rect 3169 43972 9468 43988
rect 3169 43908 9384 43972
rect 9448 43908 9468 43972
rect 3169 43892 9468 43908
rect 3169 43828 9384 43892
rect 9448 43828 9468 43892
rect 3169 43812 9468 43828
rect 3169 43748 9384 43812
rect 9448 43748 9468 43812
rect 3169 43732 9468 43748
rect 3169 43668 9384 43732
rect 9448 43668 9468 43732
rect 3169 43652 9468 43668
rect 3169 43588 9384 43652
rect 9448 43588 9468 43652
rect 3169 43572 9468 43588
rect 3169 43508 9384 43572
rect 9448 43508 9468 43572
rect 3169 43492 9468 43508
rect 3169 43428 9384 43492
rect 9448 43428 9468 43492
rect 3169 43412 9468 43428
rect 3169 43348 9384 43412
rect 9448 43348 9468 43412
rect 3169 43332 9468 43348
rect 3169 43268 9384 43332
rect 9448 43268 9468 43332
rect 3169 43252 9468 43268
rect 3169 43188 9384 43252
rect 9448 43188 9468 43252
rect 3169 43172 9468 43188
rect 3169 43108 9384 43172
rect 9448 43108 9468 43172
rect 3169 43092 9468 43108
rect 3169 43028 9384 43092
rect 9448 43028 9468 43092
rect 3169 43012 9468 43028
rect 3169 42948 9384 43012
rect 9448 42948 9468 43012
rect 3169 42932 9468 42948
rect 3169 42868 9384 42932
rect 9448 42868 9468 42932
rect 3169 42852 9468 42868
rect 3169 42788 9384 42852
rect 9448 42788 9468 42852
rect 3169 42772 9468 42788
rect 3169 42708 9384 42772
rect 9448 42708 9468 42772
rect 3169 42692 9468 42708
rect 3169 42628 9384 42692
rect 9448 42628 9468 42692
rect 3169 42612 9468 42628
rect 3169 42548 9384 42612
rect 9448 42548 9468 42612
rect 3169 42532 9468 42548
rect 3169 42468 9384 42532
rect 9448 42468 9468 42532
rect 3169 42452 9468 42468
rect 3169 42388 9384 42452
rect 9448 42388 9468 42452
rect 3169 42372 9468 42388
rect 3169 42308 9384 42372
rect 9448 42308 9468 42372
rect 3169 42292 9468 42308
rect 3169 42228 9384 42292
rect 9448 42228 9468 42292
rect 3169 42212 9468 42228
rect 3169 42148 9384 42212
rect 9448 42148 9468 42212
rect 3169 42132 9468 42148
rect 3169 42068 9384 42132
rect 9448 42068 9468 42132
rect 3169 42052 9468 42068
rect 3169 41988 9384 42052
rect 9448 41988 9468 42052
rect 3169 41972 9468 41988
rect 3169 41908 9384 41972
rect 9448 41908 9468 41972
rect 3169 41892 9468 41908
rect 3169 41828 9384 41892
rect 9448 41828 9468 41892
rect 3169 41812 9468 41828
rect 3169 41748 9384 41812
rect 9448 41748 9468 41812
rect 3169 41732 9468 41748
rect 3169 41668 9384 41732
rect 9448 41668 9468 41732
rect 3169 41652 9468 41668
rect 3169 41588 9384 41652
rect 9448 41588 9468 41652
rect 3169 41572 9468 41588
rect 3169 41508 9384 41572
rect 9448 41508 9468 41572
rect 3169 41492 9468 41508
rect 3169 41428 9384 41492
rect 9448 41428 9468 41492
rect 3169 41412 9468 41428
rect 3169 41348 9384 41412
rect 9448 41348 9468 41412
rect 3169 41332 9468 41348
rect 3169 41268 9384 41332
rect 9448 41268 9468 41332
rect 3169 41252 9468 41268
rect 3169 41188 9384 41252
rect 9448 41188 9468 41252
rect 3169 41172 9468 41188
rect 3169 41108 9384 41172
rect 9448 41108 9468 41172
rect 3169 41092 9468 41108
rect 3169 41028 9384 41092
rect 9448 41028 9468 41092
rect 3169 41000 9468 41028
rect 9488 47172 15787 47200
rect 9488 47108 15703 47172
rect 15767 47108 15787 47172
rect 9488 47092 15787 47108
rect 9488 47028 15703 47092
rect 15767 47028 15787 47092
rect 9488 47012 15787 47028
rect 9488 46948 15703 47012
rect 15767 46948 15787 47012
rect 9488 46932 15787 46948
rect 9488 46868 15703 46932
rect 15767 46868 15787 46932
rect 9488 46852 15787 46868
rect 9488 46788 15703 46852
rect 15767 46788 15787 46852
rect 9488 46772 15787 46788
rect 9488 46708 15703 46772
rect 15767 46708 15787 46772
rect 9488 46692 15787 46708
rect 9488 46628 15703 46692
rect 15767 46628 15787 46692
rect 9488 46612 15787 46628
rect 9488 46548 15703 46612
rect 15767 46548 15787 46612
rect 9488 46532 15787 46548
rect 9488 46468 15703 46532
rect 15767 46468 15787 46532
rect 9488 46452 15787 46468
rect 9488 46388 15703 46452
rect 15767 46388 15787 46452
rect 9488 46372 15787 46388
rect 9488 46308 15703 46372
rect 15767 46308 15787 46372
rect 9488 46292 15787 46308
rect 9488 46228 15703 46292
rect 15767 46228 15787 46292
rect 9488 46212 15787 46228
rect 9488 46148 15703 46212
rect 15767 46148 15787 46212
rect 9488 46132 15787 46148
rect 9488 46068 15703 46132
rect 15767 46068 15787 46132
rect 9488 46052 15787 46068
rect 9488 45988 15703 46052
rect 15767 45988 15787 46052
rect 9488 45972 15787 45988
rect 9488 45908 15703 45972
rect 15767 45908 15787 45972
rect 9488 45892 15787 45908
rect 9488 45828 15703 45892
rect 15767 45828 15787 45892
rect 9488 45812 15787 45828
rect 9488 45748 15703 45812
rect 15767 45748 15787 45812
rect 9488 45732 15787 45748
rect 9488 45668 15703 45732
rect 15767 45668 15787 45732
rect 9488 45652 15787 45668
rect 9488 45588 15703 45652
rect 15767 45588 15787 45652
rect 9488 45572 15787 45588
rect 9488 45508 15703 45572
rect 15767 45508 15787 45572
rect 9488 45492 15787 45508
rect 9488 45428 15703 45492
rect 15767 45428 15787 45492
rect 9488 45412 15787 45428
rect 9488 45348 15703 45412
rect 15767 45348 15787 45412
rect 9488 45332 15787 45348
rect 9488 45268 15703 45332
rect 15767 45268 15787 45332
rect 9488 45252 15787 45268
rect 9488 45188 15703 45252
rect 15767 45188 15787 45252
rect 9488 45172 15787 45188
rect 9488 45108 15703 45172
rect 15767 45108 15787 45172
rect 9488 45092 15787 45108
rect 9488 45028 15703 45092
rect 15767 45028 15787 45092
rect 9488 45012 15787 45028
rect 9488 44948 15703 45012
rect 15767 44948 15787 45012
rect 9488 44932 15787 44948
rect 9488 44868 15703 44932
rect 15767 44868 15787 44932
rect 9488 44852 15787 44868
rect 9488 44788 15703 44852
rect 15767 44788 15787 44852
rect 9488 44772 15787 44788
rect 9488 44708 15703 44772
rect 15767 44708 15787 44772
rect 9488 44692 15787 44708
rect 9488 44628 15703 44692
rect 15767 44628 15787 44692
rect 9488 44612 15787 44628
rect 9488 44548 15703 44612
rect 15767 44548 15787 44612
rect 9488 44532 15787 44548
rect 9488 44468 15703 44532
rect 15767 44468 15787 44532
rect 9488 44452 15787 44468
rect 9488 44388 15703 44452
rect 15767 44388 15787 44452
rect 9488 44372 15787 44388
rect 9488 44308 15703 44372
rect 15767 44308 15787 44372
rect 9488 44292 15787 44308
rect 9488 44228 15703 44292
rect 15767 44228 15787 44292
rect 9488 44212 15787 44228
rect 9488 44148 15703 44212
rect 15767 44148 15787 44212
rect 9488 44132 15787 44148
rect 9488 44068 15703 44132
rect 15767 44068 15787 44132
rect 9488 44052 15787 44068
rect 9488 43988 15703 44052
rect 15767 43988 15787 44052
rect 9488 43972 15787 43988
rect 9488 43908 15703 43972
rect 15767 43908 15787 43972
rect 9488 43892 15787 43908
rect 9488 43828 15703 43892
rect 15767 43828 15787 43892
rect 9488 43812 15787 43828
rect 9488 43748 15703 43812
rect 15767 43748 15787 43812
rect 9488 43732 15787 43748
rect 9488 43668 15703 43732
rect 15767 43668 15787 43732
rect 9488 43652 15787 43668
rect 9488 43588 15703 43652
rect 15767 43588 15787 43652
rect 9488 43572 15787 43588
rect 9488 43508 15703 43572
rect 15767 43508 15787 43572
rect 9488 43492 15787 43508
rect 9488 43428 15703 43492
rect 15767 43428 15787 43492
rect 9488 43412 15787 43428
rect 9488 43348 15703 43412
rect 15767 43348 15787 43412
rect 9488 43332 15787 43348
rect 9488 43268 15703 43332
rect 15767 43268 15787 43332
rect 9488 43252 15787 43268
rect 9488 43188 15703 43252
rect 15767 43188 15787 43252
rect 9488 43172 15787 43188
rect 9488 43108 15703 43172
rect 15767 43108 15787 43172
rect 9488 43092 15787 43108
rect 9488 43028 15703 43092
rect 15767 43028 15787 43092
rect 9488 43012 15787 43028
rect 9488 42948 15703 43012
rect 15767 42948 15787 43012
rect 9488 42932 15787 42948
rect 9488 42868 15703 42932
rect 15767 42868 15787 42932
rect 9488 42852 15787 42868
rect 9488 42788 15703 42852
rect 15767 42788 15787 42852
rect 9488 42772 15787 42788
rect 9488 42708 15703 42772
rect 15767 42708 15787 42772
rect 9488 42692 15787 42708
rect 9488 42628 15703 42692
rect 15767 42628 15787 42692
rect 9488 42612 15787 42628
rect 9488 42548 15703 42612
rect 15767 42548 15787 42612
rect 9488 42532 15787 42548
rect 9488 42468 15703 42532
rect 15767 42468 15787 42532
rect 9488 42452 15787 42468
rect 9488 42388 15703 42452
rect 15767 42388 15787 42452
rect 9488 42372 15787 42388
rect 9488 42308 15703 42372
rect 15767 42308 15787 42372
rect 9488 42292 15787 42308
rect 9488 42228 15703 42292
rect 15767 42228 15787 42292
rect 9488 42212 15787 42228
rect 9488 42148 15703 42212
rect 15767 42148 15787 42212
rect 9488 42132 15787 42148
rect 9488 42068 15703 42132
rect 15767 42068 15787 42132
rect 9488 42052 15787 42068
rect 9488 41988 15703 42052
rect 15767 41988 15787 42052
rect 9488 41972 15787 41988
rect 9488 41908 15703 41972
rect 15767 41908 15787 41972
rect 9488 41892 15787 41908
rect 9488 41828 15703 41892
rect 15767 41828 15787 41892
rect 9488 41812 15787 41828
rect 9488 41748 15703 41812
rect 15767 41748 15787 41812
rect 9488 41732 15787 41748
rect 9488 41668 15703 41732
rect 15767 41668 15787 41732
rect 9488 41652 15787 41668
rect 9488 41588 15703 41652
rect 15767 41588 15787 41652
rect 9488 41572 15787 41588
rect 9488 41508 15703 41572
rect 15767 41508 15787 41572
rect 9488 41492 15787 41508
rect 9488 41428 15703 41492
rect 15767 41428 15787 41492
rect 9488 41412 15787 41428
rect 9488 41348 15703 41412
rect 15767 41348 15787 41412
rect 9488 41332 15787 41348
rect 9488 41268 15703 41332
rect 15767 41268 15787 41332
rect 9488 41252 15787 41268
rect 9488 41188 15703 41252
rect 15767 41188 15787 41252
rect 9488 41172 15787 41188
rect 9488 41108 15703 41172
rect 15767 41108 15787 41172
rect 9488 41092 15787 41108
rect 9488 41028 15703 41092
rect 15767 41028 15787 41092
rect 9488 41000 15787 41028
rect 15807 47172 22106 47200
rect 15807 47108 22022 47172
rect 22086 47108 22106 47172
rect 15807 47092 22106 47108
rect 15807 47028 22022 47092
rect 22086 47028 22106 47092
rect 15807 47012 22106 47028
rect 15807 46948 22022 47012
rect 22086 46948 22106 47012
rect 15807 46932 22106 46948
rect 15807 46868 22022 46932
rect 22086 46868 22106 46932
rect 15807 46852 22106 46868
rect 15807 46788 22022 46852
rect 22086 46788 22106 46852
rect 15807 46772 22106 46788
rect 15807 46708 22022 46772
rect 22086 46708 22106 46772
rect 15807 46692 22106 46708
rect 15807 46628 22022 46692
rect 22086 46628 22106 46692
rect 15807 46612 22106 46628
rect 15807 46548 22022 46612
rect 22086 46548 22106 46612
rect 15807 46532 22106 46548
rect 15807 46468 22022 46532
rect 22086 46468 22106 46532
rect 15807 46452 22106 46468
rect 15807 46388 22022 46452
rect 22086 46388 22106 46452
rect 15807 46372 22106 46388
rect 15807 46308 22022 46372
rect 22086 46308 22106 46372
rect 15807 46292 22106 46308
rect 15807 46228 22022 46292
rect 22086 46228 22106 46292
rect 15807 46212 22106 46228
rect 15807 46148 22022 46212
rect 22086 46148 22106 46212
rect 15807 46132 22106 46148
rect 15807 46068 22022 46132
rect 22086 46068 22106 46132
rect 15807 46052 22106 46068
rect 15807 45988 22022 46052
rect 22086 45988 22106 46052
rect 15807 45972 22106 45988
rect 15807 45908 22022 45972
rect 22086 45908 22106 45972
rect 15807 45892 22106 45908
rect 15807 45828 22022 45892
rect 22086 45828 22106 45892
rect 15807 45812 22106 45828
rect 15807 45748 22022 45812
rect 22086 45748 22106 45812
rect 15807 45732 22106 45748
rect 15807 45668 22022 45732
rect 22086 45668 22106 45732
rect 15807 45652 22106 45668
rect 15807 45588 22022 45652
rect 22086 45588 22106 45652
rect 15807 45572 22106 45588
rect 15807 45508 22022 45572
rect 22086 45508 22106 45572
rect 15807 45492 22106 45508
rect 15807 45428 22022 45492
rect 22086 45428 22106 45492
rect 15807 45412 22106 45428
rect 15807 45348 22022 45412
rect 22086 45348 22106 45412
rect 15807 45332 22106 45348
rect 15807 45268 22022 45332
rect 22086 45268 22106 45332
rect 15807 45252 22106 45268
rect 15807 45188 22022 45252
rect 22086 45188 22106 45252
rect 15807 45172 22106 45188
rect 15807 45108 22022 45172
rect 22086 45108 22106 45172
rect 15807 45092 22106 45108
rect 15807 45028 22022 45092
rect 22086 45028 22106 45092
rect 15807 45012 22106 45028
rect 15807 44948 22022 45012
rect 22086 44948 22106 45012
rect 15807 44932 22106 44948
rect 15807 44868 22022 44932
rect 22086 44868 22106 44932
rect 15807 44852 22106 44868
rect 15807 44788 22022 44852
rect 22086 44788 22106 44852
rect 15807 44772 22106 44788
rect 15807 44708 22022 44772
rect 22086 44708 22106 44772
rect 15807 44692 22106 44708
rect 15807 44628 22022 44692
rect 22086 44628 22106 44692
rect 15807 44612 22106 44628
rect 15807 44548 22022 44612
rect 22086 44548 22106 44612
rect 15807 44532 22106 44548
rect 15807 44468 22022 44532
rect 22086 44468 22106 44532
rect 15807 44452 22106 44468
rect 15807 44388 22022 44452
rect 22086 44388 22106 44452
rect 15807 44372 22106 44388
rect 15807 44308 22022 44372
rect 22086 44308 22106 44372
rect 15807 44292 22106 44308
rect 15807 44228 22022 44292
rect 22086 44228 22106 44292
rect 15807 44212 22106 44228
rect 15807 44148 22022 44212
rect 22086 44148 22106 44212
rect 15807 44132 22106 44148
rect 15807 44068 22022 44132
rect 22086 44068 22106 44132
rect 15807 44052 22106 44068
rect 15807 43988 22022 44052
rect 22086 43988 22106 44052
rect 15807 43972 22106 43988
rect 15807 43908 22022 43972
rect 22086 43908 22106 43972
rect 15807 43892 22106 43908
rect 15807 43828 22022 43892
rect 22086 43828 22106 43892
rect 15807 43812 22106 43828
rect 15807 43748 22022 43812
rect 22086 43748 22106 43812
rect 15807 43732 22106 43748
rect 15807 43668 22022 43732
rect 22086 43668 22106 43732
rect 15807 43652 22106 43668
rect 15807 43588 22022 43652
rect 22086 43588 22106 43652
rect 15807 43572 22106 43588
rect 15807 43508 22022 43572
rect 22086 43508 22106 43572
rect 15807 43492 22106 43508
rect 15807 43428 22022 43492
rect 22086 43428 22106 43492
rect 15807 43412 22106 43428
rect 15807 43348 22022 43412
rect 22086 43348 22106 43412
rect 15807 43332 22106 43348
rect 15807 43268 22022 43332
rect 22086 43268 22106 43332
rect 15807 43252 22106 43268
rect 15807 43188 22022 43252
rect 22086 43188 22106 43252
rect 15807 43172 22106 43188
rect 15807 43108 22022 43172
rect 22086 43108 22106 43172
rect 15807 43092 22106 43108
rect 15807 43028 22022 43092
rect 22086 43028 22106 43092
rect 15807 43012 22106 43028
rect 15807 42948 22022 43012
rect 22086 42948 22106 43012
rect 15807 42932 22106 42948
rect 15807 42868 22022 42932
rect 22086 42868 22106 42932
rect 15807 42852 22106 42868
rect 15807 42788 22022 42852
rect 22086 42788 22106 42852
rect 15807 42772 22106 42788
rect 15807 42708 22022 42772
rect 22086 42708 22106 42772
rect 15807 42692 22106 42708
rect 15807 42628 22022 42692
rect 22086 42628 22106 42692
rect 15807 42612 22106 42628
rect 15807 42548 22022 42612
rect 22086 42548 22106 42612
rect 15807 42532 22106 42548
rect 15807 42468 22022 42532
rect 22086 42468 22106 42532
rect 15807 42452 22106 42468
rect 15807 42388 22022 42452
rect 22086 42388 22106 42452
rect 15807 42372 22106 42388
rect 15807 42308 22022 42372
rect 22086 42308 22106 42372
rect 15807 42292 22106 42308
rect 15807 42228 22022 42292
rect 22086 42228 22106 42292
rect 15807 42212 22106 42228
rect 15807 42148 22022 42212
rect 22086 42148 22106 42212
rect 15807 42132 22106 42148
rect 15807 42068 22022 42132
rect 22086 42068 22106 42132
rect 15807 42052 22106 42068
rect 15807 41988 22022 42052
rect 22086 41988 22106 42052
rect 15807 41972 22106 41988
rect 15807 41908 22022 41972
rect 22086 41908 22106 41972
rect 15807 41892 22106 41908
rect 15807 41828 22022 41892
rect 22086 41828 22106 41892
rect 15807 41812 22106 41828
rect 15807 41748 22022 41812
rect 22086 41748 22106 41812
rect 15807 41732 22106 41748
rect 15807 41668 22022 41732
rect 22086 41668 22106 41732
rect 15807 41652 22106 41668
rect 15807 41588 22022 41652
rect 22086 41588 22106 41652
rect 15807 41572 22106 41588
rect 15807 41508 22022 41572
rect 22086 41508 22106 41572
rect 15807 41492 22106 41508
rect 15807 41428 22022 41492
rect 22086 41428 22106 41492
rect 15807 41412 22106 41428
rect 15807 41348 22022 41412
rect 22086 41348 22106 41412
rect 15807 41332 22106 41348
rect 15807 41268 22022 41332
rect 22086 41268 22106 41332
rect 15807 41252 22106 41268
rect 15807 41188 22022 41252
rect 22086 41188 22106 41252
rect 15807 41172 22106 41188
rect 15807 41108 22022 41172
rect 22086 41108 22106 41172
rect 15807 41092 22106 41108
rect 15807 41028 22022 41092
rect 22086 41028 22106 41092
rect 15807 41000 22106 41028
rect 22126 47172 28425 47200
rect 22126 47108 28341 47172
rect 28405 47108 28425 47172
rect 22126 47092 28425 47108
rect 22126 47028 28341 47092
rect 28405 47028 28425 47092
rect 22126 47012 28425 47028
rect 22126 46948 28341 47012
rect 28405 46948 28425 47012
rect 22126 46932 28425 46948
rect 22126 46868 28341 46932
rect 28405 46868 28425 46932
rect 22126 46852 28425 46868
rect 22126 46788 28341 46852
rect 28405 46788 28425 46852
rect 22126 46772 28425 46788
rect 22126 46708 28341 46772
rect 28405 46708 28425 46772
rect 22126 46692 28425 46708
rect 22126 46628 28341 46692
rect 28405 46628 28425 46692
rect 22126 46612 28425 46628
rect 22126 46548 28341 46612
rect 28405 46548 28425 46612
rect 22126 46532 28425 46548
rect 22126 46468 28341 46532
rect 28405 46468 28425 46532
rect 22126 46452 28425 46468
rect 22126 46388 28341 46452
rect 28405 46388 28425 46452
rect 22126 46372 28425 46388
rect 22126 46308 28341 46372
rect 28405 46308 28425 46372
rect 22126 46292 28425 46308
rect 22126 46228 28341 46292
rect 28405 46228 28425 46292
rect 22126 46212 28425 46228
rect 22126 46148 28341 46212
rect 28405 46148 28425 46212
rect 22126 46132 28425 46148
rect 22126 46068 28341 46132
rect 28405 46068 28425 46132
rect 22126 46052 28425 46068
rect 22126 45988 28341 46052
rect 28405 45988 28425 46052
rect 22126 45972 28425 45988
rect 22126 45908 28341 45972
rect 28405 45908 28425 45972
rect 22126 45892 28425 45908
rect 22126 45828 28341 45892
rect 28405 45828 28425 45892
rect 22126 45812 28425 45828
rect 22126 45748 28341 45812
rect 28405 45748 28425 45812
rect 22126 45732 28425 45748
rect 22126 45668 28341 45732
rect 28405 45668 28425 45732
rect 22126 45652 28425 45668
rect 22126 45588 28341 45652
rect 28405 45588 28425 45652
rect 22126 45572 28425 45588
rect 22126 45508 28341 45572
rect 28405 45508 28425 45572
rect 22126 45492 28425 45508
rect 22126 45428 28341 45492
rect 28405 45428 28425 45492
rect 22126 45412 28425 45428
rect 22126 45348 28341 45412
rect 28405 45348 28425 45412
rect 22126 45332 28425 45348
rect 22126 45268 28341 45332
rect 28405 45268 28425 45332
rect 22126 45252 28425 45268
rect 22126 45188 28341 45252
rect 28405 45188 28425 45252
rect 22126 45172 28425 45188
rect 22126 45108 28341 45172
rect 28405 45108 28425 45172
rect 22126 45092 28425 45108
rect 22126 45028 28341 45092
rect 28405 45028 28425 45092
rect 22126 45012 28425 45028
rect 22126 44948 28341 45012
rect 28405 44948 28425 45012
rect 22126 44932 28425 44948
rect 22126 44868 28341 44932
rect 28405 44868 28425 44932
rect 22126 44852 28425 44868
rect 22126 44788 28341 44852
rect 28405 44788 28425 44852
rect 22126 44772 28425 44788
rect 22126 44708 28341 44772
rect 28405 44708 28425 44772
rect 22126 44692 28425 44708
rect 22126 44628 28341 44692
rect 28405 44628 28425 44692
rect 22126 44612 28425 44628
rect 22126 44548 28341 44612
rect 28405 44548 28425 44612
rect 22126 44532 28425 44548
rect 22126 44468 28341 44532
rect 28405 44468 28425 44532
rect 22126 44452 28425 44468
rect 22126 44388 28341 44452
rect 28405 44388 28425 44452
rect 22126 44372 28425 44388
rect 22126 44308 28341 44372
rect 28405 44308 28425 44372
rect 22126 44292 28425 44308
rect 22126 44228 28341 44292
rect 28405 44228 28425 44292
rect 22126 44212 28425 44228
rect 22126 44148 28341 44212
rect 28405 44148 28425 44212
rect 22126 44132 28425 44148
rect 22126 44068 28341 44132
rect 28405 44068 28425 44132
rect 22126 44052 28425 44068
rect 22126 43988 28341 44052
rect 28405 43988 28425 44052
rect 22126 43972 28425 43988
rect 22126 43908 28341 43972
rect 28405 43908 28425 43972
rect 22126 43892 28425 43908
rect 22126 43828 28341 43892
rect 28405 43828 28425 43892
rect 22126 43812 28425 43828
rect 22126 43748 28341 43812
rect 28405 43748 28425 43812
rect 22126 43732 28425 43748
rect 22126 43668 28341 43732
rect 28405 43668 28425 43732
rect 22126 43652 28425 43668
rect 22126 43588 28341 43652
rect 28405 43588 28425 43652
rect 22126 43572 28425 43588
rect 22126 43508 28341 43572
rect 28405 43508 28425 43572
rect 22126 43492 28425 43508
rect 22126 43428 28341 43492
rect 28405 43428 28425 43492
rect 22126 43412 28425 43428
rect 22126 43348 28341 43412
rect 28405 43348 28425 43412
rect 22126 43332 28425 43348
rect 22126 43268 28341 43332
rect 28405 43268 28425 43332
rect 22126 43252 28425 43268
rect 22126 43188 28341 43252
rect 28405 43188 28425 43252
rect 22126 43172 28425 43188
rect 22126 43108 28341 43172
rect 28405 43108 28425 43172
rect 22126 43092 28425 43108
rect 22126 43028 28341 43092
rect 28405 43028 28425 43092
rect 22126 43012 28425 43028
rect 22126 42948 28341 43012
rect 28405 42948 28425 43012
rect 22126 42932 28425 42948
rect 22126 42868 28341 42932
rect 28405 42868 28425 42932
rect 22126 42852 28425 42868
rect 22126 42788 28341 42852
rect 28405 42788 28425 42852
rect 22126 42772 28425 42788
rect 22126 42708 28341 42772
rect 28405 42708 28425 42772
rect 22126 42692 28425 42708
rect 22126 42628 28341 42692
rect 28405 42628 28425 42692
rect 22126 42612 28425 42628
rect 22126 42548 28341 42612
rect 28405 42548 28425 42612
rect 22126 42532 28425 42548
rect 22126 42468 28341 42532
rect 28405 42468 28425 42532
rect 22126 42452 28425 42468
rect 22126 42388 28341 42452
rect 28405 42388 28425 42452
rect 22126 42372 28425 42388
rect 22126 42308 28341 42372
rect 28405 42308 28425 42372
rect 22126 42292 28425 42308
rect 22126 42228 28341 42292
rect 28405 42228 28425 42292
rect 22126 42212 28425 42228
rect 22126 42148 28341 42212
rect 28405 42148 28425 42212
rect 22126 42132 28425 42148
rect 22126 42068 28341 42132
rect 28405 42068 28425 42132
rect 22126 42052 28425 42068
rect 22126 41988 28341 42052
rect 28405 41988 28425 42052
rect 22126 41972 28425 41988
rect 22126 41908 28341 41972
rect 28405 41908 28425 41972
rect 22126 41892 28425 41908
rect 22126 41828 28341 41892
rect 28405 41828 28425 41892
rect 22126 41812 28425 41828
rect 22126 41748 28341 41812
rect 28405 41748 28425 41812
rect 22126 41732 28425 41748
rect 22126 41668 28341 41732
rect 28405 41668 28425 41732
rect 22126 41652 28425 41668
rect 22126 41588 28341 41652
rect 28405 41588 28425 41652
rect 22126 41572 28425 41588
rect 22126 41508 28341 41572
rect 28405 41508 28425 41572
rect 22126 41492 28425 41508
rect 22126 41428 28341 41492
rect 28405 41428 28425 41492
rect 22126 41412 28425 41428
rect 22126 41348 28341 41412
rect 28405 41348 28425 41412
rect 22126 41332 28425 41348
rect 22126 41268 28341 41332
rect 28405 41268 28425 41332
rect 22126 41252 28425 41268
rect 22126 41188 28341 41252
rect 28405 41188 28425 41252
rect 22126 41172 28425 41188
rect 22126 41108 28341 41172
rect 28405 41108 28425 41172
rect 22126 41092 28425 41108
rect 22126 41028 28341 41092
rect 28405 41028 28425 41092
rect 22126 41000 28425 41028
rect 28445 47172 34744 47200
rect 28445 47108 34660 47172
rect 34724 47108 34744 47172
rect 28445 47092 34744 47108
rect 28445 47028 34660 47092
rect 34724 47028 34744 47092
rect 28445 47012 34744 47028
rect 28445 46948 34660 47012
rect 34724 46948 34744 47012
rect 28445 46932 34744 46948
rect 28445 46868 34660 46932
rect 34724 46868 34744 46932
rect 28445 46852 34744 46868
rect 28445 46788 34660 46852
rect 34724 46788 34744 46852
rect 28445 46772 34744 46788
rect 28445 46708 34660 46772
rect 34724 46708 34744 46772
rect 28445 46692 34744 46708
rect 28445 46628 34660 46692
rect 34724 46628 34744 46692
rect 28445 46612 34744 46628
rect 28445 46548 34660 46612
rect 34724 46548 34744 46612
rect 28445 46532 34744 46548
rect 28445 46468 34660 46532
rect 34724 46468 34744 46532
rect 28445 46452 34744 46468
rect 28445 46388 34660 46452
rect 34724 46388 34744 46452
rect 28445 46372 34744 46388
rect 28445 46308 34660 46372
rect 34724 46308 34744 46372
rect 28445 46292 34744 46308
rect 28445 46228 34660 46292
rect 34724 46228 34744 46292
rect 28445 46212 34744 46228
rect 28445 46148 34660 46212
rect 34724 46148 34744 46212
rect 28445 46132 34744 46148
rect 28445 46068 34660 46132
rect 34724 46068 34744 46132
rect 28445 46052 34744 46068
rect 28445 45988 34660 46052
rect 34724 45988 34744 46052
rect 28445 45972 34744 45988
rect 28445 45908 34660 45972
rect 34724 45908 34744 45972
rect 28445 45892 34744 45908
rect 28445 45828 34660 45892
rect 34724 45828 34744 45892
rect 28445 45812 34744 45828
rect 28445 45748 34660 45812
rect 34724 45748 34744 45812
rect 28445 45732 34744 45748
rect 28445 45668 34660 45732
rect 34724 45668 34744 45732
rect 28445 45652 34744 45668
rect 28445 45588 34660 45652
rect 34724 45588 34744 45652
rect 28445 45572 34744 45588
rect 28445 45508 34660 45572
rect 34724 45508 34744 45572
rect 28445 45492 34744 45508
rect 28445 45428 34660 45492
rect 34724 45428 34744 45492
rect 28445 45412 34744 45428
rect 28445 45348 34660 45412
rect 34724 45348 34744 45412
rect 28445 45332 34744 45348
rect 28445 45268 34660 45332
rect 34724 45268 34744 45332
rect 28445 45252 34744 45268
rect 28445 45188 34660 45252
rect 34724 45188 34744 45252
rect 28445 45172 34744 45188
rect 28445 45108 34660 45172
rect 34724 45108 34744 45172
rect 28445 45092 34744 45108
rect 28445 45028 34660 45092
rect 34724 45028 34744 45092
rect 28445 45012 34744 45028
rect 28445 44948 34660 45012
rect 34724 44948 34744 45012
rect 28445 44932 34744 44948
rect 28445 44868 34660 44932
rect 34724 44868 34744 44932
rect 28445 44852 34744 44868
rect 28445 44788 34660 44852
rect 34724 44788 34744 44852
rect 28445 44772 34744 44788
rect 28445 44708 34660 44772
rect 34724 44708 34744 44772
rect 28445 44692 34744 44708
rect 28445 44628 34660 44692
rect 34724 44628 34744 44692
rect 28445 44612 34744 44628
rect 28445 44548 34660 44612
rect 34724 44548 34744 44612
rect 28445 44532 34744 44548
rect 28445 44468 34660 44532
rect 34724 44468 34744 44532
rect 28445 44452 34744 44468
rect 28445 44388 34660 44452
rect 34724 44388 34744 44452
rect 28445 44372 34744 44388
rect 28445 44308 34660 44372
rect 34724 44308 34744 44372
rect 28445 44292 34744 44308
rect 28445 44228 34660 44292
rect 34724 44228 34744 44292
rect 28445 44212 34744 44228
rect 28445 44148 34660 44212
rect 34724 44148 34744 44212
rect 28445 44132 34744 44148
rect 28445 44068 34660 44132
rect 34724 44068 34744 44132
rect 28445 44052 34744 44068
rect 28445 43988 34660 44052
rect 34724 43988 34744 44052
rect 28445 43972 34744 43988
rect 28445 43908 34660 43972
rect 34724 43908 34744 43972
rect 28445 43892 34744 43908
rect 28445 43828 34660 43892
rect 34724 43828 34744 43892
rect 28445 43812 34744 43828
rect 28445 43748 34660 43812
rect 34724 43748 34744 43812
rect 28445 43732 34744 43748
rect 28445 43668 34660 43732
rect 34724 43668 34744 43732
rect 28445 43652 34744 43668
rect 28445 43588 34660 43652
rect 34724 43588 34744 43652
rect 28445 43572 34744 43588
rect 28445 43508 34660 43572
rect 34724 43508 34744 43572
rect 28445 43492 34744 43508
rect 28445 43428 34660 43492
rect 34724 43428 34744 43492
rect 28445 43412 34744 43428
rect 28445 43348 34660 43412
rect 34724 43348 34744 43412
rect 28445 43332 34744 43348
rect 28445 43268 34660 43332
rect 34724 43268 34744 43332
rect 28445 43252 34744 43268
rect 28445 43188 34660 43252
rect 34724 43188 34744 43252
rect 28445 43172 34744 43188
rect 28445 43108 34660 43172
rect 34724 43108 34744 43172
rect 28445 43092 34744 43108
rect 28445 43028 34660 43092
rect 34724 43028 34744 43092
rect 28445 43012 34744 43028
rect 28445 42948 34660 43012
rect 34724 42948 34744 43012
rect 28445 42932 34744 42948
rect 28445 42868 34660 42932
rect 34724 42868 34744 42932
rect 28445 42852 34744 42868
rect 28445 42788 34660 42852
rect 34724 42788 34744 42852
rect 28445 42772 34744 42788
rect 28445 42708 34660 42772
rect 34724 42708 34744 42772
rect 28445 42692 34744 42708
rect 28445 42628 34660 42692
rect 34724 42628 34744 42692
rect 28445 42612 34744 42628
rect 28445 42548 34660 42612
rect 34724 42548 34744 42612
rect 28445 42532 34744 42548
rect 28445 42468 34660 42532
rect 34724 42468 34744 42532
rect 28445 42452 34744 42468
rect 28445 42388 34660 42452
rect 34724 42388 34744 42452
rect 28445 42372 34744 42388
rect 28445 42308 34660 42372
rect 34724 42308 34744 42372
rect 28445 42292 34744 42308
rect 28445 42228 34660 42292
rect 34724 42228 34744 42292
rect 28445 42212 34744 42228
rect 28445 42148 34660 42212
rect 34724 42148 34744 42212
rect 28445 42132 34744 42148
rect 28445 42068 34660 42132
rect 34724 42068 34744 42132
rect 28445 42052 34744 42068
rect 28445 41988 34660 42052
rect 34724 41988 34744 42052
rect 28445 41972 34744 41988
rect 28445 41908 34660 41972
rect 34724 41908 34744 41972
rect 28445 41892 34744 41908
rect 28445 41828 34660 41892
rect 34724 41828 34744 41892
rect 28445 41812 34744 41828
rect 28445 41748 34660 41812
rect 34724 41748 34744 41812
rect 28445 41732 34744 41748
rect 28445 41668 34660 41732
rect 34724 41668 34744 41732
rect 28445 41652 34744 41668
rect 28445 41588 34660 41652
rect 34724 41588 34744 41652
rect 28445 41572 34744 41588
rect 28445 41508 34660 41572
rect 34724 41508 34744 41572
rect 28445 41492 34744 41508
rect 28445 41428 34660 41492
rect 34724 41428 34744 41492
rect 28445 41412 34744 41428
rect 28445 41348 34660 41412
rect 34724 41348 34744 41412
rect 28445 41332 34744 41348
rect 28445 41268 34660 41332
rect 34724 41268 34744 41332
rect 28445 41252 34744 41268
rect 28445 41188 34660 41252
rect 34724 41188 34744 41252
rect 28445 41172 34744 41188
rect 28445 41108 34660 41172
rect 34724 41108 34744 41172
rect 28445 41092 34744 41108
rect 28445 41028 34660 41092
rect 34724 41028 34744 41092
rect 28445 41000 34744 41028
rect 34764 47172 41063 47200
rect 34764 47108 40979 47172
rect 41043 47108 41063 47172
rect 34764 47092 41063 47108
rect 34764 47028 40979 47092
rect 41043 47028 41063 47092
rect 34764 47012 41063 47028
rect 34764 46948 40979 47012
rect 41043 46948 41063 47012
rect 34764 46932 41063 46948
rect 34764 46868 40979 46932
rect 41043 46868 41063 46932
rect 34764 46852 41063 46868
rect 34764 46788 40979 46852
rect 41043 46788 41063 46852
rect 34764 46772 41063 46788
rect 34764 46708 40979 46772
rect 41043 46708 41063 46772
rect 34764 46692 41063 46708
rect 34764 46628 40979 46692
rect 41043 46628 41063 46692
rect 34764 46612 41063 46628
rect 34764 46548 40979 46612
rect 41043 46548 41063 46612
rect 34764 46532 41063 46548
rect 34764 46468 40979 46532
rect 41043 46468 41063 46532
rect 34764 46452 41063 46468
rect 34764 46388 40979 46452
rect 41043 46388 41063 46452
rect 34764 46372 41063 46388
rect 34764 46308 40979 46372
rect 41043 46308 41063 46372
rect 34764 46292 41063 46308
rect 34764 46228 40979 46292
rect 41043 46228 41063 46292
rect 34764 46212 41063 46228
rect 34764 46148 40979 46212
rect 41043 46148 41063 46212
rect 34764 46132 41063 46148
rect 34764 46068 40979 46132
rect 41043 46068 41063 46132
rect 34764 46052 41063 46068
rect 34764 45988 40979 46052
rect 41043 45988 41063 46052
rect 34764 45972 41063 45988
rect 34764 45908 40979 45972
rect 41043 45908 41063 45972
rect 34764 45892 41063 45908
rect 34764 45828 40979 45892
rect 41043 45828 41063 45892
rect 34764 45812 41063 45828
rect 34764 45748 40979 45812
rect 41043 45748 41063 45812
rect 34764 45732 41063 45748
rect 34764 45668 40979 45732
rect 41043 45668 41063 45732
rect 34764 45652 41063 45668
rect 34764 45588 40979 45652
rect 41043 45588 41063 45652
rect 34764 45572 41063 45588
rect 34764 45508 40979 45572
rect 41043 45508 41063 45572
rect 34764 45492 41063 45508
rect 34764 45428 40979 45492
rect 41043 45428 41063 45492
rect 34764 45412 41063 45428
rect 34764 45348 40979 45412
rect 41043 45348 41063 45412
rect 34764 45332 41063 45348
rect 34764 45268 40979 45332
rect 41043 45268 41063 45332
rect 34764 45252 41063 45268
rect 34764 45188 40979 45252
rect 41043 45188 41063 45252
rect 34764 45172 41063 45188
rect 34764 45108 40979 45172
rect 41043 45108 41063 45172
rect 34764 45092 41063 45108
rect 34764 45028 40979 45092
rect 41043 45028 41063 45092
rect 34764 45012 41063 45028
rect 34764 44948 40979 45012
rect 41043 44948 41063 45012
rect 34764 44932 41063 44948
rect 34764 44868 40979 44932
rect 41043 44868 41063 44932
rect 34764 44852 41063 44868
rect 34764 44788 40979 44852
rect 41043 44788 41063 44852
rect 34764 44772 41063 44788
rect 34764 44708 40979 44772
rect 41043 44708 41063 44772
rect 34764 44692 41063 44708
rect 34764 44628 40979 44692
rect 41043 44628 41063 44692
rect 34764 44612 41063 44628
rect 34764 44548 40979 44612
rect 41043 44548 41063 44612
rect 34764 44532 41063 44548
rect 34764 44468 40979 44532
rect 41043 44468 41063 44532
rect 34764 44452 41063 44468
rect 34764 44388 40979 44452
rect 41043 44388 41063 44452
rect 34764 44372 41063 44388
rect 34764 44308 40979 44372
rect 41043 44308 41063 44372
rect 34764 44292 41063 44308
rect 34764 44228 40979 44292
rect 41043 44228 41063 44292
rect 34764 44212 41063 44228
rect 34764 44148 40979 44212
rect 41043 44148 41063 44212
rect 34764 44132 41063 44148
rect 34764 44068 40979 44132
rect 41043 44068 41063 44132
rect 34764 44052 41063 44068
rect 34764 43988 40979 44052
rect 41043 43988 41063 44052
rect 34764 43972 41063 43988
rect 34764 43908 40979 43972
rect 41043 43908 41063 43972
rect 34764 43892 41063 43908
rect 34764 43828 40979 43892
rect 41043 43828 41063 43892
rect 34764 43812 41063 43828
rect 34764 43748 40979 43812
rect 41043 43748 41063 43812
rect 34764 43732 41063 43748
rect 34764 43668 40979 43732
rect 41043 43668 41063 43732
rect 34764 43652 41063 43668
rect 34764 43588 40979 43652
rect 41043 43588 41063 43652
rect 34764 43572 41063 43588
rect 34764 43508 40979 43572
rect 41043 43508 41063 43572
rect 34764 43492 41063 43508
rect 34764 43428 40979 43492
rect 41043 43428 41063 43492
rect 34764 43412 41063 43428
rect 34764 43348 40979 43412
rect 41043 43348 41063 43412
rect 34764 43332 41063 43348
rect 34764 43268 40979 43332
rect 41043 43268 41063 43332
rect 34764 43252 41063 43268
rect 34764 43188 40979 43252
rect 41043 43188 41063 43252
rect 34764 43172 41063 43188
rect 34764 43108 40979 43172
rect 41043 43108 41063 43172
rect 34764 43092 41063 43108
rect 34764 43028 40979 43092
rect 41043 43028 41063 43092
rect 34764 43012 41063 43028
rect 34764 42948 40979 43012
rect 41043 42948 41063 43012
rect 34764 42932 41063 42948
rect 34764 42868 40979 42932
rect 41043 42868 41063 42932
rect 34764 42852 41063 42868
rect 34764 42788 40979 42852
rect 41043 42788 41063 42852
rect 34764 42772 41063 42788
rect 34764 42708 40979 42772
rect 41043 42708 41063 42772
rect 34764 42692 41063 42708
rect 34764 42628 40979 42692
rect 41043 42628 41063 42692
rect 34764 42612 41063 42628
rect 34764 42548 40979 42612
rect 41043 42548 41063 42612
rect 34764 42532 41063 42548
rect 34764 42468 40979 42532
rect 41043 42468 41063 42532
rect 34764 42452 41063 42468
rect 34764 42388 40979 42452
rect 41043 42388 41063 42452
rect 34764 42372 41063 42388
rect 34764 42308 40979 42372
rect 41043 42308 41063 42372
rect 34764 42292 41063 42308
rect 34764 42228 40979 42292
rect 41043 42228 41063 42292
rect 34764 42212 41063 42228
rect 34764 42148 40979 42212
rect 41043 42148 41063 42212
rect 34764 42132 41063 42148
rect 34764 42068 40979 42132
rect 41043 42068 41063 42132
rect 34764 42052 41063 42068
rect 34764 41988 40979 42052
rect 41043 41988 41063 42052
rect 34764 41972 41063 41988
rect 34764 41908 40979 41972
rect 41043 41908 41063 41972
rect 34764 41892 41063 41908
rect 34764 41828 40979 41892
rect 41043 41828 41063 41892
rect 34764 41812 41063 41828
rect 34764 41748 40979 41812
rect 41043 41748 41063 41812
rect 34764 41732 41063 41748
rect 34764 41668 40979 41732
rect 41043 41668 41063 41732
rect 34764 41652 41063 41668
rect 34764 41588 40979 41652
rect 41043 41588 41063 41652
rect 34764 41572 41063 41588
rect 34764 41508 40979 41572
rect 41043 41508 41063 41572
rect 34764 41492 41063 41508
rect 34764 41428 40979 41492
rect 41043 41428 41063 41492
rect 34764 41412 41063 41428
rect 34764 41348 40979 41412
rect 41043 41348 41063 41412
rect 34764 41332 41063 41348
rect 34764 41268 40979 41332
rect 41043 41268 41063 41332
rect 34764 41252 41063 41268
rect 34764 41188 40979 41252
rect 41043 41188 41063 41252
rect 34764 41172 41063 41188
rect 34764 41108 40979 41172
rect 41043 41108 41063 41172
rect 34764 41092 41063 41108
rect 34764 41028 40979 41092
rect 41043 41028 41063 41092
rect 34764 41000 41063 41028
rect 41083 47172 47382 47200
rect 41083 47108 47298 47172
rect 47362 47108 47382 47172
rect 41083 47092 47382 47108
rect 41083 47028 47298 47092
rect 47362 47028 47382 47092
rect 41083 47012 47382 47028
rect 41083 46948 47298 47012
rect 47362 46948 47382 47012
rect 41083 46932 47382 46948
rect 41083 46868 47298 46932
rect 47362 46868 47382 46932
rect 41083 46852 47382 46868
rect 41083 46788 47298 46852
rect 47362 46788 47382 46852
rect 41083 46772 47382 46788
rect 41083 46708 47298 46772
rect 47362 46708 47382 46772
rect 41083 46692 47382 46708
rect 41083 46628 47298 46692
rect 47362 46628 47382 46692
rect 41083 46612 47382 46628
rect 41083 46548 47298 46612
rect 47362 46548 47382 46612
rect 41083 46532 47382 46548
rect 41083 46468 47298 46532
rect 47362 46468 47382 46532
rect 41083 46452 47382 46468
rect 41083 46388 47298 46452
rect 47362 46388 47382 46452
rect 41083 46372 47382 46388
rect 41083 46308 47298 46372
rect 47362 46308 47382 46372
rect 41083 46292 47382 46308
rect 41083 46228 47298 46292
rect 47362 46228 47382 46292
rect 41083 46212 47382 46228
rect 41083 46148 47298 46212
rect 47362 46148 47382 46212
rect 41083 46132 47382 46148
rect 41083 46068 47298 46132
rect 47362 46068 47382 46132
rect 41083 46052 47382 46068
rect 41083 45988 47298 46052
rect 47362 45988 47382 46052
rect 41083 45972 47382 45988
rect 41083 45908 47298 45972
rect 47362 45908 47382 45972
rect 41083 45892 47382 45908
rect 41083 45828 47298 45892
rect 47362 45828 47382 45892
rect 41083 45812 47382 45828
rect 41083 45748 47298 45812
rect 47362 45748 47382 45812
rect 41083 45732 47382 45748
rect 41083 45668 47298 45732
rect 47362 45668 47382 45732
rect 41083 45652 47382 45668
rect 41083 45588 47298 45652
rect 47362 45588 47382 45652
rect 41083 45572 47382 45588
rect 41083 45508 47298 45572
rect 47362 45508 47382 45572
rect 41083 45492 47382 45508
rect 41083 45428 47298 45492
rect 47362 45428 47382 45492
rect 41083 45412 47382 45428
rect 41083 45348 47298 45412
rect 47362 45348 47382 45412
rect 41083 45332 47382 45348
rect 41083 45268 47298 45332
rect 47362 45268 47382 45332
rect 41083 45252 47382 45268
rect 41083 45188 47298 45252
rect 47362 45188 47382 45252
rect 41083 45172 47382 45188
rect 41083 45108 47298 45172
rect 47362 45108 47382 45172
rect 41083 45092 47382 45108
rect 41083 45028 47298 45092
rect 47362 45028 47382 45092
rect 41083 45012 47382 45028
rect 41083 44948 47298 45012
rect 47362 44948 47382 45012
rect 41083 44932 47382 44948
rect 41083 44868 47298 44932
rect 47362 44868 47382 44932
rect 41083 44852 47382 44868
rect 41083 44788 47298 44852
rect 47362 44788 47382 44852
rect 41083 44772 47382 44788
rect 41083 44708 47298 44772
rect 47362 44708 47382 44772
rect 41083 44692 47382 44708
rect 41083 44628 47298 44692
rect 47362 44628 47382 44692
rect 41083 44612 47382 44628
rect 41083 44548 47298 44612
rect 47362 44548 47382 44612
rect 41083 44532 47382 44548
rect 41083 44468 47298 44532
rect 47362 44468 47382 44532
rect 41083 44452 47382 44468
rect 41083 44388 47298 44452
rect 47362 44388 47382 44452
rect 41083 44372 47382 44388
rect 41083 44308 47298 44372
rect 47362 44308 47382 44372
rect 41083 44292 47382 44308
rect 41083 44228 47298 44292
rect 47362 44228 47382 44292
rect 41083 44212 47382 44228
rect 41083 44148 47298 44212
rect 47362 44148 47382 44212
rect 41083 44132 47382 44148
rect 41083 44068 47298 44132
rect 47362 44068 47382 44132
rect 41083 44052 47382 44068
rect 41083 43988 47298 44052
rect 47362 43988 47382 44052
rect 41083 43972 47382 43988
rect 41083 43908 47298 43972
rect 47362 43908 47382 43972
rect 41083 43892 47382 43908
rect 41083 43828 47298 43892
rect 47362 43828 47382 43892
rect 41083 43812 47382 43828
rect 41083 43748 47298 43812
rect 47362 43748 47382 43812
rect 41083 43732 47382 43748
rect 41083 43668 47298 43732
rect 47362 43668 47382 43732
rect 41083 43652 47382 43668
rect 41083 43588 47298 43652
rect 47362 43588 47382 43652
rect 41083 43572 47382 43588
rect 41083 43508 47298 43572
rect 47362 43508 47382 43572
rect 41083 43492 47382 43508
rect 41083 43428 47298 43492
rect 47362 43428 47382 43492
rect 41083 43412 47382 43428
rect 41083 43348 47298 43412
rect 47362 43348 47382 43412
rect 41083 43332 47382 43348
rect 41083 43268 47298 43332
rect 47362 43268 47382 43332
rect 41083 43252 47382 43268
rect 41083 43188 47298 43252
rect 47362 43188 47382 43252
rect 41083 43172 47382 43188
rect 41083 43108 47298 43172
rect 47362 43108 47382 43172
rect 41083 43092 47382 43108
rect 41083 43028 47298 43092
rect 47362 43028 47382 43092
rect 41083 43012 47382 43028
rect 41083 42948 47298 43012
rect 47362 42948 47382 43012
rect 41083 42932 47382 42948
rect 41083 42868 47298 42932
rect 47362 42868 47382 42932
rect 41083 42852 47382 42868
rect 41083 42788 47298 42852
rect 47362 42788 47382 42852
rect 41083 42772 47382 42788
rect 41083 42708 47298 42772
rect 47362 42708 47382 42772
rect 41083 42692 47382 42708
rect 41083 42628 47298 42692
rect 47362 42628 47382 42692
rect 41083 42612 47382 42628
rect 41083 42548 47298 42612
rect 47362 42548 47382 42612
rect 41083 42532 47382 42548
rect 41083 42468 47298 42532
rect 47362 42468 47382 42532
rect 41083 42452 47382 42468
rect 41083 42388 47298 42452
rect 47362 42388 47382 42452
rect 41083 42372 47382 42388
rect 41083 42308 47298 42372
rect 47362 42308 47382 42372
rect 41083 42292 47382 42308
rect 41083 42228 47298 42292
rect 47362 42228 47382 42292
rect 41083 42212 47382 42228
rect 41083 42148 47298 42212
rect 47362 42148 47382 42212
rect 41083 42132 47382 42148
rect 41083 42068 47298 42132
rect 47362 42068 47382 42132
rect 41083 42052 47382 42068
rect 41083 41988 47298 42052
rect 47362 41988 47382 42052
rect 41083 41972 47382 41988
rect 41083 41908 47298 41972
rect 47362 41908 47382 41972
rect 41083 41892 47382 41908
rect 41083 41828 47298 41892
rect 47362 41828 47382 41892
rect 41083 41812 47382 41828
rect 41083 41748 47298 41812
rect 47362 41748 47382 41812
rect 41083 41732 47382 41748
rect 41083 41668 47298 41732
rect 47362 41668 47382 41732
rect 41083 41652 47382 41668
rect 41083 41588 47298 41652
rect 47362 41588 47382 41652
rect 41083 41572 47382 41588
rect 41083 41508 47298 41572
rect 47362 41508 47382 41572
rect 41083 41492 47382 41508
rect 41083 41428 47298 41492
rect 47362 41428 47382 41492
rect 41083 41412 47382 41428
rect 41083 41348 47298 41412
rect 47362 41348 47382 41412
rect 41083 41332 47382 41348
rect 41083 41268 47298 41332
rect 47362 41268 47382 41332
rect 41083 41252 47382 41268
rect 41083 41188 47298 41252
rect 47362 41188 47382 41252
rect 41083 41172 47382 41188
rect 41083 41108 47298 41172
rect 47362 41108 47382 41172
rect 41083 41092 47382 41108
rect 41083 41028 47298 41092
rect 47362 41028 47382 41092
rect 41083 41000 47382 41028
rect -47383 40872 -41084 40900
rect -47383 40808 -41168 40872
rect -41104 40808 -41084 40872
rect -47383 40792 -41084 40808
rect -47383 40728 -41168 40792
rect -41104 40728 -41084 40792
rect -47383 40712 -41084 40728
rect -47383 40648 -41168 40712
rect -41104 40648 -41084 40712
rect -47383 40632 -41084 40648
rect -47383 40568 -41168 40632
rect -41104 40568 -41084 40632
rect -47383 40552 -41084 40568
rect -47383 40488 -41168 40552
rect -41104 40488 -41084 40552
rect -47383 40472 -41084 40488
rect -47383 40408 -41168 40472
rect -41104 40408 -41084 40472
rect -47383 40392 -41084 40408
rect -47383 40328 -41168 40392
rect -41104 40328 -41084 40392
rect -47383 40312 -41084 40328
rect -47383 40248 -41168 40312
rect -41104 40248 -41084 40312
rect -47383 40232 -41084 40248
rect -47383 40168 -41168 40232
rect -41104 40168 -41084 40232
rect -47383 40152 -41084 40168
rect -47383 40088 -41168 40152
rect -41104 40088 -41084 40152
rect -47383 40072 -41084 40088
rect -47383 40008 -41168 40072
rect -41104 40008 -41084 40072
rect -47383 39992 -41084 40008
rect -47383 39928 -41168 39992
rect -41104 39928 -41084 39992
rect -47383 39912 -41084 39928
rect -47383 39848 -41168 39912
rect -41104 39848 -41084 39912
rect -47383 39832 -41084 39848
rect -47383 39768 -41168 39832
rect -41104 39768 -41084 39832
rect -47383 39752 -41084 39768
rect -47383 39688 -41168 39752
rect -41104 39688 -41084 39752
rect -47383 39672 -41084 39688
rect -47383 39608 -41168 39672
rect -41104 39608 -41084 39672
rect -47383 39592 -41084 39608
rect -47383 39528 -41168 39592
rect -41104 39528 -41084 39592
rect -47383 39512 -41084 39528
rect -47383 39448 -41168 39512
rect -41104 39448 -41084 39512
rect -47383 39432 -41084 39448
rect -47383 39368 -41168 39432
rect -41104 39368 -41084 39432
rect -47383 39352 -41084 39368
rect -47383 39288 -41168 39352
rect -41104 39288 -41084 39352
rect -47383 39272 -41084 39288
rect -47383 39208 -41168 39272
rect -41104 39208 -41084 39272
rect -47383 39192 -41084 39208
rect -47383 39128 -41168 39192
rect -41104 39128 -41084 39192
rect -47383 39112 -41084 39128
rect -47383 39048 -41168 39112
rect -41104 39048 -41084 39112
rect -47383 39032 -41084 39048
rect -47383 38968 -41168 39032
rect -41104 38968 -41084 39032
rect -47383 38952 -41084 38968
rect -47383 38888 -41168 38952
rect -41104 38888 -41084 38952
rect -47383 38872 -41084 38888
rect -47383 38808 -41168 38872
rect -41104 38808 -41084 38872
rect -47383 38792 -41084 38808
rect -47383 38728 -41168 38792
rect -41104 38728 -41084 38792
rect -47383 38712 -41084 38728
rect -47383 38648 -41168 38712
rect -41104 38648 -41084 38712
rect -47383 38632 -41084 38648
rect -47383 38568 -41168 38632
rect -41104 38568 -41084 38632
rect -47383 38552 -41084 38568
rect -47383 38488 -41168 38552
rect -41104 38488 -41084 38552
rect -47383 38472 -41084 38488
rect -47383 38408 -41168 38472
rect -41104 38408 -41084 38472
rect -47383 38392 -41084 38408
rect -47383 38328 -41168 38392
rect -41104 38328 -41084 38392
rect -47383 38312 -41084 38328
rect -47383 38248 -41168 38312
rect -41104 38248 -41084 38312
rect -47383 38232 -41084 38248
rect -47383 38168 -41168 38232
rect -41104 38168 -41084 38232
rect -47383 38152 -41084 38168
rect -47383 38088 -41168 38152
rect -41104 38088 -41084 38152
rect -47383 38072 -41084 38088
rect -47383 38008 -41168 38072
rect -41104 38008 -41084 38072
rect -47383 37992 -41084 38008
rect -47383 37928 -41168 37992
rect -41104 37928 -41084 37992
rect -47383 37912 -41084 37928
rect -47383 37848 -41168 37912
rect -41104 37848 -41084 37912
rect -47383 37832 -41084 37848
rect -47383 37768 -41168 37832
rect -41104 37768 -41084 37832
rect -47383 37752 -41084 37768
rect -47383 37688 -41168 37752
rect -41104 37688 -41084 37752
rect -47383 37672 -41084 37688
rect -47383 37608 -41168 37672
rect -41104 37608 -41084 37672
rect -47383 37592 -41084 37608
rect -47383 37528 -41168 37592
rect -41104 37528 -41084 37592
rect -47383 37512 -41084 37528
rect -47383 37448 -41168 37512
rect -41104 37448 -41084 37512
rect -47383 37432 -41084 37448
rect -47383 37368 -41168 37432
rect -41104 37368 -41084 37432
rect -47383 37352 -41084 37368
rect -47383 37288 -41168 37352
rect -41104 37288 -41084 37352
rect -47383 37272 -41084 37288
rect -47383 37208 -41168 37272
rect -41104 37208 -41084 37272
rect -47383 37192 -41084 37208
rect -47383 37128 -41168 37192
rect -41104 37128 -41084 37192
rect -47383 37112 -41084 37128
rect -47383 37048 -41168 37112
rect -41104 37048 -41084 37112
rect -47383 37032 -41084 37048
rect -47383 36968 -41168 37032
rect -41104 36968 -41084 37032
rect -47383 36952 -41084 36968
rect -47383 36888 -41168 36952
rect -41104 36888 -41084 36952
rect -47383 36872 -41084 36888
rect -47383 36808 -41168 36872
rect -41104 36808 -41084 36872
rect -47383 36792 -41084 36808
rect -47383 36728 -41168 36792
rect -41104 36728 -41084 36792
rect -47383 36712 -41084 36728
rect -47383 36648 -41168 36712
rect -41104 36648 -41084 36712
rect -47383 36632 -41084 36648
rect -47383 36568 -41168 36632
rect -41104 36568 -41084 36632
rect -47383 36552 -41084 36568
rect -47383 36488 -41168 36552
rect -41104 36488 -41084 36552
rect -47383 36472 -41084 36488
rect -47383 36408 -41168 36472
rect -41104 36408 -41084 36472
rect -47383 36392 -41084 36408
rect -47383 36328 -41168 36392
rect -41104 36328 -41084 36392
rect -47383 36312 -41084 36328
rect -47383 36248 -41168 36312
rect -41104 36248 -41084 36312
rect -47383 36232 -41084 36248
rect -47383 36168 -41168 36232
rect -41104 36168 -41084 36232
rect -47383 36152 -41084 36168
rect -47383 36088 -41168 36152
rect -41104 36088 -41084 36152
rect -47383 36072 -41084 36088
rect -47383 36008 -41168 36072
rect -41104 36008 -41084 36072
rect -47383 35992 -41084 36008
rect -47383 35928 -41168 35992
rect -41104 35928 -41084 35992
rect -47383 35912 -41084 35928
rect -47383 35848 -41168 35912
rect -41104 35848 -41084 35912
rect -47383 35832 -41084 35848
rect -47383 35768 -41168 35832
rect -41104 35768 -41084 35832
rect -47383 35752 -41084 35768
rect -47383 35688 -41168 35752
rect -41104 35688 -41084 35752
rect -47383 35672 -41084 35688
rect -47383 35608 -41168 35672
rect -41104 35608 -41084 35672
rect -47383 35592 -41084 35608
rect -47383 35528 -41168 35592
rect -41104 35528 -41084 35592
rect -47383 35512 -41084 35528
rect -47383 35448 -41168 35512
rect -41104 35448 -41084 35512
rect -47383 35432 -41084 35448
rect -47383 35368 -41168 35432
rect -41104 35368 -41084 35432
rect -47383 35352 -41084 35368
rect -47383 35288 -41168 35352
rect -41104 35288 -41084 35352
rect -47383 35272 -41084 35288
rect -47383 35208 -41168 35272
rect -41104 35208 -41084 35272
rect -47383 35192 -41084 35208
rect -47383 35128 -41168 35192
rect -41104 35128 -41084 35192
rect -47383 35112 -41084 35128
rect -47383 35048 -41168 35112
rect -41104 35048 -41084 35112
rect -47383 35032 -41084 35048
rect -47383 34968 -41168 35032
rect -41104 34968 -41084 35032
rect -47383 34952 -41084 34968
rect -47383 34888 -41168 34952
rect -41104 34888 -41084 34952
rect -47383 34872 -41084 34888
rect -47383 34808 -41168 34872
rect -41104 34808 -41084 34872
rect -47383 34792 -41084 34808
rect -47383 34728 -41168 34792
rect -41104 34728 -41084 34792
rect -47383 34700 -41084 34728
rect -41064 40872 -34765 40900
rect -41064 40808 -34849 40872
rect -34785 40808 -34765 40872
rect -41064 40792 -34765 40808
rect -41064 40728 -34849 40792
rect -34785 40728 -34765 40792
rect -41064 40712 -34765 40728
rect -41064 40648 -34849 40712
rect -34785 40648 -34765 40712
rect -41064 40632 -34765 40648
rect -41064 40568 -34849 40632
rect -34785 40568 -34765 40632
rect -41064 40552 -34765 40568
rect -41064 40488 -34849 40552
rect -34785 40488 -34765 40552
rect -41064 40472 -34765 40488
rect -41064 40408 -34849 40472
rect -34785 40408 -34765 40472
rect -41064 40392 -34765 40408
rect -41064 40328 -34849 40392
rect -34785 40328 -34765 40392
rect -41064 40312 -34765 40328
rect -41064 40248 -34849 40312
rect -34785 40248 -34765 40312
rect -41064 40232 -34765 40248
rect -41064 40168 -34849 40232
rect -34785 40168 -34765 40232
rect -41064 40152 -34765 40168
rect -41064 40088 -34849 40152
rect -34785 40088 -34765 40152
rect -41064 40072 -34765 40088
rect -41064 40008 -34849 40072
rect -34785 40008 -34765 40072
rect -41064 39992 -34765 40008
rect -41064 39928 -34849 39992
rect -34785 39928 -34765 39992
rect -41064 39912 -34765 39928
rect -41064 39848 -34849 39912
rect -34785 39848 -34765 39912
rect -41064 39832 -34765 39848
rect -41064 39768 -34849 39832
rect -34785 39768 -34765 39832
rect -41064 39752 -34765 39768
rect -41064 39688 -34849 39752
rect -34785 39688 -34765 39752
rect -41064 39672 -34765 39688
rect -41064 39608 -34849 39672
rect -34785 39608 -34765 39672
rect -41064 39592 -34765 39608
rect -41064 39528 -34849 39592
rect -34785 39528 -34765 39592
rect -41064 39512 -34765 39528
rect -41064 39448 -34849 39512
rect -34785 39448 -34765 39512
rect -41064 39432 -34765 39448
rect -41064 39368 -34849 39432
rect -34785 39368 -34765 39432
rect -41064 39352 -34765 39368
rect -41064 39288 -34849 39352
rect -34785 39288 -34765 39352
rect -41064 39272 -34765 39288
rect -41064 39208 -34849 39272
rect -34785 39208 -34765 39272
rect -41064 39192 -34765 39208
rect -41064 39128 -34849 39192
rect -34785 39128 -34765 39192
rect -41064 39112 -34765 39128
rect -41064 39048 -34849 39112
rect -34785 39048 -34765 39112
rect -41064 39032 -34765 39048
rect -41064 38968 -34849 39032
rect -34785 38968 -34765 39032
rect -41064 38952 -34765 38968
rect -41064 38888 -34849 38952
rect -34785 38888 -34765 38952
rect -41064 38872 -34765 38888
rect -41064 38808 -34849 38872
rect -34785 38808 -34765 38872
rect -41064 38792 -34765 38808
rect -41064 38728 -34849 38792
rect -34785 38728 -34765 38792
rect -41064 38712 -34765 38728
rect -41064 38648 -34849 38712
rect -34785 38648 -34765 38712
rect -41064 38632 -34765 38648
rect -41064 38568 -34849 38632
rect -34785 38568 -34765 38632
rect -41064 38552 -34765 38568
rect -41064 38488 -34849 38552
rect -34785 38488 -34765 38552
rect -41064 38472 -34765 38488
rect -41064 38408 -34849 38472
rect -34785 38408 -34765 38472
rect -41064 38392 -34765 38408
rect -41064 38328 -34849 38392
rect -34785 38328 -34765 38392
rect -41064 38312 -34765 38328
rect -41064 38248 -34849 38312
rect -34785 38248 -34765 38312
rect -41064 38232 -34765 38248
rect -41064 38168 -34849 38232
rect -34785 38168 -34765 38232
rect -41064 38152 -34765 38168
rect -41064 38088 -34849 38152
rect -34785 38088 -34765 38152
rect -41064 38072 -34765 38088
rect -41064 38008 -34849 38072
rect -34785 38008 -34765 38072
rect -41064 37992 -34765 38008
rect -41064 37928 -34849 37992
rect -34785 37928 -34765 37992
rect -41064 37912 -34765 37928
rect -41064 37848 -34849 37912
rect -34785 37848 -34765 37912
rect -41064 37832 -34765 37848
rect -41064 37768 -34849 37832
rect -34785 37768 -34765 37832
rect -41064 37752 -34765 37768
rect -41064 37688 -34849 37752
rect -34785 37688 -34765 37752
rect -41064 37672 -34765 37688
rect -41064 37608 -34849 37672
rect -34785 37608 -34765 37672
rect -41064 37592 -34765 37608
rect -41064 37528 -34849 37592
rect -34785 37528 -34765 37592
rect -41064 37512 -34765 37528
rect -41064 37448 -34849 37512
rect -34785 37448 -34765 37512
rect -41064 37432 -34765 37448
rect -41064 37368 -34849 37432
rect -34785 37368 -34765 37432
rect -41064 37352 -34765 37368
rect -41064 37288 -34849 37352
rect -34785 37288 -34765 37352
rect -41064 37272 -34765 37288
rect -41064 37208 -34849 37272
rect -34785 37208 -34765 37272
rect -41064 37192 -34765 37208
rect -41064 37128 -34849 37192
rect -34785 37128 -34765 37192
rect -41064 37112 -34765 37128
rect -41064 37048 -34849 37112
rect -34785 37048 -34765 37112
rect -41064 37032 -34765 37048
rect -41064 36968 -34849 37032
rect -34785 36968 -34765 37032
rect -41064 36952 -34765 36968
rect -41064 36888 -34849 36952
rect -34785 36888 -34765 36952
rect -41064 36872 -34765 36888
rect -41064 36808 -34849 36872
rect -34785 36808 -34765 36872
rect -41064 36792 -34765 36808
rect -41064 36728 -34849 36792
rect -34785 36728 -34765 36792
rect -41064 36712 -34765 36728
rect -41064 36648 -34849 36712
rect -34785 36648 -34765 36712
rect -41064 36632 -34765 36648
rect -41064 36568 -34849 36632
rect -34785 36568 -34765 36632
rect -41064 36552 -34765 36568
rect -41064 36488 -34849 36552
rect -34785 36488 -34765 36552
rect -41064 36472 -34765 36488
rect -41064 36408 -34849 36472
rect -34785 36408 -34765 36472
rect -41064 36392 -34765 36408
rect -41064 36328 -34849 36392
rect -34785 36328 -34765 36392
rect -41064 36312 -34765 36328
rect -41064 36248 -34849 36312
rect -34785 36248 -34765 36312
rect -41064 36232 -34765 36248
rect -41064 36168 -34849 36232
rect -34785 36168 -34765 36232
rect -41064 36152 -34765 36168
rect -41064 36088 -34849 36152
rect -34785 36088 -34765 36152
rect -41064 36072 -34765 36088
rect -41064 36008 -34849 36072
rect -34785 36008 -34765 36072
rect -41064 35992 -34765 36008
rect -41064 35928 -34849 35992
rect -34785 35928 -34765 35992
rect -41064 35912 -34765 35928
rect -41064 35848 -34849 35912
rect -34785 35848 -34765 35912
rect -41064 35832 -34765 35848
rect -41064 35768 -34849 35832
rect -34785 35768 -34765 35832
rect -41064 35752 -34765 35768
rect -41064 35688 -34849 35752
rect -34785 35688 -34765 35752
rect -41064 35672 -34765 35688
rect -41064 35608 -34849 35672
rect -34785 35608 -34765 35672
rect -41064 35592 -34765 35608
rect -41064 35528 -34849 35592
rect -34785 35528 -34765 35592
rect -41064 35512 -34765 35528
rect -41064 35448 -34849 35512
rect -34785 35448 -34765 35512
rect -41064 35432 -34765 35448
rect -41064 35368 -34849 35432
rect -34785 35368 -34765 35432
rect -41064 35352 -34765 35368
rect -41064 35288 -34849 35352
rect -34785 35288 -34765 35352
rect -41064 35272 -34765 35288
rect -41064 35208 -34849 35272
rect -34785 35208 -34765 35272
rect -41064 35192 -34765 35208
rect -41064 35128 -34849 35192
rect -34785 35128 -34765 35192
rect -41064 35112 -34765 35128
rect -41064 35048 -34849 35112
rect -34785 35048 -34765 35112
rect -41064 35032 -34765 35048
rect -41064 34968 -34849 35032
rect -34785 34968 -34765 35032
rect -41064 34952 -34765 34968
rect -41064 34888 -34849 34952
rect -34785 34888 -34765 34952
rect -41064 34872 -34765 34888
rect -41064 34808 -34849 34872
rect -34785 34808 -34765 34872
rect -41064 34792 -34765 34808
rect -41064 34728 -34849 34792
rect -34785 34728 -34765 34792
rect -41064 34700 -34765 34728
rect -34745 40872 -28446 40900
rect -34745 40808 -28530 40872
rect -28466 40808 -28446 40872
rect -34745 40792 -28446 40808
rect -34745 40728 -28530 40792
rect -28466 40728 -28446 40792
rect -34745 40712 -28446 40728
rect -34745 40648 -28530 40712
rect -28466 40648 -28446 40712
rect -34745 40632 -28446 40648
rect -34745 40568 -28530 40632
rect -28466 40568 -28446 40632
rect -34745 40552 -28446 40568
rect -34745 40488 -28530 40552
rect -28466 40488 -28446 40552
rect -34745 40472 -28446 40488
rect -34745 40408 -28530 40472
rect -28466 40408 -28446 40472
rect -34745 40392 -28446 40408
rect -34745 40328 -28530 40392
rect -28466 40328 -28446 40392
rect -34745 40312 -28446 40328
rect -34745 40248 -28530 40312
rect -28466 40248 -28446 40312
rect -34745 40232 -28446 40248
rect -34745 40168 -28530 40232
rect -28466 40168 -28446 40232
rect -34745 40152 -28446 40168
rect -34745 40088 -28530 40152
rect -28466 40088 -28446 40152
rect -34745 40072 -28446 40088
rect -34745 40008 -28530 40072
rect -28466 40008 -28446 40072
rect -34745 39992 -28446 40008
rect -34745 39928 -28530 39992
rect -28466 39928 -28446 39992
rect -34745 39912 -28446 39928
rect -34745 39848 -28530 39912
rect -28466 39848 -28446 39912
rect -34745 39832 -28446 39848
rect -34745 39768 -28530 39832
rect -28466 39768 -28446 39832
rect -34745 39752 -28446 39768
rect -34745 39688 -28530 39752
rect -28466 39688 -28446 39752
rect -34745 39672 -28446 39688
rect -34745 39608 -28530 39672
rect -28466 39608 -28446 39672
rect -34745 39592 -28446 39608
rect -34745 39528 -28530 39592
rect -28466 39528 -28446 39592
rect -34745 39512 -28446 39528
rect -34745 39448 -28530 39512
rect -28466 39448 -28446 39512
rect -34745 39432 -28446 39448
rect -34745 39368 -28530 39432
rect -28466 39368 -28446 39432
rect -34745 39352 -28446 39368
rect -34745 39288 -28530 39352
rect -28466 39288 -28446 39352
rect -34745 39272 -28446 39288
rect -34745 39208 -28530 39272
rect -28466 39208 -28446 39272
rect -34745 39192 -28446 39208
rect -34745 39128 -28530 39192
rect -28466 39128 -28446 39192
rect -34745 39112 -28446 39128
rect -34745 39048 -28530 39112
rect -28466 39048 -28446 39112
rect -34745 39032 -28446 39048
rect -34745 38968 -28530 39032
rect -28466 38968 -28446 39032
rect -34745 38952 -28446 38968
rect -34745 38888 -28530 38952
rect -28466 38888 -28446 38952
rect -34745 38872 -28446 38888
rect -34745 38808 -28530 38872
rect -28466 38808 -28446 38872
rect -34745 38792 -28446 38808
rect -34745 38728 -28530 38792
rect -28466 38728 -28446 38792
rect -34745 38712 -28446 38728
rect -34745 38648 -28530 38712
rect -28466 38648 -28446 38712
rect -34745 38632 -28446 38648
rect -34745 38568 -28530 38632
rect -28466 38568 -28446 38632
rect -34745 38552 -28446 38568
rect -34745 38488 -28530 38552
rect -28466 38488 -28446 38552
rect -34745 38472 -28446 38488
rect -34745 38408 -28530 38472
rect -28466 38408 -28446 38472
rect -34745 38392 -28446 38408
rect -34745 38328 -28530 38392
rect -28466 38328 -28446 38392
rect -34745 38312 -28446 38328
rect -34745 38248 -28530 38312
rect -28466 38248 -28446 38312
rect -34745 38232 -28446 38248
rect -34745 38168 -28530 38232
rect -28466 38168 -28446 38232
rect -34745 38152 -28446 38168
rect -34745 38088 -28530 38152
rect -28466 38088 -28446 38152
rect -34745 38072 -28446 38088
rect -34745 38008 -28530 38072
rect -28466 38008 -28446 38072
rect -34745 37992 -28446 38008
rect -34745 37928 -28530 37992
rect -28466 37928 -28446 37992
rect -34745 37912 -28446 37928
rect -34745 37848 -28530 37912
rect -28466 37848 -28446 37912
rect -34745 37832 -28446 37848
rect -34745 37768 -28530 37832
rect -28466 37768 -28446 37832
rect -34745 37752 -28446 37768
rect -34745 37688 -28530 37752
rect -28466 37688 -28446 37752
rect -34745 37672 -28446 37688
rect -34745 37608 -28530 37672
rect -28466 37608 -28446 37672
rect -34745 37592 -28446 37608
rect -34745 37528 -28530 37592
rect -28466 37528 -28446 37592
rect -34745 37512 -28446 37528
rect -34745 37448 -28530 37512
rect -28466 37448 -28446 37512
rect -34745 37432 -28446 37448
rect -34745 37368 -28530 37432
rect -28466 37368 -28446 37432
rect -34745 37352 -28446 37368
rect -34745 37288 -28530 37352
rect -28466 37288 -28446 37352
rect -34745 37272 -28446 37288
rect -34745 37208 -28530 37272
rect -28466 37208 -28446 37272
rect -34745 37192 -28446 37208
rect -34745 37128 -28530 37192
rect -28466 37128 -28446 37192
rect -34745 37112 -28446 37128
rect -34745 37048 -28530 37112
rect -28466 37048 -28446 37112
rect -34745 37032 -28446 37048
rect -34745 36968 -28530 37032
rect -28466 36968 -28446 37032
rect -34745 36952 -28446 36968
rect -34745 36888 -28530 36952
rect -28466 36888 -28446 36952
rect -34745 36872 -28446 36888
rect -34745 36808 -28530 36872
rect -28466 36808 -28446 36872
rect -34745 36792 -28446 36808
rect -34745 36728 -28530 36792
rect -28466 36728 -28446 36792
rect -34745 36712 -28446 36728
rect -34745 36648 -28530 36712
rect -28466 36648 -28446 36712
rect -34745 36632 -28446 36648
rect -34745 36568 -28530 36632
rect -28466 36568 -28446 36632
rect -34745 36552 -28446 36568
rect -34745 36488 -28530 36552
rect -28466 36488 -28446 36552
rect -34745 36472 -28446 36488
rect -34745 36408 -28530 36472
rect -28466 36408 -28446 36472
rect -34745 36392 -28446 36408
rect -34745 36328 -28530 36392
rect -28466 36328 -28446 36392
rect -34745 36312 -28446 36328
rect -34745 36248 -28530 36312
rect -28466 36248 -28446 36312
rect -34745 36232 -28446 36248
rect -34745 36168 -28530 36232
rect -28466 36168 -28446 36232
rect -34745 36152 -28446 36168
rect -34745 36088 -28530 36152
rect -28466 36088 -28446 36152
rect -34745 36072 -28446 36088
rect -34745 36008 -28530 36072
rect -28466 36008 -28446 36072
rect -34745 35992 -28446 36008
rect -34745 35928 -28530 35992
rect -28466 35928 -28446 35992
rect -34745 35912 -28446 35928
rect -34745 35848 -28530 35912
rect -28466 35848 -28446 35912
rect -34745 35832 -28446 35848
rect -34745 35768 -28530 35832
rect -28466 35768 -28446 35832
rect -34745 35752 -28446 35768
rect -34745 35688 -28530 35752
rect -28466 35688 -28446 35752
rect -34745 35672 -28446 35688
rect -34745 35608 -28530 35672
rect -28466 35608 -28446 35672
rect -34745 35592 -28446 35608
rect -34745 35528 -28530 35592
rect -28466 35528 -28446 35592
rect -34745 35512 -28446 35528
rect -34745 35448 -28530 35512
rect -28466 35448 -28446 35512
rect -34745 35432 -28446 35448
rect -34745 35368 -28530 35432
rect -28466 35368 -28446 35432
rect -34745 35352 -28446 35368
rect -34745 35288 -28530 35352
rect -28466 35288 -28446 35352
rect -34745 35272 -28446 35288
rect -34745 35208 -28530 35272
rect -28466 35208 -28446 35272
rect -34745 35192 -28446 35208
rect -34745 35128 -28530 35192
rect -28466 35128 -28446 35192
rect -34745 35112 -28446 35128
rect -34745 35048 -28530 35112
rect -28466 35048 -28446 35112
rect -34745 35032 -28446 35048
rect -34745 34968 -28530 35032
rect -28466 34968 -28446 35032
rect -34745 34952 -28446 34968
rect -34745 34888 -28530 34952
rect -28466 34888 -28446 34952
rect -34745 34872 -28446 34888
rect -34745 34808 -28530 34872
rect -28466 34808 -28446 34872
rect -34745 34792 -28446 34808
rect -34745 34728 -28530 34792
rect -28466 34728 -28446 34792
rect -34745 34700 -28446 34728
rect -28426 40872 -22127 40900
rect -28426 40808 -22211 40872
rect -22147 40808 -22127 40872
rect -28426 40792 -22127 40808
rect -28426 40728 -22211 40792
rect -22147 40728 -22127 40792
rect -28426 40712 -22127 40728
rect -28426 40648 -22211 40712
rect -22147 40648 -22127 40712
rect -28426 40632 -22127 40648
rect -28426 40568 -22211 40632
rect -22147 40568 -22127 40632
rect -28426 40552 -22127 40568
rect -28426 40488 -22211 40552
rect -22147 40488 -22127 40552
rect -28426 40472 -22127 40488
rect -28426 40408 -22211 40472
rect -22147 40408 -22127 40472
rect -28426 40392 -22127 40408
rect -28426 40328 -22211 40392
rect -22147 40328 -22127 40392
rect -28426 40312 -22127 40328
rect -28426 40248 -22211 40312
rect -22147 40248 -22127 40312
rect -28426 40232 -22127 40248
rect -28426 40168 -22211 40232
rect -22147 40168 -22127 40232
rect -28426 40152 -22127 40168
rect -28426 40088 -22211 40152
rect -22147 40088 -22127 40152
rect -28426 40072 -22127 40088
rect -28426 40008 -22211 40072
rect -22147 40008 -22127 40072
rect -28426 39992 -22127 40008
rect -28426 39928 -22211 39992
rect -22147 39928 -22127 39992
rect -28426 39912 -22127 39928
rect -28426 39848 -22211 39912
rect -22147 39848 -22127 39912
rect -28426 39832 -22127 39848
rect -28426 39768 -22211 39832
rect -22147 39768 -22127 39832
rect -28426 39752 -22127 39768
rect -28426 39688 -22211 39752
rect -22147 39688 -22127 39752
rect -28426 39672 -22127 39688
rect -28426 39608 -22211 39672
rect -22147 39608 -22127 39672
rect -28426 39592 -22127 39608
rect -28426 39528 -22211 39592
rect -22147 39528 -22127 39592
rect -28426 39512 -22127 39528
rect -28426 39448 -22211 39512
rect -22147 39448 -22127 39512
rect -28426 39432 -22127 39448
rect -28426 39368 -22211 39432
rect -22147 39368 -22127 39432
rect -28426 39352 -22127 39368
rect -28426 39288 -22211 39352
rect -22147 39288 -22127 39352
rect -28426 39272 -22127 39288
rect -28426 39208 -22211 39272
rect -22147 39208 -22127 39272
rect -28426 39192 -22127 39208
rect -28426 39128 -22211 39192
rect -22147 39128 -22127 39192
rect -28426 39112 -22127 39128
rect -28426 39048 -22211 39112
rect -22147 39048 -22127 39112
rect -28426 39032 -22127 39048
rect -28426 38968 -22211 39032
rect -22147 38968 -22127 39032
rect -28426 38952 -22127 38968
rect -28426 38888 -22211 38952
rect -22147 38888 -22127 38952
rect -28426 38872 -22127 38888
rect -28426 38808 -22211 38872
rect -22147 38808 -22127 38872
rect -28426 38792 -22127 38808
rect -28426 38728 -22211 38792
rect -22147 38728 -22127 38792
rect -28426 38712 -22127 38728
rect -28426 38648 -22211 38712
rect -22147 38648 -22127 38712
rect -28426 38632 -22127 38648
rect -28426 38568 -22211 38632
rect -22147 38568 -22127 38632
rect -28426 38552 -22127 38568
rect -28426 38488 -22211 38552
rect -22147 38488 -22127 38552
rect -28426 38472 -22127 38488
rect -28426 38408 -22211 38472
rect -22147 38408 -22127 38472
rect -28426 38392 -22127 38408
rect -28426 38328 -22211 38392
rect -22147 38328 -22127 38392
rect -28426 38312 -22127 38328
rect -28426 38248 -22211 38312
rect -22147 38248 -22127 38312
rect -28426 38232 -22127 38248
rect -28426 38168 -22211 38232
rect -22147 38168 -22127 38232
rect -28426 38152 -22127 38168
rect -28426 38088 -22211 38152
rect -22147 38088 -22127 38152
rect -28426 38072 -22127 38088
rect -28426 38008 -22211 38072
rect -22147 38008 -22127 38072
rect -28426 37992 -22127 38008
rect -28426 37928 -22211 37992
rect -22147 37928 -22127 37992
rect -28426 37912 -22127 37928
rect -28426 37848 -22211 37912
rect -22147 37848 -22127 37912
rect -28426 37832 -22127 37848
rect -28426 37768 -22211 37832
rect -22147 37768 -22127 37832
rect -28426 37752 -22127 37768
rect -28426 37688 -22211 37752
rect -22147 37688 -22127 37752
rect -28426 37672 -22127 37688
rect -28426 37608 -22211 37672
rect -22147 37608 -22127 37672
rect -28426 37592 -22127 37608
rect -28426 37528 -22211 37592
rect -22147 37528 -22127 37592
rect -28426 37512 -22127 37528
rect -28426 37448 -22211 37512
rect -22147 37448 -22127 37512
rect -28426 37432 -22127 37448
rect -28426 37368 -22211 37432
rect -22147 37368 -22127 37432
rect -28426 37352 -22127 37368
rect -28426 37288 -22211 37352
rect -22147 37288 -22127 37352
rect -28426 37272 -22127 37288
rect -28426 37208 -22211 37272
rect -22147 37208 -22127 37272
rect -28426 37192 -22127 37208
rect -28426 37128 -22211 37192
rect -22147 37128 -22127 37192
rect -28426 37112 -22127 37128
rect -28426 37048 -22211 37112
rect -22147 37048 -22127 37112
rect -28426 37032 -22127 37048
rect -28426 36968 -22211 37032
rect -22147 36968 -22127 37032
rect -28426 36952 -22127 36968
rect -28426 36888 -22211 36952
rect -22147 36888 -22127 36952
rect -28426 36872 -22127 36888
rect -28426 36808 -22211 36872
rect -22147 36808 -22127 36872
rect -28426 36792 -22127 36808
rect -28426 36728 -22211 36792
rect -22147 36728 -22127 36792
rect -28426 36712 -22127 36728
rect -28426 36648 -22211 36712
rect -22147 36648 -22127 36712
rect -28426 36632 -22127 36648
rect -28426 36568 -22211 36632
rect -22147 36568 -22127 36632
rect -28426 36552 -22127 36568
rect -28426 36488 -22211 36552
rect -22147 36488 -22127 36552
rect -28426 36472 -22127 36488
rect -28426 36408 -22211 36472
rect -22147 36408 -22127 36472
rect -28426 36392 -22127 36408
rect -28426 36328 -22211 36392
rect -22147 36328 -22127 36392
rect -28426 36312 -22127 36328
rect -28426 36248 -22211 36312
rect -22147 36248 -22127 36312
rect -28426 36232 -22127 36248
rect -28426 36168 -22211 36232
rect -22147 36168 -22127 36232
rect -28426 36152 -22127 36168
rect -28426 36088 -22211 36152
rect -22147 36088 -22127 36152
rect -28426 36072 -22127 36088
rect -28426 36008 -22211 36072
rect -22147 36008 -22127 36072
rect -28426 35992 -22127 36008
rect -28426 35928 -22211 35992
rect -22147 35928 -22127 35992
rect -28426 35912 -22127 35928
rect -28426 35848 -22211 35912
rect -22147 35848 -22127 35912
rect -28426 35832 -22127 35848
rect -28426 35768 -22211 35832
rect -22147 35768 -22127 35832
rect -28426 35752 -22127 35768
rect -28426 35688 -22211 35752
rect -22147 35688 -22127 35752
rect -28426 35672 -22127 35688
rect -28426 35608 -22211 35672
rect -22147 35608 -22127 35672
rect -28426 35592 -22127 35608
rect -28426 35528 -22211 35592
rect -22147 35528 -22127 35592
rect -28426 35512 -22127 35528
rect -28426 35448 -22211 35512
rect -22147 35448 -22127 35512
rect -28426 35432 -22127 35448
rect -28426 35368 -22211 35432
rect -22147 35368 -22127 35432
rect -28426 35352 -22127 35368
rect -28426 35288 -22211 35352
rect -22147 35288 -22127 35352
rect -28426 35272 -22127 35288
rect -28426 35208 -22211 35272
rect -22147 35208 -22127 35272
rect -28426 35192 -22127 35208
rect -28426 35128 -22211 35192
rect -22147 35128 -22127 35192
rect -28426 35112 -22127 35128
rect -28426 35048 -22211 35112
rect -22147 35048 -22127 35112
rect -28426 35032 -22127 35048
rect -28426 34968 -22211 35032
rect -22147 34968 -22127 35032
rect -28426 34952 -22127 34968
rect -28426 34888 -22211 34952
rect -22147 34888 -22127 34952
rect -28426 34872 -22127 34888
rect -28426 34808 -22211 34872
rect -22147 34808 -22127 34872
rect -28426 34792 -22127 34808
rect -28426 34728 -22211 34792
rect -22147 34728 -22127 34792
rect -28426 34700 -22127 34728
rect -22107 40872 -15808 40900
rect -22107 40808 -15892 40872
rect -15828 40808 -15808 40872
rect -22107 40792 -15808 40808
rect -22107 40728 -15892 40792
rect -15828 40728 -15808 40792
rect -22107 40712 -15808 40728
rect -22107 40648 -15892 40712
rect -15828 40648 -15808 40712
rect -22107 40632 -15808 40648
rect -22107 40568 -15892 40632
rect -15828 40568 -15808 40632
rect -22107 40552 -15808 40568
rect -22107 40488 -15892 40552
rect -15828 40488 -15808 40552
rect -22107 40472 -15808 40488
rect -22107 40408 -15892 40472
rect -15828 40408 -15808 40472
rect -22107 40392 -15808 40408
rect -22107 40328 -15892 40392
rect -15828 40328 -15808 40392
rect -22107 40312 -15808 40328
rect -22107 40248 -15892 40312
rect -15828 40248 -15808 40312
rect -22107 40232 -15808 40248
rect -22107 40168 -15892 40232
rect -15828 40168 -15808 40232
rect -22107 40152 -15808 40168
rect -22107 40088 -15892 40152
rect -15828 40088 -15808 40152
rect -22107 40072 -15808 40088
rect -22107 40008 -15892 40072
rect -15828 40008 -15808 40072
rect -22107 39992 -15808 40008
rect -22107 39928 -15892 39992
rect -15828 39928 -15808 39992
rect -22107 39912 -15808 39928
rect -22107 39848 -15892 39912
rect -15828 39848 -15808 39912
rect -22107 39832 -15808 39848
rect -22107 39768 -15892 39832
rect -15828 39768 -15808 39832
rect -22107 39752 -15808 39768
rect -22107 39688 -15892 39752
rect -15828 39688 -15808 39752
rect -22107 39672 -15808 39688
rect -22107 39608 -15892 39672
rect -15828 39608 -15808 39672
rect -22107 39592 -15808 39608
rect -22107 39528 -15892 39592
rect -15828 39528 -15808 39592
rect -22107 39512 -15808 39528
rect -22107 39448 -15892 39512
rect -15828 39448 -15808 39512
rect -22107 39432 -15808 39448
rect -22107 39368 -15892 39432
rect -15828 39368 -15808 39432
rect -22107 39352 -15808 39368
rect -22107 39288 -15892 39352
rect -15828 39288 -15808 39352
rect -22107 39272 -15808 39288
rect -22107 39208 -15892 39272
rect -15828 39208 -15808 39272
rect -22107 39192 -15808 39208
rect -22107 39128 -15892 39192
rect -15828 39128 -15808 39192
rect -22107 39112 -15808 39128
rect -22107 39048 -15892 39112
rect -15828 39048 -15808 39112
rect -22107 39032 -15808 39048
rect -22107 38968 -15892 39032
rect -15828 38968 -15808 39032
rect -22107 38952 -15808 38968
rect -22107 38888 -15892 38952
rect -15828 38888 -15808 38952
rect -22107 38872 -15808 38888
rect -22107 38808 -15892 38872
rect -15828 38808 -15808 38872
rect -22107 38792 -15808 38808
rect -22107 38728 -15892 38792
rect -15828 38728 -15808 38792
rect -22107 38712 -15808 38728
rect -22107 38648 -15892 38712
rect -15828 38648 -15808 38712
rect -22107 38632 -15808 38648
rect -22107 38568 -15892 38632
rect -15828 38568 -15808 38632
rect -22107 38552 -15808 38568
rect -22107 38488 -15892 38552
rect -15828 38488 -15808 38552
rect -22107 38472 -15808 38488
rect -22107 38408 -15892 38472
rect -15828 38408 -15808 38472
rect -22107 38392 -15808 38408
rect -22107 38328 -15892 38392
rect -15828 38328 -15808 38392
rect -22107 38312 -15808 38328
rect -22107 38248 -15892 38312
rect -15828 38248 -15808 38312
rect -22107 38232 -15808 38248
rect -22107 38168 -15892 38232
rect -15828 38168 -15808 38232
rect -22107 38152 -15808 38168
rect -22107 38088 -15892 38152
rect -15828 38088 -15808 38152
rect -22107 38072 -15808 38088
rect -22107 38008 -15892 38072
rect -15828 38008 -15808 38072
rect -22107 37992 -15808 38008
rect -22107 37928 -15892 37992
rect -15828 37928 -15808 37992
rect -22107 37912 -15808 37928
rect -22107 37848 -15892 37912
rect -15828 37848 -15808 37912
rect -22107 37832 -15808 37848
rect -22107 37768 -15892 37832
rect -15828 37768 -15808 37832
rect -22107 37752 -15808 37768
rect -22107 37688 -15892 37752
rect -15828 37688 -15808 37752
rect -22107 37672 -15808 37688
rect -22107 37608 -15892 37672
rect -15828 37608 -15808 37672
rect -22107 37592 -15808 37608
rect -22107 37528 -15892 37592
rect -15828 37528 -15808 37592
rect -22107 37512 -15808 37528
rect -22107 37448 -15892 37512
rect -15828 37448 -15808 37512
rect -22107 37432 -15808 37448
rect -22107 37368 -15892 37432
rect -15828 37368 -15808 37432
rect -22107 37352 -15808 37368
rect -22107 37288 -15892 37352
rect -15828 37288 -15808 37352
rect -22107 37272 -15808 37288
rect -22107 37208 -15892 37272
rect -15828 37208 -15808 37272
rect -22107 37192 -15808 37208
rect -22107 37128 -15892 37192
rect -15828 37128 -15808 37192
rect -22107 37112 -15808 37128
rect -22107 37048 -15892 37112
rect -15828 37048 -15808 37112
rect -22107 37032 -15808 37048
rect -22107 36968 -15892 37032
rect -15828 36968 -15808 37032
rect -22107 36952 -15808 36968
rect -22107 36888 -15892 36952
rect -15828 36888 -15808 36952
rect -22107 36872 -15808 36888
rect -22107 36808 -15892 36872
rect -15828 36808 -15808 36872
rect -22107 36792 -15808 36808
rect -22107 36728 -15892 36792
rect -15828 36728 -15808 36792
rect -22107 36712 -15808 36728
rect -22107 36648 -15892 36712
rect -15828 36648 -15808 36712
rect -22107 36632 -15808 36648
rect -22107 36568 -15892 36632
rect -15828 36568 -15808 36632
rect -22107 36552 -15808 36568
rect -22107 36488 -15892 36552
rect -15828 36488 -15808 36552
rect -22107 36472 -15808 36488
rect -22107 36408 -15892 36472
rect -15828 36408 -15808 36472
rect -22107 36392 -15808 36408
rect -22107 36328 -15892 36392
rect -15828 36328 -15808 36392
rect -22107 36312 -15808 36328
rect -22107 36248 -15892 36312
rect -15828 36248 -15808 36312
rect -22107 36232 -15808 36248
rect -22107 36168 -15892 36232
rect -15828 36168 -15808 36232
rect -22107 36152 -15808 36168
rect -22107 36088 -15892 36152
rect -15828 36088 -15808 36152
rect -22107 36072 -15808 36088
rect -22107 36008 -15892 36072
rect -15828 36008 -15808 36072
rect -22107 35992 -15808 36008
rect -22107 35928 -15892 35992
rect -15828 35928 -15808 35992
rect -22107 35912 -15808 35928
rect -22107 35848 -15892 35912
rect -15828 35848 -15808 35912
rect -22107 35832 -15808 35848
rect -22107 35768 -15892 35832
rect -15828 35768 -15808 35832
rect -22107 35752 -15808 35768
rect -22107 35688 -15892 35752
rect -15828 35688 -15808 35752
rect -22107 35672 -15808 35688
rect -22107 35608 -15892 35672
rect -15828 35608 -15808 35672
rect -22107 35592 -15808 35608
rect -22107 35528 -15892 35592
rect -15828 35528 -15808 35592
rect -22107 35512 -15808 35528
rect -22107 35448 -15892 35512
rect -15828 35448 -15808 35512
rect -22107 35432 -15808 35448
rect -22107 35368 -15892 35432
rect -15828 35368 -15808 35432
rect -22107 35352 -15808 35368
rect -22107 35288 -15892 35352
rect -15828 35288 -15808 35352
rect -22107 35272 -15808 35288
rect -22107 35208 -15892 35272
rect -15828 35208 -15808 35272
rect -22107 35192 -15808 35208
rect -22107 35128 -15892 35192
rect -15828 35128 -15808 35192
rect -22107 35112 -15808 35128
rect -22107 35048 -15892 35112
rect -15828 35048 -15808 35112
rect -22107 35032 -15808 35048
rect -22107 34968 -15892 35032
rect -15828 34968 -15808 35032
rect -22107 34952 -15808 34968
rect -22107 34888 -15892 34952
rect -15828 34888 -15808 34952
rect -22107 34872 -15808 34888
rect -22107 34808 -15892 34872
rect -15828 34808 -15808 34872
rect -22107 34792 -15808 34808
rect -22107 34728 -15892 34792
rect -15828 34728 -15808 34792
rect -22107 34700 -15808 34728
rect -15788 40872 -9489 40900
rect -15788 40808 -9573 40872
rect -9509 40808 -9489 40872
rect -15788 40792 -9489 40808
rect -15788 40728 -9573 40792
rect -9509 40728 -9489 40792
rect -15788 40712 -9489 40728
rect -15788 40648 -9573 40712
rect -9509 40648 -9489 40712
rect -15788 40632 -9489 40648
rect -15788 40568 -9573 40632
rect -9509 40568 -9489 40632
rect -15788 40552 -9489 40568
rect -15788 40488 -9573 40552
rect -9509 40488 -9489 40552
rect -15788 40472 -9489 40488
rect -15788 40408 -9573 40472
rect -9509 40408 -9489 40472
rect -15788 40392 -9489 40408
rect -15788 40328 -9573 40392
rect -9509 40328 -9489 40392
rect -15788 40312 -9489 40328
rect -15788 40248 -9573 40312
rect -9509 40248 -9489 40312
rect -15788 40232 -9489 40248
rect -15788 40168 -9573 40232
rect -9509 40168 -9489 40232
rect -15788 40152 -9489 40168
rect -15788 40088 -9573 40152
rect -9509 40088 -9489 40152
rect -15788 40072 -9489 40088
rect -15788 40008 -9573 40072
rect -9509 40008 -9489 40072
rect -15788 39992 -9489 40008
rect -15788 39928 -9573 39992
rect -9509 39928 -9489 39992
rect -15788 39912 -9489 39928
rect -15788 39848 -9573 39912
rect -9509 39848 -9489 39912
rect -15788 39832 -9489 39848
rect -15788 39768 -9573 39832
rect -9509 39768 -9489 39832
rect -15788 39752 -9489 39768
rect -15788 39688 -9573 39752
rect -9509 39688 -9489 39752
rect -15788 39672 -9489 39688
rect -15788 39608 -9573 39672
rect -9509 39608 -9489 39672
rect -15788 39592 -9489 39608
rect -15788 39528 -9573 39592
rect -9509 39528 -9489 39592
rect -15788 39512 -9489 39528
rect -15788 39448 -9573 39512
rect -9509 39448 -9489 39512
rect -15788 39432 -9489 39448
rect -15788 39368 -9573 39432
rect -9509 39368 -9489 39432
rect -15788 39352 -9489 39368
rect -15788 39288 -9573 39352
rect -9509 39288 -9489 39352
rect -15788 39272 -9489 39288
rect -15788 39208 -9573 39272
rect -9509 39208 -9489 39272
rect -15788 39192 -9489 39208
rect -15788 39128 -9573 39192
rect -9509 39128 -9489 39192
rect -15788 39112 -9489 39128
rect -15788 39048 -9573 39112
rect -9509 39048 -9489 39112
rect -15788 39032 -9489 39048
rect -15788 38968 -9573 39032
rect -9509 38968 -9489 39032
rect -15788 38952 -9489 38968
rect -15788 38888 -9573 38952
rect -9509 38888 -9489 38952
rect -15788 38872 -9489 38888
rect -15788 38808 -9573 38872
rect -9509 38808 -9489 38872
rect -15788 38792 -9489 38808
rect -15788 38728 -9573 38792
rect -9509 38728 -9489 38792
rect -15788 38712 -9489 38728
rect -15788 38648 -9573 38712
rect -9509 38648 -9489 38712
rect -15788 38632 -9489 38648
rect -15788 38568 -9573 38632
rect -9509 38568 -9489 38632
rect -15788 38552 -9489 38568
rect -15788 38488 -9573 38552
rect -9509 38488 -9489 38552
rect -15788 38472 -9489 38488
rect -15788 38408 -9573 38472
rect -9509 38408 -9489 38472
rect -15788 38392 -9489 38408
rect -15788 38328 -9573 38392
rect -9509 38328 -9489 38392
rect -15788 38312 -9489 38328
rect -15788 38248 -9573 38312
rect -9509 38248 -9489 38312
rect -15788 38232 -9489 38248
rect -15788 38168 -9573 38232
rect -9509 38168 -9489 38232
rect -15788 38152 -9489 38168
rect -15788 38088 -9573 38152
rect -9509 38088 -9489 38152
rect -15788 38072 -9489 38088
rect -15788 38008 -9573 38072
rect -9509 38008 -9489 38072
rect -15788 37992 -9489 38008
rect -15788 37928 -9573 37992
rect -9509 37928 -9489 37992
rect -15788 37912 -9489 37928
rect -15788 37848 -9573 37912
rect -9509 37848 -9489 37912
rect -15788 37832 -9489 37848
rect -15788 37768 -9573 37832
rect -9509 37768 -9489 37832
rect -15788 37752 -9489 37768
rect -15788 37688 -9573 37752
rect -9509 37688 -9489 37752
rect -15788 37672 -9489 37688
rect -15788 37608 -9573 37672
rect -9509 37608 -9489 37672
rect -15788 37592 -9489 37608
rect -15788 37528 -9573 37592
rect -9509 37528 -9489 37592
rect -15788 37512 -9489 37528
rect -15788 37448 -9573 37512
rect -9509 37448 -9489 37512
rect -15788 37432 -9489 37448
rect -15788 37368 -9573 37432
rect -9509 37368 -9489 37432
rect -15788 37352 -9489 37368
rect -15788 37288 -9573 37352
rect -9509 37288 -9489 37352
rect -15788 37272 -9489 37288
rect -15788 37208 -9573 37272
rect -9509 37208 -9489 37272
rect -15788 37192 -9489 37208
rect -15788 37128 -9573 37192
rect -9509 37128 -9489 37192
rect -15788 37112 -9489 37128
rect -15788 37048 -9573 37112
rect -9509 37048 -9489 37112
rect -15788 37032 -9489 37048
rect -15788 36968 -9573 37032
rect -9509 36968 -9489 37032
rect -15788 36952 -9489 36968
rect -15788 36888 -9573 36952
rect -9509 36888 -9489 36952
rect -15788 36872 -9489 36888
rect -15788 36808 -9573 36872
rect -9509 36808 -9489 36872
rect -15788 36792 -9489 36808
rect -15788 36728 -9573 36792
rect -9509 36728 -9489 36792
rect -15788 36712 -9489 36728
rect -15788 36648 -9573 36712
rect -9509 36648 -9489 36712
rect -15788 36632 -9489 36648
rect -15788 36568 -9573 36632
rect -9509 36568 -9489 36632
rect -15788 36552 -9489 36568
rect -15788 36488 -9573 36552
rect -9509 36488 -9489 36552
rect -15788 36472 -9489 36488
rect -15788 36408 -9573 36472
rect -9509 36408 -9489 36472
rect -15788 36392 -9489 36408
rect -15788 36328 -9573 36392
rect -9509 36328 -9489 36392
rect -15788 36312 -9489 36328
rect -15788 36248 -9573 36312
rect -9509 36248 -9489 36312
rect -15788 36232 -9489 36248
rect -15788 36168 -9573 36232
rect -9509 36168 -9489 36232
rect -15788 36152 -9489 36168
rect -15788 36088 -9573 36152
rect -9509 36088 -9489 36152
rect -15788 36072 -9489 36088
rect -15788 36008 -9573 36072
rect -9509 36008 -9489 36072
rect -15788 35992 -9489 36008
rect -15788 35928 -9573 35992
rect -9509 35928 -9489 35992
rect -15788 35912 -9489 35928
rect -15788 35848 -9573 35912
rect -9509 35848 -9489 35912
rect -15788 35832 -9489 35848
rect -15788 35768 -9573 35832
rect -9509 35768 -9489 35832
rect -15788 35752 -9489 35768
rect -15788 35688 -9573 35752
rect -9509 35688 -9489 35752
rect -15788 35672 -9489 35688
rect -15788 35608 -9573 35672
rect -9509 35608 -9489 35672
rect -15788 35592 -9489 35608
rect -15788 35528 -9573 35592
rect -9509 35528 -9489 35592
rect -15788 35512 -9489 35528
rect -15788 35448 -9573 35512
rect -9509 35448 -9489 35512
rect -15788 35432 -9489 35448
rect -15788 35368 -9573 35432
rect -9509 35368 -9489 35432
rect -15788 35352 -9489 35368
rect -15788 35288 -9573 35352
rect -9509 35288 -9489 35352
rect -15788 35272 -9489 35288
rect -15788 35208 -9573 35272
rect -9509 35208 -9489 35272
rect -15788 35192 -9489 35208
rect -15788 35128 -9573 35192
rect -9509 35128 -9489 35192
rect -15788 35112 -9489 35128
rect -15788 35048 -9573 35112
rect -9509 35048 -9489 35112
rect -15788 35032 -9489 35048
rect -15788 34968 -9573 35032
rect -9509 34968 -9489 35032
rect -15788 34952 -9489 34968
rect -15788 34888 -9573 34952
rect -9509 34888 -9489 34952
rect -15788 34872 -9489 34888
rect -15788 34808 -9573 34872
rect -9509 34808 -9489 34872
rect -15788 34792 -9489 34808
rect -15788 34728 -9573 34792
rect -9509 34728 -9489 34792
rect -15788 34700 -9489 34728
rect -9469 40872 -3170 40900
rect -9469 40808 -3254 40872
rect -3190 40808 -3170 40872
rect -9469 40792 -3170 40808
rect -9469 40728 -3254 40792
rect -3190 40728 -3170 40792
rect -9469 40712 -3170 40728
rect -9469 40648 -3254 40712
rect -3190 40648 -3170 40712
rect -9469 40632 -3170 40648
rect -9469 40568 -3254 40632
rect -3190 40568 -3170 40632
rect -9469 40552 -3170 40568
rect -9469 40488 -3254 40552
rect -3190 40488 -3170 40552
rect -9469 40472 -3170 40488
rect -9469 40408 -3254 40472
rect -3190 40408 -3170 40472
rect -9469 40392 -3170 40408
rect -9469 40328 -3254 40392
rect -3190 40328 -3170 40392
rect -9469 40312 -3170 40328
rect -9469 40248 -3254 40312
rect -3190 40248 -3170 40312
rect -9469 40232 -3170 40248
rect -9469 40168 -3254 40232
rect -3190 40168 -3170 40232
rect -9469 40152 -3170 40168
rect -9469 40088 -3254 40152
rect -3190 40088 -3170 40152
rect -9469 40072 -3170 40088
rect -9469 40008 -3254 40072
rect -3190 40008 -3170 40072
rect -9469 39992 -3170 40008
rect -9469 39928 -3254 39992
rect -3190 39928 -3170 39992
rect -9469 39912 -3170 39928
rect -9469 39848 -3254 39912
rect -3190 39848 -3170 39912
rect -9469 39832 -3170 39848
rect -9469 39768 -3254 39832
rect -3190 39768 -3170 39832
rect -9469 39752 -3170 39768
rect -9469 39688 -3254 39752
rect -3190 39688 -3170 39752
rect -9469 39672 -3170 39688
rect -9469 39608 -3254 39672
rect -3190 39608 -3170 39672
rect -9469 39592 -3170 39608
rect -9469 39528 -3254 39592
rect -3190 39528 -3170 39592
rect -9469 39512 -3170 39528
rect -9469 39448 -3254 39512
rect -3190 39448 -3170 39512
rect -9469 39432 -3170 39448
rect -9469 39368 -3254 39432
rect -3190 39368 -3170 39432
rect -9469 39352 -3170 39368
rect -9469 39288 -3254 39352
rect -3190 39288 -3170 39352
rect -9469 39272 -3170 39288
rect -9469 39208 -3254 39272
rect -3190 39208 -3170 39272
rect -9469 39192 -3170 39208
rect -9469 39128 -3254 39192
rect -3190 39128 -3170 39192
rect -9469 39112 -3170 39128
rect -9469 39048 -3254 39112
rect -3190 39048 -3170 39112
rect -9469 39032 -3170 39048
rect -9469 38968 -3254 39032
rect -3190 38968 -3170 39032
rect -9469 38952 -3170 38968
rect -9469 38888 -3254 38952
rect -3190 38888 -3170 38952
rect -9469 38872 -3170 38888
rect -9469 38808 -3254 38872
rect -3190 38808 -3170 38872
rect -9469 38792 -3170 38808
rect -9469 38728 -3254 38792
rect -3190 38728 -3170 38792
rect -9469 38712 -3170 38728
rect -9469 38648 -3254 38712
rect -3190 38648 -3170 38712
rect -9469 38632 -3170 38648
rect -9469 38568 -3254 38632
rect -3190 38568 -3170 38632
rect -9469 38552 -3170 38568
rect -9469 38488 -3254 38552
rect -3190 38488 -3170 38552
rect -9469 38472 -3170 38488
rect -9469 38408 -3254 38472
rect -3190 38408 -3170 38472
rect -9469 38392 -3170 38408
rect -9469 38328 -3254 38392
rect -3190 38328 -3170 38392
rect -9469 38312 -3170 38328
rect -9469 38248 -3254 38312
rect -3190 38248 -3170 38312
rect -9469 38232 -3170 38248
rect -9469 38168 -3254 38232
rect -3190 38168 -3170 38232
rect -9469 38152 -3170 38168
rect -9469 38088 -3254 38152
rect -3190 38088 -3170 38152
rect -9469 38072 -3170 38088
rect -9469 38008 -3254 38072
rect -3190 38008 -3170 38072
rect -9469 37992 -3170 38008
rect -9469 37928 -3254 37992
rect -3190 37928 -3170 37992
rect -9469 37912 -3170 37928
rect -9469 37848 -3254 37912
rect -3190 37848 -3170 37912
rect -9469 37832 -3170 37848
rect -9469 37768 -3254 37832
rect -3190 37768 -3170 37832
rect -9469 37752 -3170 37768
rect -9469 37688 -3254 37752
rect -3190 37688 -3170 37752
rect -9469 37672 -3170 37688
rect -9469 37608 -3254 37672
rect -3190 37608 -3170 37672
rect -9469 37592 -3170 37608
rect -9469 37528 -3254 37592
rect -3190 37528 -3170 37592
rect -9469 37512 -3170 37528
rect -9469 37448 -3254 37512
rect -3190 37448 -3170 37512
rect -9469 37432 -3170 37448
rect -9469 37368 -3254 37432
rect -3190 37368 -3170 37432
rect -9469 37352 -3170 37368
rect -9469 37288 -3254 37352
rect -3190 37288 -3170 37352
rect -9469 37272 -3170 37288
rect -9469 37208 -3254 37272
rect -3190 37208 -3170 37272
rect -9469 37192 -3170 37208
rect -9469 37128 -3254 37192
rect -3190 37128 -3170 37192
rect -9469 37112 -3170 37128
rect -9469 37048 -3254 37112
rect -3190 37048 -3170 37112
rect -9469 37032 -3170 37048
rect -9469 36968 -3254 37032
rect -3190 36968 -3170 37032
rect -9469 36952 -3170 36968
rect -9469 36888 -3254 36952
rect -3190 36888 -3170 36952
rect -9469 36872 -3170 36888
rect -9469 36808 -3254 36872
rect -3190 36808 -3170 36872
rect -9469 36792 -3170 36808
rect -9469 36728 -3254 36792
rect -3190 36728 -3170 36792
rect -9469 36712 -3170 36728
rect -9469 36648 -3254 36712
rect -3190 36648 -3170 36712
rect -9469 36632 -3170 36648
rect -9469 36568 -3254 36632
rect -3190 36568 -3170 36632
rect -9469 36552 -3170 36568
rect -9469 36488 -3254 36552
rect -3190 36488 -3170 36552
rect -9469 36472 -3170 36488
rect -9469 36408 -3254 36472
rect -3190 36408 -3170 36472
rect -9469 36392 -3170 36408
rect -9469 36328 -3254 36392
rect -3190 36328 -3170 36392
rect -9469 36312 -3170 36328
rect -9469 36248 -3254 36312
rect -3190 36248 -3170 36312
rect -9469 36232 -3170 36248
rect -9469 36168 -3254 36232
rect -3190 36168 -3170 36232
rect -9469 36152 -3170 36168
rect -9469 36088 -3254 36152
rect -3190 36088 -3170 36152
rect -9469 36072 -3170 36088
rect -9469 36008 -3254 36072
rect -3190 36008 -3170 36072
rect -9469 35992 -3170 36008
rect -9469 35928 -3254 35992
rect -3190 35928 -3170 35992
rect -9469 35912 -3170 35928
rect -9469 35848 -3254 35912
rect -3190 35848 -3170 35912
rect -9469 35832 -3170 35848
rect -9469 35768 -3254 35832
rect -3190 35768 -3170 35832
rect -9469 35752 -3170 35768
rect -9469 35688 -3254 35752
rect -3190 35688 -3170 35752
rect -9469 35672 -3170 35688
rect -9469 35608 -3254 35672
rect -3190 35608 -3170 35672
rect -9469 35592 -3170 35608
rect -9469 35528 -3254 35592
rect -3190 35528 -3170 35592
rect -9469 35512 -3170 35528
rect -9469 35448 -3254 35512
rect -3190 35448 -3170 35512
rect -9469 35432 -3170 35448
rect -9469 35368 -3254 35432
rect -3190 35368 -3170 35432
rect -9469 35352 -3170 35368
rect -9469 35288 -3254 35352
rect -3190 35288 -3170 35352
rect -9469 35272 -3170 35288
rect -9469 35208 -3254 35272
rect -3190 35208 -3170 35272
rect -9469 35192 -3170 35208
rect -9469 35128 -3254 35192
rect -3190 35128 -3170 35192
rect -9469 35112 -3170 35128
rect -9469 35048 -3254 35112
rect -3190 35048 -3170 35112
rect -9469 35032 -3170 35048
rect -9469 34968 -3254 35032
rect -3190 34968 -3170 35032
rect -9469 34952 -3170 34968
rect -9469 34888 -3254 34952
rect -3190 34888 -3170 34952
rect -9469 34872 -3170 34888
rect -9469 34808 -3254 34872
rect -3190 34808 -3170 34872
rect -9469 34792 -3170 34808
rect -9469 34728 -3254 34792
rect -3190 34728 -3170 34792
rect -9469 34700 -3170 34728
rect -3150 40872 3149 40900
rect -3150 40808 3065 40872
rect 3129 40808 3149 40872
rect -3150 40792 3149 40808
rect -3150 40728 3065 40792
rect 3129 40728 3149 40792
rect -3150 40712 3149 40728
rect -3150 40648 3065 40712
rect 3129 40648 3149 40712
rect -3150 40632 3149 40648
rect -3150 40568 3065 40632
rect 3129 40568 3149 40632
rect -3150 40552 3149 40568
rect -3150 40488 3065 40552
rect 3129 40488 3149 40552
rect -3150 40472 3149 40488
rect -3150 40408 3065 40472
rect 3129 40408 3149 40472
rect -3150 40392 3149 40408
rect -3150 40328 3065 40392
rect 3129 40328 3149 40392
rect -3150 40312 3149 40328
rect -3150 40248 3065 40312
rect 3129 40248 3149 40312
rect -3150 40232 3149 40248
rect -3150 40168 3065 40232
rect 3129 40168 3149 40232
rect -3150 40152 3149 40168
rect -3150 40088 3065 40152
rect 3129 40088 3149 40152
rect -3150 40072 3149 40088
rect -3150 40008 3065 40072
rect 3129 40008 3149 40072
rect -3150 39992 3149 40008
rect -3150 39928 3065 39992
rect 3129 39928 3149 39992
rect -3150 39912 3149 39928
rect -3150 39848 3065 39912
rect 3129 39848 3149 39912
rect -3150 39832 3149 39848
rect -3150 39768 3065 39832
rect 3129 39768 3149 39832
rect -3150 39752 3149 39768
rect -3150 39688 3065 39752
rect 3129 39688 3149 39752
rect -3150 39672 3149 39688
rect -3150 39608 3065 39672
rect 3129 39608 3149 39672
rect -3150 39592 3149 39608
rect -3150 39528 3065 39592
rect 3129 39528 3149 39592
rect -3150 39512 3149 39528
rect -3150 39448 3065 39512
rect 3129 39448 3149 39512
rect -3150 39432 3149 39448
rect -3150 39368 3065 39432
rect 3129 39368 3149 39432
rect -3150 39352 3149 39368
rect -3150 39288 3065 39352
rect 3129 39288 3149 39352
rect -3150 39272 3149 39288
rect -3150 39208 3065 39272
rect 3129 39208 3149 39272
rect -3150 39192 3149 39208
rect -3150 39128 3065 39192
rect 3129 39128 3149 39192
rect -3150 39112 3149 39128
rect -3150 39048 3065 39112
rect 3129 39048 3149 39112
rect -3150 39032 3149 39048
rect -3150 38968 3065 39032
rect 3129 38968 3149 39032
rect -3150 38952 3149 38968
rect -3150 38888 3065 38952
rect 3129 38888 3149 38952
rect -3150 38872 3149 38888
rect -3150 38808 3065 38872
rect 3129 38808 3149 38872
rect -3150 38792 3149 38808
rect -3150 38728 3065 38792
rect 3129 38728 3149 38792
rect -3150 38712 3149 38728
rect -3150 38648 3065 38712
rect 3129 38648 3149 38712
rect -3150 38632 3149 38648
rect -3150 38568 3065 38632
rect 3129 38568 3149 38632
rect -3150 38552 3149 38568
rect -3150 38488 3065 38552
rect 3129 38488 3149 38552
rect -3150 38472 3149 38488
rect -3150 38408 3065 38472
rect 3129 38408 3149 38472
rect -3150 38392 3149 38408
rect -3150 38328 3065 38392
rect 3129 38328 3149 38392
rect -3150 38312 3149 38328
rect -3150 38248 3065 38312
rect 3129 38248 3149 38312
rect -3150 38232 3149 38248
rect -3150 38168 3065 38232
rect 3129 38168 3149 38232
rect -3150 38152 3149 38168
rect -3150 38088 3065 38152
rect 3129 38088 3149 38152
rect -3150 38072 3149 38088
rect -3150 38008 3065 38072
rect 3129 38008 3149 38072
rect -3150 37992 3149 38008
rect -3150 37928 3065 37992
rect 3129 37928 3149 37992
rect -3150 37912 3149 37928
rect -3150 37848 3065 37912
rect 3129 37848 3149 37912
rect -3150 37832 3149 37848
rect -3150 37768 3065 37832
rect 3129 37768 3149 37832
rect -3150 37752 3149 37768
rect -3150 37688 3065 37752
rect 3129 37688 3149 37752
rect -3150 37672 3149 37688
rect -3150 37608 3065 37672
rect 3129 37608 3149 37672
rect -3150 37592 3149 37608
rect -3150 37528 3065 37592
rect 3129 37528 3149 37592
rect -3150 37512 3149 37528
rect -3150 37448 3065 37512
rect 3129 37448 3149 37512
rect -3150 37432 3149 37448
rect -3150 37368 3065 37432
rect 3129 37368 3149 37432
rect -3150 37352 3149 37368
rect -3150 37288 3065 37352
rect 3129 37288 3149 37352
rect -3150 37272 3149 37288
rect -3150 37208 3065 37272
rect 3129 37208 3149 37272
rect -3150 37192 3149 37208
rect -3150 37128 3065 37192
rect 3129 37128 3149 37192
rect -3150 37112 3149 37128
rect -3150 37048 3065 37112
rect 3129 37048 3149 37112
rect -3150 37032 3149 37048
rect -3150 36968 3065 37032
rect 3129 36968 3149 37032
rect -3150 36952 3149 36968
rect -3150 36888 3065 36952
rect 3129 36888 3149 36952
rect -3150 36872 3149 36888
rect -3150 36808 3065 36872
rect 3129 36808 3149 36872
rect -3150 36792 3149 36808
rect -3150 36728 3065 36792
rect 3129 36728 3149 36792
rect -3150 36712 3149 36728
rect -3150 36648 3065 36712
rect 3129 36648 3149 36712
rect -3150 36632 3149 36648
rect -3150 36568 3065 36632
rect 3129 36568 3149 36632
rect -3150 36552 3149 36568
rect -3150 36488 3065 36552
rect 3129 36488 3149 36552
rect -3150 36472 3149 36488
rect -3150 36408 3065 36472
rect 3129 36408 3149 36472
rect -3150 36392 3149 36408
rect -3150 36328 3065 36392
rect 3129 36328 3149 36392
rect -3150 36312 3149 36328
rect -3150 36248 3065 36312
rect 3129 36248 3149 36312
rect -3150 36232 3149 36248
rect -3150 36168 3065 36232
rect 3129 36168 3149 36232
rect -3150 36152 3149 36168
rect -3150 36088 3065 36152
rect 3129 36088 3149 36152
rect -3150 36072 3149 36088
rect -3150 36008 3065 36072
rect 3129 36008 3149 36072
rect -3150 35992 3149 36008
rect -3150 35928 3065 35992
rect 3129 35928 3149 35992
rect -3150 35912 3149 35928
rect -3150 35848 3065 35912
rect 3129 35848 3149 35912
rect -3150 35832 3149 35848
rect -3150 35768 3065 35832
rect 3129 35768 3149 35832
rect -3150 35752 3149 35768
rect -3150 35688 3065 35752
rect 3129 35688 3149 35752
rect -3150 35672 3149 35688
rect -3150 35608 3065 35672
rect 3129 35608 3149 35672
rect -3150 35592 3149 35608
rect -3150 35528 3065 35592
rect 3129 35528 3149 35592
rect -3150 35512 3149 35528
rect -3150 35448 3065 35512
rect 3129 35448 3149 35512
rect -3150 35432 3149 35448
rect -3150 35368 3065 35432
rect 3129 35368 3149 35432
rect -3150 35352 3149 35368
rect -3150 35288 3065 35352
rect 3129 35288 3149 35352
rect -3150 35272 3149 35288
rect -3150 35208 3065 35272
rect 3129 35208 3149 35272
rect -3150 35192 3149 35208
rect -3150 35128 3065 35192
rect 3129 35128 3149 35192
rect -3150 35112 3149 35128
rect -3150 35048 3065 35112
rect 3129 35048 3149 35112
rect -3150 35032 3149 35048
rect -3150 34968 3065 35032
rect 3129 34968 3149 35032
rect -3150 34952 3149 34968
rect -3150 34888 3065 34952
rect 3129 34888 3149 34952
rect -3150 34872 3149 34888
rect -3150 34808 3065 34872
rect 3129 34808 3149 34872
rect -3150 34792 3149 34808
rect -3150 34728 3065 34792
rect 3129 34728 3149 34792
rect -3150 34700 3149 34728
rect 3169 40872 9468 40900
rect 3169 40808 9384 40872
rect 9448 40808 9468 40872
rect 3169 40792 9468 40808
rect 3169 40728 9384 40792
rect 9448 40728 9468 40792
rect 3169 40712 9468 40728
rect 3169 40648 9384 40712
rect 9448 40648 9468 40712
rect 3169 40632 9468 40648
rect 3169 40568 9384 40632
rect 9448 40568 9468 40632
rect 3169 40552 9468 40568
rect 3169 40488 9384 40552
rect 9448 40488 9468 40552
rect 3169 40472 9468 40488
rect 3169 40408 9384 40472
rect 9448 40408 9468 40472
rect 3169 40392 9468 40408
rect 3169 40328 9384 40392
rect 9448 40328 9468 40392
rect 3169 40312 9468 40328
rect 3169 40248 9384 40312
rect 9448 40248 9468 40312
rect 3169 40232 9468 40248
rect 3169 40168 9384 40232
rect 9448 40168 9468 40232
rect 3169 40152 9468 40168
rect 3169 40088 9384 40152
rect 9448 40088 9468 40152
rect 3169 40072 9468 40088
rect 3169 40008 9384 40072
rect 9448 40008 9468 40072
rect 3169 39992 9468 40008
rect 3169 39928 9384 39992
rect 9448 39928 9468 39992
rect 3169 39912 9468 39928
rect 3169 39848 9384 39912
rect 9448 39848 9468 39912
rect 3169 39832 9468 39848
rect 3169 39768 9384 39832
rect 9448 39768 9468 39832
rect 3169 39752 9468 39768
rect 3169 39688 9384 39752
rect 9448 39688 9468 39752
rect 3169 39672 9468 39688
rect 3169 39608 9384 39672
rect 9448 39608 9468 39672
rect 3169 39592 9468 39608
rect 3169 39528 9384 39592
rect 9448 39528 9468 39592
rect 3169 39512 9468 39528
rect 3169 39448 9384 39512
rect 9448 39448 9468 39512
rect 3169 39432 9468 39448
rect 3169 39368 9384 39432
rect 9448 39368 9468 39432
rect 3169 39352 9468 39368
rect 3169 39288 9384 39352
rect 9448 39288 9468 39352
rect 3169 39272 9468 39288
rect 3169 39208 9384 39272
rect 9448 39208 9468 39272
rect 3169 39192 9468 39208
rect 3169 39128 9384 39192
rect 9448 39128 9468 39192
rect 3169 39112 9468 39128
rect 3169 39048 9384 39112
rect 9448 39048 9468 39112
rect 3169 39032 9468 39048
rect 3169 38968 9384 39032
rect 9448 38968 9468 39032
rect 3169 38952 9468 38968
rect 3169 38888 9384 38952
rect 9448 38888 9468 38952
rect 3169 38872 9468 38888
rect 3169 38808 9384 38872
rect 9448 38808 9468 38872
rect 3169 38792 9468 38808
rect 3169 38728 9384 38792
rect 9448 38728 9468 38792
rect 3169 38712 9468 38728
rect 3169 38648 9384 38712
rect 9448 38648 9468 38712
rect 3169 38632 9468 38648
rect 3169 38568 9384 38632
rect 9448 38568 9468 38632
rect 3169 38552 9468 38568
rect 3169 38488 9384 38552
rect 9448 38488 9468 38552
rect 3169 38472 9468 38488
rect 3169 38408 9384 38472
rect 9448 38408 9468 38472
rect 3169 38392 9468 38408
rect 3169 38328 9384 38392
rect 9448 38328 9468 38392
rect 3169 38312 9468 38328
rect 3169 38248 9384 38312
rect 9448 38248 9468 38312
rect 3169 38232 9468 38248
rect 3169 38168 9384 38232
rect 9448 38168 9468 38232
rect 3169 38152 9468 38168
rect 3169 38088 9384 38152
rect 9448 38088 9468 38152
rect 3169 38072 9468 38088
rect 3169 38008 9384 38072
rect 9448 38008 9468 38072
rect 3169 37992 9468 38008
rect 3169 37928 9384 37992
rect 9448 37928 9468 37992
rect 3169 37912 9468 37928
rect 3169 37848 9384 37912
rect 9448 37848 9468 37912
rect 3169 37832 9468 37848
rect 3169 37768 9384 37832
rect 9448 37768 9468 37832
rect 3169 37752 9468 37768
rect 3169 37688 9384 37752
rect 9448 37688 9468 37752
rect 3169 37672 9468 37688
rect 3169 37608 9384 37672
rect 9448 37608 9468 37672
rect 3169 37592 9468 37608
rect 3169 37528 9384 37592
rect 9448 37528 9468 37592
rect 3169 37512 9468 37528
rect 3169 37448 9384 37512
rect 9448 37448 9468 37512
rect 3169 37432 9468 37448
rect 3169 37368 9384 37432
rect 9448 37368 9468 37432
rect 3169 37352 9468 37368
rect 3169 37288 9384 37352
rect 9448 37288 9468 37352
rect 3169 37272 9468 37288
rect 3169 37208 9384 37272
rect 9448 37208 9468 37272
rect 3169 37192 9468 37208
rect 3169 37128 9384 37192
rect 9448 37128 9468 37192
rect 3169 37112 9468 37128
rect 3169 37048 9384 37112
rect 9448 37048 9468 37112
rect 3169 37032 9468 37048
rect 3169 36968 9384 37032
rect 9448 36968 9468 37032
rect 3169 36952 9468 36968
rect 3169 36888 9384 36952
rect 9448 36888 9468 36952
rect 3169 36872 9468 36888
rect 3169 36808 9384 36872
rect 9448 36808 9468 36872
rect 3169 36792 9468 36808
rect 3169 36728 9384 36792
rect 9448 36728 9468 36792
rect 3169 36712 9468 36728
rect 3169 36648 9384 36712
rect 9448 36648 9468 36712
rect 3169 36632 9468 36648
rect 3169 36568 9384 36632
rect 9448 36568 9468 36632
rect 3169 36552 9468 36568
rect 3169 36488 9384 36552
rect 9448 36488 9468 36552
rect 3169 36472 9468 36488
rect 3169 36408 9384 36472
rect 9448 36408 9468 36472
rect 3169 36392 9468 36408
rect 3169 36328 9384 36392
rect 9448 36328 9468 36392
rect 3169 36312 9468 36328
rect 3169 36248 9384 36312
rect 9448 36248 9468 36312
rect 3169 36232 9468 36248
rect 3169 36168 9384 36232
rect 9448 36168 9468 36232
rect 3169 36152 9468 36168
rect 3169 36088 9384 36152
rect 9448 36088 9468 36152
rect 3169 36072 9468 36088
rect 3169 36008 9384 36072
rect 9448 36008 9468 36072
rect 3169 35992 9468 36008
rect 3169 35928 9384 35992
rect 9448 35928 9468 35992
rect 3169 35912 9468 35928
rect 3169 35848 9384 35912
rect 9448 35848 9468 35912
rect 3169 35832 9468 35848
rect 3169 35768 9384 35832
rect 9448 35768 9468 35832
rect 3169 35752 9468 35768
rect 3169 35688 9384 35752
rect 9448 35688 9468 35752
rect 3169 35672 9468 35688
rect 3169 35608 9384 35672
rect 9448 35608 9468 35672
rect 3169 35592 9468 35608
rect 3169 35528 9384 35592
rect 9448 35528 9468 35592
rect 3169 35512 9468 35528
rect 3169 35448 9384 35512
rect 9448 35448 9468 35512
rect 3169 35432 9468 35448
rect 3169 35368 9384 35432
rect 9448 35368 9468 35432
rect 3169 35352 9468 35368
rect 3169 35288 9384 35352
rect 9448 35288 9468 35352
rect 3169 35272 9468 35288
rect 3169 35208 9384 35272
rect 9448 35208 9468 35272
rect 3169 35192 9468 35208
rect 3169 35128 9384 35192
rect 9448 35128 9468 35192
rect 3169 35112 9468 35128
rect 3169 35048 9384 35112
rect 9448 35048 9468 35112
rect 3169 35032 9468 35048
rect 3169 34968 9384 35032
rect 9448 34968 9468 35032
rect 3169 34952 9468 34968
rect 3169 34888 9384 34952
rect 9448 34888 9468 34952
rect 3169 34872 9468 34888
rect 3169 34808 9384 34872
rect 9448 34808 9468 34872
rect 3169 34792 9468 34808
rect 3169 34728 9384 34792
rect 9448 34728 9468 34792
rect 3169 34700 9468 34728
rect 9488 40872 15787 40900
rect 9488 40808 15703 40872
rect 15767 40808 15787 40872
rect 9488 40792 15787 40808
rect 9488 40728 15703 40792
rect 15767 40728 15787 40792
rect 9488 40712 15787 40728
rect 9488 40648 15703 40712
rect 15767 40648 15787 40712
rect 9488 40632 15787 40648
rect 9488 40568 15703 40632
rect 15767 40568 15787 40632
rect 9488 40552 15787 40568
rect 9488 40488 15703 40552
rect 15767 40488 15787 40552
rect 9488 40472 15787 40488
rect 9488 40408 15703 40472
rect 15767 40408 15787 40472
rect 9488 40392 15787 40408
rect 9488 40328 15703 40392
rect 15767 40328 15787 40392
rect 9488 40312 15787 40328
rect 9488 40248 15703 40312
rect 15767 40248 15787 40312
rect 9488 40232 15787 40248
rect 9488 40168 15703 40232
rect 15767 40168 15787 40232
rect 9488 40152 15787 40168
rect 9488 40088 15703 40152
rect 15767 40088 15787 40152
rect 9488 40072 15787 40088
rect 9488 40008 15703 40072
rect 15767 40008 15787 40072
rect 9488 39992 15787 40008
rect 9488 39928 15703 39992
rect 15767 39928 15787 39992
rect 9488 39912 15787 39928
rect 9488 39848 15703 39912
rect 15767 39848 15787 39912
rect 9488 39832 15787 39848
rect 9488 39768 15703 39832
rect 15767 39768 15787 39832
rect 9488 39752 15787 39768
rect 9488 39688 15703 39752
rect 15767 39688 15787 39752
rect 9488 39672 15787 39688
rect 9488 39608 15703 39672
rect 15767 39608 15787 39672
rect 9488 39592 15787 39608
rect 9488 39528 15703 39592
rect 15767 39528 15787 39592
rect 9488 39512 15787 39528
rect 9488 39448 15703 39512
rect 15767 39448 15787 39512
rect 9488 39432 15787 39448
rect 9488 39368 15703 39432
rect 15767 39368 15787 39432
rect 9488 39352 15787 39368
rect 9488 39288 15703 39352
rect 15767 39288 15787 39352
rect 9488 39272 15787 39288
rect 9488 39208 15703 39272
rect 15767 39208 15787 39272
rect 9488 39192 15787 39208
rect 9488 39128 15703 39192
rect 15767 39128 15787 39192
rect 9488 39112 15787 39128
rect 9488 39048 15703 39112
rect 15767 39048 15787 39112
rect 9488 39032 15787 39048
rect 9488 38968 15703 39032
rect 15767 38968 15787 39032
rect 9488 38952 15787 38968
rect 9488 38888 15703 38952
rect 15767 38888 15787 38952
rect 9488 38872 15787 38888
rect 9488 38808 15703 38872
rect 15767 38808 15787 38872
rect 9488 38792 15787 38808
rect 9488 38728 15703 38792
rect 15767 38728 15787 38792
rect 9488 38712 15787 38728
rect 9488 38648 15703 38712
rect 15767 38648 15787 38712
rect 9488 38632 15787 38648
rect 9488 38568 15703 38632
rect 15767 38568 15787 38632
rect 9488 38552 15787 38568
rect 9488 38488 15703 38552
rect 15767 38488 15787 38552
rect 9488 38472 15787 38488
rect 9488 38408 15703 38472
rect 15767 38408 15787 38472
rect 9488 38392 15787 38408
rect 9488 38328 15703 38392
rect 15767 38328 15787 38392
rect 9488 38312 15787 38328
rect 9488 38248 15703 38312
rect 15767 38248 15787 38312
rect 9488 38232 15787 38248
rect 9488 38168 15703 38232
rect 15767 38168 15787 38232
rect 9488 38152 15787 38168
rect 9488 38088 15703 38152
rect 15767 38088 15787 38152
rect 9488 38072 15787 38088
rect 9488 38008 15703 38072
rect 15767 38008 15787 38072
rect 9488 37992 15787 38008
rect 9488 37928 15703 37992
rect 15767 37928 15787 37992
rect 9488 37912 15787 37928
rect 9488 37848 15703 37912
rect 15767 37848 15787 37912
rect 9488 37832 15787 37848
rect 9488 37768 15703 37832
rect 15767 37768 15787 37832
rect 9488 37752 15787 37768
rect 9488 37688 15703 37752
rect 15767 37688 15787 37752
rect 9488 37672 15787 37688
rect 9488 37608 15703 37672
rect 15767 37608 15787 37672
rect 9488 37592 15787 37608
rect 9488 37528 15703 37592
rect 15767 37528 15787 37592
rect 9488 37512 15787 37528
rect 9488 37448 15703 37512
rect 15767 37448 15787 37512
rect 9488 37432 15787 37448
rect 9488 37368 15703 37432
rect 15767 37368 15787 37432
rect 9488 37352 15787 37368
rect 9488 37288 15703 37352
rect 15767 37288 15787 37352
rect 9488 37272 15787 37288
rect 9488 37208 15703 37272
rect 15767 37208 15787 37272
rect 9488 37192 15787 37208
rect 9488 37128 15703 37192
rect 15767 37128 15787 37192
rect 9488 37112 15787 37128
rect 9488 37048 15703 37112
rect 15767 37048 15787 37112
rect 9488 37032 15787 37048
rect 9488 36968 15703 37032
rect 15767 36968 15787 37032
rect 9488 36952 15787 36968
rect 9488 36888 15703 36952
rect 15767 36888 15787 36952
rect 9488 36872 15787 36888
rect 9488 36808 15703 36872
rect 15767 36808 15787 36872
rect 9488 36792 15787 36808
rect 9488 36728 15703 36792
rect 15767 36728 15787 36792
rect 9488 36712 15787 36728
rect 9488 36648 15703 36712
rect 15767 36648 15787 36712
rect 9488 36632 15787 36648
rect 9488 36568 15703 36632
rect 15767 36568 15787 36632
rect 9488 36552 15787 36568
rect 9488 36488 15703 36552
rect 15767 36488 15787 36552
rect 9488 36472 15787 36488
rect 9488 36408 15703 36472
rect 15767 36408 15787 36472
rect 9488 36392 15787 36408
rect 9488 36328 15703 36392
rect 15767 36328 15787 36392
rect 9488 36312 15787 36328
rect 9488 36248 15703 36312
rect 15767 36248 15787 36312
rect 9488 36232 15787 36248
rect 9488 36168 15703 36232
rect 15767 36168 15787 36232
rect 9488 36152 15787 36168
rect 9488 36088 15703 36152
rect 15767 36088 15787 36152
rect 9488 36072 15787 36088
rect 9488 36008 15703 36072
rect 15767 36008 15787 36072
rect 9488 35992 15787 36008
rect 9488 35928 15703 35992
rect 15767 35928 15787 35992
rect 9488 35912 15787 35928
rect 9488 35848 15703 35912
rect 15767 35848 15787 35912
rect 9488 35832 15787 35848
rect 9488 35768 15703 35832
rect 15767 35768 15787 35832
rect 9488 35752 15787 35768
rect 9488 35688 15703 35752
rect 15767 35688 15787 35752
rect 9488 35672 15787 35688
rect 9488 35608 15703 35672
rect 15767 35608 15787 35672
rect 9488 35592 15787 35608
rect 9488 35528 15703 35592
rect 15767 35528 15787 35592
rect 9488 35512 15787 35528
rect 9488 35448 15703 35512
rect 15767 35448 15787 35512
rect 9488 35432 15787 35448
rect 9488 35368 15703 35432
rect 15767 35368 15787 35432
rect 9488 35352 15787 35368
rect 9488 35288 15703 35352
rect 15767 35288 15787 35352
rect 9488 35272 15787 35288
rect 9488 35208 15703 35272
rect 15767 35208 15787 35272
rect 9488 35192 15787 35208
rect 9488 35128 15703 35192
rect 15767 35128 15787 35192
rect 9488 35112 15787 35128
rect 9488 35048 15703 35112
rect 15767 35048 15787 35112
rect 9488 35032 15787 35048
rect 9488 34968 15703 35032
rect 15767 34968 15787 35032
rect 9488 34952 15787 34968
rect 9488 34888 15703 34952
rect 15767 34888 15787 34952
rect 9488 34872 15787 34888
rect 9488 34808 15703 34872
rect 15767 34808 15787 34872
rect 9488 34792 15787 34808
rect 9488 34728 15703 34792
rect 15767 34728 15787 34792
rect 9488 34700 15787 34728
rect 15807 40872 22106 40900
rect 15807 40808 22022 40872
rect 22086 40808 22106 40872
rect 15807 40792 22106 40808
rect 15807 40728 22022 40792
rect 22086 40728 22106 40792
rect 15807 40712 22106 40728
rect 15807 40648 22022 40712
rect 22086 40648 22106 40712
rect 15807 40632 22106 40648
rect 15807 40568 22022 40632
rect 22086 40568 22106 40632
rect 15807 40552 22106 40568
rect 15807 40488 22022 40552
rect 22086 40488 22106 40552
rect 15807 40472 22106 40488
rect 15807 40408 22022 40472
rect 22086 40408 22106 40472
rect 15807 40392 22106 40408
rect 15807 40328 22022 40392
rect 22086 40328 22106 40392
rect 15807 40312 22106 40328
rect 15807 40248 22022 40312
rect 22086 40248 22106 40312
rect 15807 40232 22106 40248
rect 15807 40168 22022 40232
rect 22086 40168 22106 40232
rect 15807 40152 22106 40168
rect 15807 40088 22022 40152
rect 22086 40088 22106 40152
rect 15807 40072 22106 40088
rect 15807 40008 22022 40072
rect 22086 40008 22106 40072
rect 15807 39992 22106 40008
rect 15807 39928 22022 39992
rect 22086 39928 22106 39992
rect 15807 39912 22106 39928
rect 15807 39848 22022 39912
rect 22086 39848 22106 39912
rect 15807 39832 22106 39848
rect 15807 39768 22022 39832
rect 22086 39768 22106 39832
rect 15807 39752 22106 39768
rect 15807 39688 22022 39752
rect 22086 39688 22106 39752
rect 15807 39672 22106 39688
rect 15807 39608 22022 39672
rect 22086 39608 22106 39672
rect 15807 39592 22106 39608
rect 15807 39528 22022 39592
rect 22086 39528 22106 39592
rect 15807 39512 22106 39528
rect 15807 39448 22022 39512
rect 22086 39448 22106 39512
rect 15807 39432 22106 39448
rect 15807 39368 22022 39432
rect 22086 39368 22106 39432
rect 15807 39352 22106 39368
rect 15807 39288 22022 39352
rect 22086 39288 22106 39352
rect 15807 39272 22106 39288
rect 15807 39208 22022 39272
rect 22086 39208 22106 39272
rect 15807 39192 22106 39208
rect 15807 39128 22022 39192
rect 22086 39128 22106 39192
rect 15807 39112 22106 39128
rect 15807 39048 22022 39112
rect 22086 39048 22106 39112
rect 15807 39032 22106 39048
rect 15807 38968 22022 39032
rect 22086 38968 22106 39032
rect 15807 38952 22106 38968
rect 15807 38888 22022 38952
rect 22086 38888 22106 38952
rect 15807 38872 22106 38888
rect 15807 38808 22022 38872
rect 22086 38808 22106 38872
rect 15807 38792 22106 38808
rect 15807 38728 22022 38792
rect 22086 38728 22106 38792
rect 15807 38712 22106 38728
rect 15807 38648 22022 38712
rect 22086 38648 22106 38712
rect 15807 38632 22106 38648
rect 15807 38568 22022 38632
rect 22086 38568 22106 38632
rect 15807 38552 22106 38568
rect 15807 38488 22022 38552
rect 22086 38488 22106 38552
rect 15807 38472 22106 38488
rect 15807 38408 22022 38472
rect 22086 38408 22106 38472
rect 15807 38392 22106 38408
rect 15807 38328 22022 38392
rect 22086 38328 22106 38392
rect 15807 38312 22106 38328
rect 15807 38248 22022 38312
rect 22086 38248 22106 38312
rect 15807 38232 22106 38248
rect 15807 38168 22022 38232
rect 22086 38168 22106 38232
rect 15807 38152 22106 38168
rect 15807 38088 22022 38152
rect 22086 38088 22106 38152
rect 15807 38072 22106 38088
rect 15807 38008 22022 38072
rect 22086 38008 22106 38072
rect 15807 37992 22106 38008
rect 15807 37928 22022 37992
rect 22086 37928 22106 37992
rect 15807 37912 22106 37928
rect 15807 37848 22022 37912
rect 22086 37848 22106 37912
rect 15807 37832 22106 37848
rect 15807 37768 22022 37832
rect 22086 37768 22106 37832
rect 15807 37752 22106 37768
rect 15807 37688 22022 37752
rect 22086 37688 22106 37752
rect 15807 37672 22106 37688
rect 15807 37608 22022 37672
rect 22086 37608 22106 37672
rect 15807 37592 22106 37608
rect 15807 37528 22022 37592
rect 22086 37528 22106 37592
rect 15807 37512 22106 37528
rect 15807 37448 22022 37512
rect 22086 37448 22106 37512
rect 15807 37432 22106 37448
rect 15807 37368 22022 37432
rect 22086 37368 22106 37432
rect 15807 37352 22106 37368
rect 15807 37288 22022 37352
rect 22086 37288 22106 37352
rect 15807 37272 22106 37288
rect 15807 37208 22022 37272
rect 22086 37208 22106 37272
rect 15807 37192 22106 37208
rect 15807 37128 22022 37192
rect 22086 37128 22106 37192
rect 15807 37112 22106 37128
rect 15807 37048 22022 37112
rect 22086 37048 22106 37112
rect 15807 37032 22106 37048
rect 15807 36968 22022 37032
rect 22086 36968 22106 37032
rect 15807 36952 22106 36968
rect 15807 36888 22022 36952
rect 22086 36888 22106 36952
rect 15807 36872 22106 36888
rect 15807 36808 22022 36872
rect 22086 36808 22106 36872
rect 15807 36792 22106 36808
rect 15807 36728 22022 36792
rect 22086 36728 22106 36792
rect 15807 36712 22106 36728
rect 15807 36648 22022 36712
rect 22086 36648 22106 36712
rect 15807 36632 22106 36648
rect 15807 36568 22022 36632
rect 22086 36568 22106 36632
rect 15807 36552 22106 36568
rect 15807 36488 22022 36552
rect 22086 36488 22106 36552
rect 15807 36472 22106 36488
rect 15807 36408 22022 36472
rect 22086 36408 22106 36472
rect 15807 36392 22106 36408
rect 15807 36328 22022 36392
rect 22086 36328 22106 36392
rect 15807 36312 22106 36328
rect 15807 36248 22022 36312
rect 22086 36248 22106 36312
rect 15807 36232 22106 36248
rect 15807 36168 22022 36232
rect 22086 36168 22106 36232
rect 15807 36152 22106 36168
rect 15807 36088 22022 36152
rect 22086 36088 22106 36152
rect 15807 36072 22106 36088
rect 15807 36008 22022 36072
rect 22086 36008 22106 36072
rect 15807 35992 22106 36008
rect 15807 35928 22022 35992
rect 22086 35928 22106 35992
rect 15807 35912 22106 35928
rect 15807 35848 22022 35912
rect 22086 35848 22106 35912
rect 15807 35832 22106 35848
rect 15807 35768 22022 35832
rect 22086 35768 22106 35832
rect 15807 35752 22106 35768
rect 15807 35688 22022 35752
rect 22086 35688 22106 35752
rect 15807 35672 22106 35688
rect 15807 35608 22022 35672
rect 22086 35608 22106 35672
rect 15807 35592 22106 35608
rect 15807 35528 22022 35592
rect 22086 35528 22106 35592
rect 15807 35512 22106 35528
rect 15807 35448 22022 35512
rect 22086 35448 22106 35512
rect 15807 35432 22106 35448
rect 15807 35368 22022 35432
rect 22086 35368 22106 35432
rect 15807 35352 22106 35368
rect 15807 35288 22022 35352
rect 22086 35288 22106 35352
rect 15807 35272 22106 35288
rect 15807 35208 22022 35272
rect 22086 35208 22106 35272
rect 15807 35192 22106 35208
rect 15807 35128 22022 35192
rect 22086 35128 22106 35192
rect 15807 35112 22106 35128
rect 15807 35048 22022 35112
rect 22086 35048 22106 35112
rect 15807 35032 22106 35048
rect 15807 34968 22022 35032
rect 22086 34968 22106 35032
rect 15807 34952 22106 34968
rect 15807 34888 22022 34952
rect 22086 34888 22106 34952
rect 15807 34872 22106 34888
rect 15807 34808 22022 34872
rect 22086 34808 22106 34872
rect 15807 34792 22106 34808
rect 15807 34728 22022 34792
rect 22086 34728 22106 34792
rect 15807 34700 22106 34728
rect 22126 40872 28425 40900
rect 22126 40808 28341 40872
rect 28405 40808 28425 40872
rect 22126 40792 28425 40808
rect 22126 40728 28341 40792
rect 28405 40728 28425 40792
rect 22126 40712 28425 40728
rect 22126 40648 28341 40712
rect 28405 40648 28425 40712
rect 22126 40632 28425 40648
rect 22126 40568 28341 40632
rect 28405 40568 28425 40632
rect 22126 40552 28425 40568
rect 22126 40488 28341 40552
rect 28405 40488 28425 40552
rect 22126 40472 28425 40488
rect 22126 40408 28341 40472
rect 28405 40408 28425 40472
rect 22126 40392 28425 40408
rect 22126 40328 28341 40392
rect 28405 40328 28425 40392
rect 22126 40312 28425 40328
rect 22126 40248 28341 40312
rect 28405 40248 28425 40312
rect 22126 40232 28425 40248
rect 22126 40168 28341 40232
rect 28405 40168 28425 40232
rect 22126 40152 28425 40168
rect 22126 40088 28341 40152
rect 28405 40088 28425 40152
rect 22126 40072 28425 40088
rect 22126 40008 28341 40072
rect 28405 40008 28425 40072
rect 22126 39992 28425 40008
rect 22126 39928 28341 39992
rect 28405 39928 28425 39992
rect 22126 39912 28425 39928
rect 22126 39848 28341 39912
rect 28405 39848 28425 39912
rect 22126 39832 28425 39848
rect 22126 39768 28341 39832
rect 28405 39768 28425 39832
rect 22126 39752 28425 39768
rect 22126 39688 28341 39752
rect 28405 39688 28425 39752
rect 22126 39672 28425 39688
rect 22126 39608 28341 39672
rect 28405 39608 28425 39672
rect 22126 39592 28425 39608
rect 22126 39528 28341 39592
rect 28405 39528 28425 39592
rect 22126 39512 28425 39528
rect 22126 39448 28341 39512
rect 28405 39448 28425 39512
rect 22126 39432 28425 39448
rect 22126 39368 28341 39432
rect 28405 39368 28425 39432
rect 22126 39352 28425 39368
rect 22126 39288 28341 39352
rect 28405 39288 28425 39352
rect 22126 39272 28425 39288
rect 22126 39208 28341 39272
rect 28405 39208 28425 39272
rect 22126 39192 28425 39208
rect 22126 39128 28341 39192
rect 28405 39128 28425 39192
rect 22126 39112 28425 39128
rect 22126 39048 28341 39112
rect 28405 39048 28425 39112
rect 22126 39032 28425 39048
rect 22126 38968 28341 39032
rect 28405 38968 28425 39032
rect 22126 38952 28425 38968
rect 22126 38888 28341 38952
rect 28405 38888 28425 38952
rect 22126 38872 28425 38888
rect 22126 38808 28341 38872
rect 28405 38808 28425 38872
rect 22126 38792 28425 38808
rect 22126 38728 28341 38792
rect 28405 38728 28425 38792
rect 22126 38712 28425 38728
rect 22126 38648 28341 38712
rect 28405 38648 28425 38712
rect 22126 38632 28425 38648
rect 22126 38568 28341 38632
rect 28405 38568 28425 38632
rect 22126 38552 28425 38568
rect 22126 38488 28341 38552
rect 28405 38488 28425 38552
rect 22126 38472 28425 38488
rect 22126 38408 28341 38472
rect 28405 38408 28425 38472
rect 22126 38392 28425 38408
rect 22126 38328 28341 38392
rect 28405 38328 28425 38392
rect 22126 38312 28425 38328
rect 22126 38248 28341 38312
rect 28405 38248 28425 38312
rect 22126 38232 28425 38248
rect 22126 38168 28341 38232
rect 28405 38168 28425 38232
rect 22126 38152 28425 38168
rect 22126 38088 28341 38152
rect 28405 38088 28425 38152
rect 22126 38072 28425 38088
rect 22126 38008 28341 38072
rect 28405 38008 28425 38072
rect 22126 37992 28425 38008
rect 22126 37928 28341 37992
rect 28405 37928 28425 37992
rect 22126 37912 28425 37928
rect 22126 37848 28341 37912
rect 28405 37848 28425 37912
rect 22126 37832 28425 37848
rect 22126 37768 28341 37832
rect 28405 37768 28425 37832
rect 22126 37752 28425 37768
rect 22126 37688 28341 37752
rect 28405 37688 28425 37752
rect 22126 37672 28425 37688
rect 22126 37608 28341 37672
rect 28405 37608 28425 37672
rect 22126 37592 28425 37608
rect 22126 37528 28341 37592
rect 28405 37528 28425 37592
rect 22126 37512 28425 37528
rect 22126 37448 28341 37512
rect 28405 37448 28425 37512
rect 22126 37432 28425 37448
rect 22126 37368 28341 37432
rect 28405 37368 28425 37432
rect 22126 37352 28425 37368
rect 22126 37288 28341 37352
rect 28405 37288 28425 37352
rect 22126 37272 28425 37288
rect 22126 37208 28341 37272
rect 28405 37208 28425 37272
rect 22126 37192 28425 37208
rect 22126 37128 28341 37192
rect 28405 37128 28425 37192
rect 22126 37112 28425 37128
rect 22126 37048 28341 37112
rect 28405 37048 28425 37112
rect 22126 37032 28425 37048
rect 22126 36968 28341 37032
rect 28405 36968 28425 37032
rect 22126 36952 28425 36968
rect 22126 36888 28341 36952
rect 28405 36888 28425 36952
rect 22126 36872 28425 36888
rect 22126 36808 28341 36872
rect 28405 36808 28425 36872
rect 22126 36792 28425 36808
rect 22126 36728 28341 36792
rect 28405 36728 28425 36792
rect 22126 36712 28425 36728
rect 22126 36648 28341 36712
rect 28405 36648 28425 36712
rect 22126 36632 28425 36648
rect 22126 36568 28341 36632
rect 28405 36568 28425 36632
rect 22126 36552 28425 36568
rect 22126 36488 28341 36552
rect 28405 36488 28425 36552
rect 22126 36472 28425 36488
rect 22126 36408 28341 36472
rect 28405 36408 28425 36472
rect 22126 36392 28425 36408
rect 22126 36328 28341 36392
rect 28405 36328 28425 36392
rect 22126 36312 28425 36328
rect 22126 36248 28341 36312
rect 28405 36248 28425 36312
rect 22126 36232 28425 36248
rect 22126 36168 28341 36232
rect 28405 36168 28425 36232
rect 22126 36152 28425 36168
rect 22126 36088 28341 36152
rect 28405 36088 28425 36152
rect 22126 36072 28425 36088
rect 22126 36008 28341 36072
rect 28405 36008 28425 36072
rect 22126 35992 28425 36008
rect 22126 35928 28341 35992
rect 28405 35928 28425 35992
rect 22126 35912 28425 35928
rect 22126 35848 28341 35912
rect 28405 35848 28425 35912
rect 22126 35832 28425 35848
rect 22126 35768 28341 35832
rect 28405 35768 28425 35832
rect 22126 35752 28425 35768
rect 22126 35688 28341 35752
rect 28405 35688 28425 35752
rect 22126 35672 28425 35688
rect 22126 35608 28341 35672
rect 28405 35608 28425 35672
rect 22126 35592 28425 35608
rect 22126 35528 28341 35592
rect 28405 35528 28425 35592
rect 22126 35512 28425 35528
rect 22126 35448 28341 35512
rect 28405 35448 28425 35512
rect 22126 35432 28425 35448
rect 22126 35368 28341 35432
rect 28405 35368 28425 35432
rect 22126 35352 28425 35368
rect 22126 35288 28341 35352
rect 28405 35288 28425 35352
rect 22126 35272 28425 35288
rect 22126 35208 28341 35272
rect 28405 35208 28425 35272
rect 22126 35192 28425 35208
rect 22126 35128 28341 35192
rect 28405 35128 28425 35192
rect 22126 35112 28425 35128
rect 22126 35048 28341 35112
rect 28405 35048 28425 35112
rect 22126 35032 28425 35048
rect 22126 34968 28341 35032
rect 28405 34968 28425 35032
rect 22126 34952 28425 34968
rect 22126 34888 28341 34952
rect 28405 34888 28425 34952
rect 22126 34872 28425 34888
rect 22126 34808 28341 34872
rect 28405 34808 28425 34872
rect 22126 34792 28425 34808
rect 22126 34728 28341 34792
rect 28405 34728 28425 34792
rect 22126 34700 28425 34728
rect 28445 40872 34744 40900
rect 28445 40808 34660 40872
rect 34724 40808 34744 40872
rect 28445 40792 34744 40808
rect 28445 40728 34660 40792
rect 34724 40728 34744 40792
rect 28445 40712 34744 40728
rect 28445 40648 34660 40712
rect 34724 40648 34744 40712
rect 28445 40632 34744 40648
rect 28445 40568 34660 40632
rect 34724 40568 34744 40632
rect 28445 40552 34744 40568
rect 28445 40488 34660 40552
rect 34724 40488 34744 40552
rect 28445 40472 34744 40488
rect 28445 40408 34660 40472
rect 34724 40408 34744 40472
rect 28445 40392 34744 40408
rect 28445 40328 34660 40392
rect 34724 40328 34744 40392
rect 28445 40312 34744 40328
rect 28445 40248 34660 40312
rect 34724 40248 34744 40312
rect 28445 40232 34744 40248
rect 28445 40168 34660 40232
rect 34724 40168 34744 40232
rect 28445 40152 34744 40168
rect 28445 40088 34660 40152
rect 34724 40088 34744 40152
rect 28445 40072 34744 40088
rect 28445 40008 34660 40072
rect 34724 40008 34744 40072
rect 28445 39992 34744 40008
rect 28445 39928 34660 39992
rect 34724 39928 34744 39992
rect 28445 39912 34744 39928
rect 28445 39848 34660 39912
rect 34724 39848 34744 39912
rect 28445 39832 34744 39848
rect 28445 39768 34660 39832
rect 34724 39768 34744 39832
rect 28445 39752 34744 39768
rect 28445 39688 34660 39752
rect 34724 39688 34744 39752
rect 28445 39672 34744 39688
rect 28445 39608 34660 39672
rect 34724 39608 34744 39672
rect 28445 39592 34744 39608
rect 28445 39528 34660 39592
rect 34724 39528 34744 39592
rect 28445 39512 34744 39528
rect 28445 39448 34660 39512
rect 34724 39448 34744 39512
rect 28445 39432 34744 39448
rect 28445 39368 34660 39432
rect 34724 39368 34744 39432
rect 28445 39352 34744 39368
rect 28445 39288 34660 39352
rect 34724 39288 34744 39352
rect 28445 39272 34744 39288
rect 28445 39208 34660 39272
rect 34724 39208 34744 39272
rect 28445 39192 34744 39208
rect 28445 39128 34660 39192
rect 34724 39128 34744 39192
rect 28445 39112 34744 39128
rect 28445 39048 34660 39112
rect 34724 39048 34744 39112
rect 28445 39032 34744 39048
rect 28445 38968 34660 39032
rect 34724 38968 34744 39032
rect 28445 38952 34744 38968
rect 28445 38888 34660 38952
rect 34724 38888 34744 38952
rect 28445 38872 34744 38888
rect 28445 38808 34660 38872
rect 34724 38808 34744 38872
rect 28445 38792 34744 38808
rect 28445 38728 34660 38792
rect 34724 38728 34744 38792
rect 28445 38712 34744 38728
rect 28445 38648 34660 38712
rect 34724 38648 34744 38712
rect 28445 38632 34744 38648
rect 28445 38568 34660 38632
rect 34724 38568 34744 38632
rect 28445 38552 34744 38568
rect 28445 38488 34660 38552
rect 34724 38488 34744 38552
rect 28445 38472 34744 38488
rect 28445 38408 34660 38472
rect 34724 38408 34744 38472
rect 28445 38392 34744 38408
rect 28445 38328 34660 38392
rect 34724 38328 34744 38392
rect 28445 38312 34744 38328
rect 28445 38248 34660 38312
rect 34724 38248 34744 38312
rect 28445 38232 34744 38248
rect 28445 38168 34660 38232
rect 34724 38168 34744 38232
rect 28445 38152 34744 38168
rect 28445 38088 34660 38152
rect 34724 38088 34744 38152
rect 28445 38072 34744 38088
rect 28445 38008 34660 38072
rect 34724 38008 34744 38072
rect 28445 37992 34744 38008
rect 28445 37928 34660 37992
rect 34724 37928 34744 37992
rect 28445 37912 34744 37928
rect 28445 37848 34660 37912
rect 34724 37848 34744 37912
rect 28445 37832 34744 37848
rect 28445 37768 34660 37832
rect 34724 37768 34744 37832
rect 28445 37752 34744 37768
rect 28445 37688 34660 37752
rect 34724 37688 34744 37752
rect 28445 37672 34744 37688
rect 28445 37608 34660 37672
rect 34724 37608 34744 37672
rect 28445 37592 34744 37608
rect 28445 37528 34660 37592
rect 34724 37528 34744 37592
rect 28445 37512 34744 37528
rect 28445 37448 34660 37512
rect 34724 37448 34744 37512
rect 28445 37432 34744 37448
rect 28445 37368 34660 37432
rect 34724 37368 34744 37432
rect 28445 37352 34744 37368
rect 28445 37288 34660 37352
rect 34724 37288 34744 37352
rect 28445 37272 34744 37288
rect 28445 37208 34660 37272
rect 34724 37208 34744 37272
rect 28445 37192 34744 37208
rect 28445 37128 34660 37192
rect 34724 37128 34744 37192
rect 28445 37112 34744 37128
rect 28445 37048 34660 37112
rect 34724 37048 34744 37112
rect 28445 37032 34744 37048
rect 28445 36968 34660 37032
rect 34724 36968 34744 37032
rect 28445 36952 34744 36968
rect 28445 36888 34660 36952
rect 34724 36888 34744 36952
rect 28445 36872 34744 36888
rect 28445 36808 34660 36872
rect 34724 36808 34744 36872
rect 28445 36792 34744 36808
rect 28445 36728 34660 36792
rect 34724 36728 34744 36792
rect 28445 36712 34744 36728
rect 28445 36648 34660 36712
rect 34724 36648 34744 36712
rect 28445 36632 34744 36648
rect 28445 36568 34660 36632
rect 34724 36568 34744 36632
rect 28445 36552 34744 36568
rect 28445 36488 34660 36552
rect 34724 36488 34744 36552
rect 28445 36472 34744 36488
rect 28445 36408 34660 36472
rect 34724 36408 34744 36472
rect 28445 36392 34744 36408
rect 28445 36328 34660 36392
rect 34724 36328 34744 36392
rect 28445 36312 34744 36328
rect 28445 36248 34660 36312
rect 34724 36248 34744 36312
rect 28445 36232 34744 36248
rect 28445 36168 34660 36232
rect 34724 36168 34744 36232
rect 28445 36152 34744 36168
rect 28445 36088 34660 36152
rect 34724 36088 34744 36152
rect 28445 36072 34744 36088
rect 28445 36008 34660 36072
rect 34724 36008 34744 36072
rect 28445 35992 34744 36008
rect 28445 35928 34660 35992
rect 34724 35928 34744 35992
rect 28445 35912 34744 35928
rect 28445 35848 34660 35912
rect 34724 35848 34744 35912
rect 28445 35832 34744 35848
rect 28445 35768 34660 35832
rect 34724 35768 34744 35832
rect 28445 35752 34744 35768
rect 28445 35688 34660 35752
rect 34724 35688 34744 35752
rect 28445 35672 34744 35688
rect 28445 35608 34660 35672
rect 34724 35608 34744 35672
rect 28445 35592 34744 35608
rect 28445 35528 34660 35592
rect 34724 35528 34744 35592
rect 28445 35512 34744 35528
rect 28445 35448 34660 35512
rect 34724 35448 34744 35512
rect 28445 35432 34744 35448
rect 28445 35368 34660 35432
rect 34724 35368 34744 35432
rect 28445 35352 34744 35368
rect 28445 35288 34660 35352
rect 34724 35288 34744 35352
rect 28445 35272 34744 35288
rect 28445 35208 34660 35272
rect 34724 35208 34744 35272
rect 28445 35192 34744 35208
rect 28445 35128 34660 35192
rect 34724 35128 34744 35192
rect 28445 35112 34744 35128
rect 28445 35048 34660 35112
rect 34724 35048 34744 35112
rect 28445 35032 34744 35048
rect 28445 34968 34660 35032
rect 34724 34968 34744 35032
rect 28445 34952 34744 34968
rect 28445 34888 34660 34952
rect 34724 34888 34744 34952
rect 28445 34872 34744 34888
rect 28445 34808 34660 34872
rect 34724 34808 34744 34872
rect 28445 34792 34744 34808
rect 28445 34728 34660 34792
rect 34724 34728 34744 34792
rect 28445 34700 34744 34728
rect 34764 40872 41063 40900
rect 34764 40808 40979 40872
rect 41043 40808 41063 40872
rect 34764 40792 41063 40808
rect 34764 40728 40979 40792
rect 41043 40728 41063 40792
rect 34764 40712 41063 40728
rect 34764 40648 40979 40712
rect 41043 40648 41063 40712
rect 34764 40632 41063 40648
rect 34764 40568 40979 40632
rect 41043 40568 41063 40632
rect 34764 40552 41063 40568
rect 34764 40488 40979 40552
rect 41043 40488 41063 40552
rect 34764 40472 41063 40488
rect 34764 40408 40979 40472
rect 41043 40408 41063 40472
rect 34764 40392 41063 40408
rect 34764 40328 40979 40392
rect 41043 40328 41063 40392
rect 34764 40312 41063 40328
rect 34764 40248 40979 40312
rect 41043 40248 41063 40312
rect 34764 40232 41063 40248
rect 34764 40168 40979 40232
rect 41043 40168 41063 40232
rect 34764 40152 41063 40168
rect 34764 40088 40979 40152
rect 41043 40088 41063 40152
rect 34764 40072 41063 40088
rect 34764 40008 40979 40072
rect 41043 40008 41063 40072
rect 34764 39992 41063 40008
rect 34764 39928 40979 39992
rect 41043 39928 41063 39992
rect 34764 39912 41063 39928
rect 34764 39848 40979 39912
rect 41043 39848 41063 39912
rect 34764 39832 41063 39848
rect 34764 39768 40979 39832
rect 41043 39768 41063 39832
rect 34764 39752 41063 39768
rect 34764 39688 40979 39752
rect 41043 39688 41063 39752
rect 34764 39672 41063 39688
rect 34764 39608 40979 39672
rect 41043 39608 41063 39672
rect 34764 39592 41063 39608
rect 34764 39528 40979 39592
rect 41043 39528 41063 39592
rect 34764 39512 41063 39528
rect 34764 39448 40979 39512
rect 41043 39448 41063 39512
rect 34764 39432 41063 39448
rect 34764 39368 40979 39432
rect 41043 39368 41063 39432
rect 34764 39352 41063 39368
rect 34764 39288 40979 39352
rect 41043 39288 41063 39352
rect 34764 39272 41063 39288
rect 34764 39208 40979 39272
rect 41043 39208 41063 39272
rect 34764 39192 41063 39208
rect 34764 39128 40979 39192
rect 41043 39128 41063 39192
rect 34764 39112 41063 39128
rect 34764 39048 40979 39112
rect 41043 39048 41063 39112
rect 34764 39032 41063 39048
rect 34764 38968 40979 39032
rect 41043 38968 41063 39032
rect 34764 38952 41063 38968
rect 34764 38888 40979 38952
rect 41043 38888 41063 38952
rect 34764 38872 41063 38888
rect 34764 38808 40979 38872
rect 41043 38808 41063 38872
rect 34764 38792 41063 38808
rect 34764 38728 40979 38792
rect 41043 38728 41063 38792
rect 34764 38712 41063 38728
rect 34764 38648 40979 38712
rect 41043 38648 41063 38712
rect 34764 38632 41063 38648
rect 34764 38568 40979 38632
rect 41043 38568 41063 38632
rect 34764 38552 41063 38568
rect 34764 38488 40979 38552
rect 41043 38488 41063 38552
rect 34764 38472 41063 38488
rect 34764 38408 40979 38472
rect 41043 38408 41063 38472
rect 34764 38392 41063 38408
rect 34764 38328 40979 38392
rect 41043 38328 41063 38392
rect 34764 38312 41063 38328
rect 34764 38248 40979 38312
rect 41043 38248 41063 38312
rect 34764 38232 41063 38248
rect 34764 38168 40979 38232
rect 41043 38168 41063 38232
rect 34764 38152 41063 38168
rect 34764 38088 40979 38152
rect 41043 38088 41063 38152
rect 34764 38072 41063 38088
rect 34764 38008 40979 38072
rect 41043 38008 41063 38072
rect 34764 37992 41063 38008
rect 34764 37928 40979 37992
rect 41043 37928 41063 37992
rect 34764 37912 41063 37928
rect 34764 37848 40979 37912
rect 41043 37848 41063 37912
rect 34764 37832 41063 37848
rect 34764 37768 40979 37832
rect 41043 37768 41063 37832
rect 34764 37752 41063 37768
rect 34764 37688 40979 37752
rect 41043 37688 41063 37752
rect 34764 37672 41063 37688
rect 34764 37608 40979 37672
rect 41043 37608 41063 37672
rect 34764 37592 41063 37608
rect 34764 37528 40979 37592
rect 41043 37528 41063 37592
rect 34764 37512 41063 37528
rect 34764 37448 40979 37512
rect 41043 37448 41063 37512
rect 34764 37432 41063 37448
rect 34764 37368 40979 37432
rect 41043 37368 41063 37432
rect 34764 37352 41063 37368
rect 34764 37288 40979 37352
rect 41043 37288 41063 37352
rect 34764 37272 41063 37288
rect 34764 37208 40979 37272
rect 41043 37208 41063 37272
rect 34764 37192 41063 37208
rect 34764 37128 40979 37192
rect 41043 37128 41063 37192
rect 34764 37112 41063 37128
rect 34764 37048 40979 37112
rect 41043 37048 41063 37112
rect 34764 37032 41063 37048
rect 34764 36968 40979 37032
rect 41043 36968 41063 37032
rect 34764 36952 41063 36968
rect 34764 36888 40979 36952
rect 41043 36888 41063 36952
rect 34764 36872 41063 36888
rect 34764 36808 40979 36872
rect 41043 36808 41063 36872
rect 34764 36792 41063 36808
rect 34764 36728 40979 36792
rect 41043 36728 41063 36792
rect 34764 36712 41063 36728
rect 34764 36648 40979 36712
rect 41043 36648 41063 36712
rect 34764 36632 41063 36648
rect 34764 36568 40979 36632
rect 41043 36568 41063 36632
rect 34764 36552 41063 36568
rect 34764 36488 40979 36552
rect 41043 36488 41063 36552
rect 34764 36472 41063 36488
rect 34764 36408 40979 36472
rect 41043 36408 41063 36472
rect 34764 36392 41063 36408
rect 34764 36328 40979 36392
rect 41043 36328 41063 36392
rect 34764 36312 41063 36328
rect 34764 36248 40979 36312
rect 41043 36248 41063 36312
rect 34764 36232 41063 36248
rect 34764 36168 40979 36232
rect 41043 36168 41063 36232
rect 34764 36152 41063 36168
rect 34764 36088 40979 36152
rect 41043 36088 41063 36152
rect 34764 36072 41063 36088
rect 34764 36008 40979 36072
rect 41043 36008 41063 36072
rect 34764 35992 41063 36008
rect 34764 35928 40979 35992
rect 41043 35928 41063 35992
rect 34764 35912 41063 35928
rect 34764 35848 40979 35912
rect 41043 35848 41063 35912
rect 34764 35832 41063 35848
rect 34764 35768 40979 35832
rect 41043 35768 41063 35832
rect 34764 35752 41063 35768
rect 34764 35688 40979 35752
rect 41043 35688 41063 35752
rect 34764 35672 41063 35688
rect 34764 35608 40979 35672
rect 41043 35608 41063 35672
rect 34764 35592 41063 35608
rect 34764 35528 40979 35592
rect 41043 35528 41063 35592
rect 34764 35512 41063 35528
rect 34764 35448 40979 35512
rect 41043 35448 41063 35512
rect 34764 35432 41063 35448
rect 34764 35368 40979 35432
rect 41043 35368 41063 35432
rect 34764 35352 41063 35368
rect 34764 35288 40979 35352
rect 41043 35288 41063 35352
rect 34764 35272 41063 35288
rect 34764 35208 40979 35272
rect 41043 35208 41063 35272
rect 34764 35192 41063 35208
rect 34764 35128 40979 35192
rect 41043 35128 41063 35192
rect 34764 35112 41063 35128
rect 34764 35048 40979 35112
rect 41043 35048 41063 35112
rect 34764 35032 41063 35048
rect 34764 34968 40979 35032
rect 41043 34968 41063 35032
rect 34764 34952 41063 34968
rect 34764 34888 40979 34952
rect 41043 34888 41063 34952
rect 34764 34872 41063 34888
rect 34764 34808 40979 34872
rect 41043 34808 41063 34872
rect 34764 34792 41063 34808
rect 34764 34728 40979 34792
rect 41043 34728 41063 34792
rect 34764 34700 41063 34728
rect 41083 40872 47382 40900
rect 41083 40808 47298 40872
rect 47362 40808 47382 40872
rect 41083 40792 47382 40808
rect 41083 40728 47298 40792
rect 47362 40728 47382 40792
rect 41083 40712 47382 40728
rect 41083 40648 47298 40712
rect 47362 40648 47382 40712
rect 41083 40632 47382 40648
rect 41083 40568 47298 40632
rect 47362 40568 47382 40632
rect 41083 40552 47382 40568
rect 41083 40488 47298 40552
rect 47362 40488 47382 40552
rect 41083 40472 47382 40488
rect 41083 40408 47298 40472
rect 47362 40408 47382 40472
rect 41083 40392 47382 40408
rect 41083 40328 47298 40392
rect 47362 40328 47382 40392
rect 41083 40312 47382 40328
rect 41083 40248 47298 40312
rect 47362 40248 47382 40312
rect 41083 40232 47382 40248
rect 41083 40168 47298 40232
rect 47362 40168 47382 40232
rect 41083 40152 47382 40168
rect 41083 40088 47298 40152
rect 47362 40088 47382 40152
rect 41083 40072 47382 40088
rect 41083 40008 47298 40072
rect 47362 40008 47382 40072
rect 41083 39992 47382 40008
rect 41083 39928 47298 39992
rect 47362 39928 47382 39992
rect 41083 39912 47382 39928
rect 41083 39848 47298 39912
rect 47362 39848 47382 39912
rect 41083 39832 47382 39848
rect 41083 39768 47298 39832
rect 47362 39768 47382 39832
rect 41083 39752 47382 39768
rect 41083 39688 47298 39752
rect 47362 39688 47382 39752
rect 41083 39672 47382 39688
rect 41083 39608 47298 39672
rect 47362 39608 47382 39672
rect 41083 39592 47382 39608
rect 41083 39528 47298 39592
rect 47362 39528 47382 39592
rect 41083 39512 47382 39528
rect 41083 39448 47298 39512
rect 47362 39448 47382 39512
rect 41083 39432 47382 39448
rect 41083 39368 47298 39432
rect 47362 39368 47382 39432
rect 41083 39352 47382 39368
rect 41083 39288 47298 39352
rect 47362 39288 47382 39352
rect 41083 39272 47382 39288
rect 41083 39208 47298 39272
rect 47362 39208 47382 39272
rect 41083 39192 47382 39208
rect 41083 39128 47298 39192
rect 47362 39128 47382 39192
rect 41083 39112 47382 39128
rect 41083 39048 47298 39112
rect 47362 39048 47382 39112
rect 41083 39032 47382 39048
rect 41083 38968 47298 39032
rect 47362 38968 47382 39032
rect 41083 38952 47382 38968
rect 41083 38888 47298 38952
rect 47362 38888 47382 38952
rect 41083 38872 47382 38888
rect 41083 38808 47298 38872
rect 47362 38808 47382 38872
rect 41083 38792 47382 38808
rect 41083 38728 47298 38792
rect 47362 38728 47382 38792
rect 41083 38712 47382 38728
rect 41083 38648 47298 38712
rect 47362 38648 47382 38712
rect 41083 38632 47382 38648
rect 41083 38568 47298 38632
rect 47362 38568 47382 38632
rect 41083 38552 47382 38568
rect 41083 38488 47298 38552
rect 47362 38488 47382 38552
rect 41083 38472 47382 38488
rect 41083 38408 47298 38472
rect 47362 38408 47382 38472
rect 41083 38392 47382 38408
rect 41083 38328 47298 38392
rect 47362 38328 47382 38392
rect 41083 38312 47382 38328
rect 41083 38248 47298 38312
rect 47362 38248 47382 38312
rect 41083 38232 47382 38248
rect 41083 38168 47298 38232
rect 47362 38168 47382 38232
rect 41083 38152 47382 38168
rect 41083 38088 47298 38152
rect 47362 38088 47382 38152
rect 41083 38072 47382 38088
rect 41083 38008 47298 38072
rect 47362 38008 47382 38072
rect 41083 37992 47382 38008
rect 41083 37928 47298 37992
rect 47362 37928 47382 37992
rect 41083 37912 47382 37928
rect 41083 37848 47298 37912
rect 47362 37848 47382 37912
rect 41083 37832 47382 37848
rect 41083 37768 47298 37832
rect 47362 37768 47382 37832
rect 41083 37752 47382 37768
rect 41083 37688 47298 37752
rect 47362 37688 47382 37752
rect 41083 37672 47382 37688
rect 41083 37608 47298 37672
rect 47362 37608 47382 37672
rect 41083 37592 47382 37608
rect 41083 37528 47298 37592
rect 47362 37528 47382 37592
rect 41083 37512 47382 37528
rect 41083 37448 47298 37512
rect 47362 37448 47382 37512
rect 41083 37432 47382 37448
rect 41083 37368 47298 37432
rect 47362 37368 47382 37432
rect 41083 37352 47382 37368
rect 41083 37288 47298 37352
rect 47362 37288 47382 37352
rect 41083 37272 47382 37288
rect 41083 37208 47298 37272
rect 47362 37208 47382 37272
rect 41083 37192 47382 37208
rect 41083 37128 47298 37192
rect 47362 37128 47382 37192
rect 41083 37112 47382 37128
rect 41083 37048 47298 37112
rect 47362 37048 47382 37112
rect 41083 37032 47382 37048
rect 41083 36968 47298 37032
rect 47362 36968 47382 37032
rect 41083 36952 47382 36968
rect 41083 36888 47298 36952
rect 47362 36888 47382 36952
rect 41083 36872 47382 36888
rect 41083 36808 47298 36872
rect 47362 36808 47382 36872
rect 41083 36792 47382 36808
rect 41083 36728 47298 36792
rect 47362 36728 47382 36792
rect 41083 36712 47382 36728
rect 41083 36648 47298 36712
rect 47362 36648 47382 36712
rect 41083 36632 47382 36648
rect 41083 36568 47298 36632
rect 47362 36568 47382 36632
rect 41083 36552 47382 36568
rect 41083 36488 47298 36552
rect 47362 36488 47382 36552
rect 41083 36472 47382 36488
rect 41083 36408 47298 36472
rect 47362 36408 47382 36472
rect 41083 36392 47382 36408
rect 41083 36328 47298 36392
rect 47362 36328 47382 36392
rect 41083 36312 47382 36328
rect 41083 36248 47298 36312
rect 47362 36248 47382 36312
rect 41083 36232 47382 36248
rect 41083 36168 47298 36232
rect 47362 36168 47382 36232
rect 41083 36152 47382 36168
rect 41083 36088 47298 36152
rect 47362 36088 47382 36152
rect 41083 36072 47382 36088
rect 41083 36008 47298 36072
rect 47362 36008 47382 36072
rect 41083 35992 47382 36008
rect 41083 35928 47298 35992
rect 47362 35928 47382 35992
rect 41083 35912 47382 35928
rect 41083 35848 47298 35912
rect 47362 35848 47382 35912
rect 41083 35832 47382 35848
rect 41083 35768 47298 35832
rect 47362 35768 47382 35832
rect 41083 35752 47382 35768
rect 41083 35688 47298 35752
rect 47362 35688 47382 35752
rect 41083 35672 47382 35688
rect 41083 35608 47298 35672
rect 47362 35608 47382 35672
rect 41083 35592 47382 35608
rect 41083 35528 47298 35592
rect 47362 35528 47382 35592
rect 41083 35512 47382 35528
rect 41083 35448 47298 35512
rect 47362 35448 47382 35512
rect 41083 35432 47382 35448
rect 41083 35368 47298 35432
rect 47362 35368 47382 35432
rect 41083 35352 47382 35368
rect 41083 35288 47298 35352
rect 47362 35288 47382 35352
rect 41083 35272 47382 35288
rect 41083 35208 47298 35272
rect 47362 35208 47382 35272
rect 41083 35192 47382 35208
rect 41083 35128 47298 35192
rect 47362 35128 47382 35192
rect 41083 35112 47382 35128
rect 41083 35048 47298 35112
rect 47362 35048 47382 35112
rect 41083 35032 47382 35048
rect 41083 34968 47298 35032
rect 47362 34968 47382 35032
rect 41083 34952 47382 34968
rect 41083 34888 47298 34952
rect 47362 34888 47382 34952
rect 41083 34872 47382 34888
rect 41083 34808 47298 34872
rect 47362 34808 47382 34872
rect 41083 34792 47382 34808
rect 41083 34728 47298 34792
rect 47362 34728 47382 34792
rect 41083 34700 47382 34728
rect -47383 34572 -41084 34600
rect -47383 34508 -41168 34572
rect -41104 34508 -41084 34572
rect -47383 34492 -41084 34508
rect -47383 34428 -41168 34492
rect -41104 34428 -41084 34492
rect -47383 34412 -41084 34428
rect -47383 34348 -41168 34412
rect -41104 34348 -41084 34412
rect -47383 34332 -41084 34348
rect -47383 34268 -41168 34332
rect -41104 34268 -41084 34332
rect -47383 34252 -41084 34268
rect -47383 34188 -41168 34252
rect -41104 34188 -41084 34252
rect -47383 34172 -41084 34188
rect -47383 34108 -41168 34172
rect -41104 34108 -41084 34172
rect -47383 34092 -41084 34108
rect -47383 34028 -41168 34092
rect -41104 34028 -41084 34092
rect -47383 34012 -41084 34028
rect -47383 33948 -41168 34012
rect -41104 33948 -41084 34012
rect -47383 33932 -41084 33948
rect -47383 33868 -41168 33932
rect -41104 33868 -41084 33932
rect -47383 33852 -41084 33868
rect -47383 33788 -41168 33852
rect -41104 33788 -41084 33852
rect -47383 33772 -41084 33788
rect -47383 33708 -41168 33772
rect -41104 33708 -41084 33772
rect -47383 33692 -41084 33708
rect -47383 33628 -41168 33692
rect -41104 33628 -41084 33692
rect -47383 33612 -41084 33628
rect -47383 33548 -41168 33612
rect -41104 33548 -41084 33612
rect -47383 33532 -41084 33548
rect -47383 33468 -41168 33532
rect -41104 33468 -41084 33532
rect -47383 33452 -41084 33468
rect -47383 33388 -41168 33452
rect -41104 33388 -41084 33452
rect -47383 33372 -41084 33388
rect -47383 33308 -41168 33372
rect -41104 33308 -41084 33372
rect -47383 33292 -41084 33308
rect -47383 33228 -41168 33292
rect -41104 33228 -41084 33292
rect -47383 33212 -41084 33228
rect -47383 33148 -41168 33212
rect -41104 33148 -41084 33212
rect -47383 33132 -41084 33148
rect -47383 33068 -41168 33132
rect -41104 33068 -41084 33132
rect -47383 33052 -41084 33068
rect -47383 32988 -41168 33052
rect -41104 32988 -41084 33052
rect -47383 32972 -41084 32988
rect -47383 32908 -41168 32972
rect -41104 32908 -41084 32972
rect -47383 32892 -41084 32908
rect -47383 32828 -41168 32892
rect -41104 32828 -41084 32892
rect -47383 32812 -41084 32828
rect -47383 32748 -41168 32812
rect -41104 32748 -41084 32812
rect -47383 32732 -41084 32748
rect -47383 32668 -41168 32732
rect -41104 32668 -41084 32732
rect -47383 32652 -41084 32668
rect -47383 32588 -41168 32652
rect -41104 32588 -41084 32652
rect -47383 32572 -41084 32588
rect -47383 32508 -41168 32572
rect -41104 32508 -41084 32572
rect -47383 32492 -41084 32508
rect -47383 32428 -41168 32492
rect -41104 32428 -41084 32492
rect -47383 32412 -41084 32428
rect -47383 32348 -41168 32412
rect -41104 32348 -41084 32412
rect -47383 32332 -41084 32348
rect -47383 32268 -41168 32332
rect -41104 32268 -41084 32332
rect -47383 32252 -41084 32268
rect -47383 32188 -41168 32252
rect -41104 32188 -41084 32252
rect -47383 32172 -41084 32188
rect -47383 32108 -41168 32172
rect -41104 32108 -41084 32172
rect -47383 32092 -41084 32108
rect -47383 32028 -41168 32092
rect -41104 32028 -41084 32092
rect -47383 32012 -41084 32028
rect -47383 31948 -41168 32012
rect -41104 31948 -41084 32012
rect -47383 31932 -41084 31948
rect -47383 31868 -41168 31932
rect -41104 31868 -41084 31932
rect -47383 31852 -41084 31868
rect -47383 31788 -41168 31852
rect -41104 31788 -41084 31852
rect -47383 31772 -41084 31788
rect -47383 31708 -41168 31772
rect -41104 31708 -41084 31772
rect -47383 31692 -41084 31708
rect -47383 31628 -41168 31692
rect -41104 31628 -41084 31692
rect -47383 31612 -41084 31628
rect -47383 31548 -41168 31612
rect -41104 31548 -41084 31612
rect -47383 31532 -41084 31548
rect -47383 31468 -41168 31532
rect -41104 31468 -41084 31532
rect -47383 31452 -41084 31468
rect -47383 31388 -41168 31452
rect -41104 31388 -41084 31452
rect -47383 31372 -41084 31388
rect -47383 31308 -41168 31372
rect -41104 31308 -41084 31372
rect -47383 31292 -41084 31308
rect -47383 31228 -41168 31292
rect -41104 31228 -41084 31292
rect -47383 31212 -41084 31228
rect -47383 31148 -41168 31212
rect -41104 31148 -41084 31212
rect -47383 31132 -41084 31148
rect -47383 31068 -41168 31132
rect -41104 31068 -41084 31132
rect -47383 31052 -41084 31068
rect -47383 30988 -41168 31052
rect -41104 30988 -41084 31052
rect -47383 30972 -41084 30988
rect -47383 30908 -41168 30972
rect -41104 30908 -41084 30972
rect -47383 30892 -41084 30908
rect -47383 30828 -41168 30892
rect -41104 30828 -41084 30892
rect -47383 30812 -41084 30828
rect -47383 30748 -41168 30812
rect -41104 30748 -41084 30812
rect -47383 30732 -41084 30748
rect -47383 30668 -41168 30732
rect -41104 30668 -41084 30732
rect -47383 30652 -41084 30668
rect -47383 30588 -41168 30652
rect -41104 30588 -41084 30652
rect -47383 30572 -41084 30588
rect -47383 30508 -41168 30572
rect -41104 30508 -41084 30572
rect -47383 30492 -41084 30508
rect -47383 30428 -41168 30492
rect -41104 30428 -41084 30492
rect -47383 30412 -41084 30428
rect -47383 30348 -41168 30412
rect -41104 30348 -41084 30412
rect -47383 30332 -41084 30348
rect -47383 30268 -41168 30332
rect -41104 30268 -41084 30332
rect -47383 30252 -41084 30268
rect -47383 30188 -41168 30252
rect -41104 30188 -41084 30252
rect -47383 30172 -41084 30188
rect -47383 30108 -41168 30172
rect -41104 30108 -41084 30172
rect -47383 30092 -41084 30108
rect -47383 30028 -41168 30092
rect -41104 30028 -41084 30092
rect -47383 30012 -41084 30028
rect -47383 29948 -41168 30012
rect -41104 29948 -41084 30012
rect -47383 29932 -41084 29948
rect -47383 29868 -41168 29932
rect -41104 29868 -41084 29932
rect -47383 29852 -41084 29868
rect -47383 29788 -41168 29852
rect -41104 29788 -41084 29852
rect -47383 29772 -41084 29788
rect -47383 29708 -41168 29772
rect -41104 29708 -41084 29772
rect -47383 29692 -41084 29708
rect -47383 29628 -41168 29692
rect -41104 29628 -41084 29692
rect -47383 29612 -41084 29628
rect -47383 29548 -41168 29612
rect -41104 29548 -41084 29612
rect -47383 29532 -41084 29548
rect -47383 29468 -41168 29532
rect -41104 29468 -41084 29532
rect -47383 29452 -41084 29468
rect -47383 29388 -41168 29452
rect -41104 29388 -41084 29452
rect -47383 29372 -41084 29388
rect -47383 29308 -41168 29372
rect -41104 29308 -41084 29372
rect -47383 29292 -41084 29308
rect -47383 29228 -41168 29292
rect -41104 29228 -41084 29292
rect -47383 29212 -41084 29228
rect -47383 29148 -41168 29212
rect -41104 29148 -41084 29212
rect -47383 29132 -41084 29148
rect -47383 29068 -41168 29132
rect -41104 29068 -41084 29132
rect -47383 29052 -41084 29068
rect -47383 28988 -41168 29052
rect -41104 28988 -41084 29052
rect -47383 28972 -41084 28988
rect -47383 28908 -41168 28972
rect -41104 28908 -41084 28972
rect -47383 28892 -41084 28908
rect -47383 28828 -41168 28892
rect -41104 28828 -41084 28892
rect -47383 28812 -41084 28828
rect -47383 28748 -41168 28812
rect -41104 28748 -41084 28812
rect -47383 28732 -41084 28748
rect -47383 28668 -41168 28732
rect -41104 28668 -41084 28732
rect -47383 28652 -41084 28668
rect -47383 28588 -41168 28652
rect -41104 28588 -41084 28652
rect -47383 28572 -41084 28588
rect -47383 28508 -41168 28572
rect -41104 28508 -41084 28572
rect -47383 28492 -41084 28508
rect -47383 28428 -41168 28492
rect -41104 28428 -41084 28492
rect -47383 28400 -41084 28428
rect -41064 34572 -34765 34600
rect -41064 34508 -34849 34572
rect -34785 34508 -34765 34572
rect -41064 34492 -34765 34508
rect -41064 34428 -34849 34492
rect -34785 34428 -34765 34492
rect -41064 34412 -34765 34428
rect -41064 34348 -34849 34412
rect -34785 34348 -34765 34412
rect -41064 34332 -34765 34348
rect -41064 34268 -34849 34332
rect -34785 34268 -34765 34332
rect -41064 34252 -34765 34268
rect -41064 34188 -34849 34252
rect -34785 34188 -34765 34252
rect -41064 34172 -34765 34188
rect -41064 34108 -34849 34172
rect -34785 34108 -34765 34172
rect -41064 34092 -34765 34108
rect -41064 34028 -34849 34092
rect -34785 34028 -34765 34092
rect -41064 34012 -34765 34028
rect -41064 33948 -34849 34012
rect -34785 33948 -34765 34012
rect -41064 33932 -34765 33948
rect -41064 33868 -34849 33932
rect -34785 33868 -34765 33932
rect -41064 33852 -34765 33868
rect -41064 33788 -34849 33852
rect -34785 33788 -34765 33852
rect -41064 33772 -34765 33788
rect -41064 33708 -34849 33772
rect -34785 33708 -34765 33772
rect -41064 33692 -34765 33708
rect -41064 33628 -34849 33692
rect -34785 33628 -34765 33692
rect -41064 33612 -34765 33628
rect -41064 33548 -34849 33612
rect -34785 33548 -34765 33612
rect -41064 33532 -34765 33548
rect -41064 33468 -34849 33532
rect -34785 33468 -34765 33532
rect -41064 33452 -34765 33468
rect -41064 33388 -34849 33452
rect -34785 33388 -34765 33452
rect -41064 33372 -34765 33388
rect -41064 33308 -34849 33372
rect -34785 33308 -34765 33372
rect -41064 33292 -34765 33308
rect -41064 33228 -34849 33292
rect -34785 33228 -34765 33292
rect -41064 33212 -34765 33228
rect -41064 33148 -34849 33212
rect -34785 33148 -34765 33212
rect -41064 33132 -34765 33148
rect -41064 33068 -34849 33132
rect -34785 33068 -34765 33132
rect -41064 33052 -34765 33068
rect -41064 32988 -34849 33052
rect -34785 32988 -34765 33052
rect -41064 32972 -34765 32988
rect -41064 32908 -34849 32972
rect -34785 32908 -34765 32972
rect -41064 32892 -34765 32908
rect -41064 32828 -34849 32892
rect -34785 32828 -34765 32892
rect -41064 32812 -34765 32828
rect -41064 32748 -34849 32812
rect -34785 32748 -34765 32812
rect -41064 32732 -34765 32748
rect -41064 32668 -34849 32732
rect -34785 32668 -34765 32732
rect -41064 32652 -34765 32668
rect -41064 32588 -34849 32652
rect -34785 32588 -34765 32652
rect -41064 32572 -34765 32588
rect -41064 32508 -34849 32572
rect -34785 32508 -34765 32572
rect -41064 32492 -34765 32508
rect -41064 32428 -34849 32492
rect -34785 32428 -34765 32492
rect -41064 32412 -34765 32428
rect -41064 32348 -34849 32412
rect -34785 32348 -34765 32412
rect -41064 32332 -34765 32348
rect -41064 32268 -34849 32332
rect -34785 32268 -34765 32332
rect -41064 32252 -34765 32268
rect -41064 32188 -34849 32252
rect -34785 32188 -34765 32252
rect -41064 32172 -34765 32188
rect -41064 32108 -34849 32172
rect -34785 32108 -34765 32172
rect -41064 32092 -34765 32108
rect -41064 32028 -34849 32092
rect -34785 32028 -34765 32092
rect -41064 32012 -34765 32028
rect -41064 31948 -34849 32012
rect -34785 31948 -34765 32012
rect -41064 31932 -34765 31948
rect -41064 31868 -34849 31932
rect -34785 31868 -34765 31932
rect -41064 31852 -34765 31868
rect -41064 31788 -34849 31852
rect -34785 31788 -34765 31852
rect -41064 31772 -34765 31788
rect -41064 31708 -34849 31772
rect -34785 31708 -34765 31772
rect -41064 31692 -34765 31708
rect -41064 31628 -34849 31692
rect -34785 31628 -34765 31692
rect -41064 31612 -34765 31628
rect -41064 31548 -34849 31612
rect -34785 31548 -34765 31612
rect -41064 31532 -34765 31548
rect -41064 31468 -34849 31532
rect -34785 31468 -34765 31532
rect -41064 31452 -34765 31468
rect -41064 31388 -34849 31452
rect -34785 31388 -34765 31452
rect -41064 31372 -34765 31388
rect -41064 31308 -34849 31372
rect -34785 31308 -34765 31372
rect -41064 31292 -34765 31308
rect -41064 31228 -34849 31292
rect -34785 31228 -34765 31292
rect -41064 31212 -34765 31228
rect -41064 31148 -34849 31212
rect -34785 31148 -34765 31212
rect -41064 31132 -34765 31148
rect -41064 31068 -34849 31132
rect -34785 31068 -34765 31132
rect -41064 31052 -34765 31068
rect -41064 30988 -34849 31052
rect -34785 30988 -34765 31052
rect -41064 30972 -34765 30988
rect -41064 30908 -34849 30972
rect -34785 30908 -34765 30972
rect -41064 30892 -34765 30908
rect -41064 30828 -34849 30892
rect -34785 30828 -34765 30892
rect -41064 30812 -34765 30828
rect -41064 30748 -34849 30812
rect -34785 30748 -34765 30812
rect -41064 30732 -34765 30748
rect -41064 30668 -34849 30732
rect -34785 30668 -34765 30732
rect -41064 30652 -34765 30668
rect -41064 30588 -34849 30652
rect -34785 30588 -34765 30652
rect -41064 30572 -34765 30588
rect -41064 30508 -34849 30572
rect -34785 30508 -34765 30572
rect -41064 30492 -34765 30508
rect -41064 30428 -34849 30492
rect -34785 30428 -34765 30492
rect -41064 30412 -34765 30428
rect -41064 30348 -34849 30412
rect -34785 30348 -34765 30412
rect -41064 30332 -34765 30348
rect -41064 30268 -34849 30332
rect -34785 30268 -34765 30332
rect -41064 30252 -34765 30268
rect -41064 30188 -34849 30252
rect -34785 30188 -34765 30252
rect -41064 30172 -34765 30188
rect -41064 30108 -34849 30172
rect -34785 30108 -34765 30172
rect -41064 30092 -34765 30108
rect -41064 30028 -34849 30092
rect -34785 30028 -34765 30092
rect -41064 30012 -34765 30028
rect -41064 29948 -34849 30012
rect -34785 29948 -34765 30012
rect -41064 29932 -34765 29948
rect -41064 29868 -34849 29932
rect -34785 29868 -34765 29932
rect -41064 29852 -34765 29868
rect -41064 29788 -34849 29852
rect -34785 29788 -34765 29852
rect -41064 29772 -34765 29788
rect -41064 29708 -34849 29772
rect -34785 29708 -34765 29772
rect -41064 29692 -34765 29708
rect -41064 29628 -34849 29692
rect -34785 29628 -34765 29692
rect -41064 29612 -34765 29628
rect -41064 29548 -34849 29612
rect -34785 29548 -34765 29612
rect -41064 29532 -34765 29548
rect -41064 29468 -34849 29532
rect -34785 29468 -34765 29532
rect -41064 29452 -34765 29468
rect -41064 29388 -34849 29452
rect -34785 29388 -34765 29452
rect -41064 29372 -34765 29388
rect -41064 29308 -34849 29372
rect -34785 29308 -34765 29372
rect -41064 29292 -34765 29308
rect -41064 29228 -34849 29292
rect -34785 29228 -34765 29292
rect -41064 29212 -34765 29228
rect -41064 29148 -34849 29212
rect -34785 29148 -34765 29212
rect -41064 29132 -34765 29148
rect -41064 29068 -34849 29132
rect -34785 29068 -34765 29132
rect -41064 29052 -34765 29068
rect -41064 28988 -34849 29052
rect -34785 28988 -34765 29052
rect -41064 28972 -34765 28988
rect -41064 28908 -34849 28972
rect -34785 28908 -34765 28972
rect -41064 28892 -34765 28908
rect -41064 28828 -34849 28892
rect -34785 28828 -34765 28892
rect -41064 28812 -34765 28828
rect -41064 28748 -34849 28812
rect -34785 28748 -34765 28812
rect -41064 28732 -34765 28748
rect -41064 28668 -34849 28732
rect -34785 28668 -34765 28732
rect -41064 28652 -34765 28668
rect -41064 28588 -34849 28652
rect -34785 28588 -34765 28652
rect -41064 28572 -34765 28588
rect -41064 28508 -34849 28572
rect -34785 28508 -34765 28572
rect -41064 28492 -34765 28508
rect -41064 28428 -34849 28492
rect -34785 28428 -34765 28492
rect -41064 28400 -34765 28428
rect -34745 34572 -28446 34600
rect -34745 34508 -28530 34572
rect -28466 34508 -28446 34572
rect -34745 34492 -28446 34508
rect -34745 34428 -28530 34492
rect -28466 34428 -28446 34492
rect -34745 34412 -28446 34428
rect -34745 34348 -28530 34412
rect -28466 34348 -28446 34412
rect -34745 34332 -28446 34348
rect -34745 34268 -28530 34332
rect -28466 34268 -28446 34332
rect -34745 34252 -28446 34268
rect -34745 34188 -28530 34252
rect -28466 34188 -28446 34252
rect -34745 34172 -28446 34188
rect -34745 34108 -28530 34172
rect -28466 34108 -28446 34172
rect -34745 34092 -28446 34108
rect -34745 34028 -28530 34092
rect -28466 34028 -28446 34092
rect -34745 34012 -28446 34028
rect -34745 33948 -28530 34012
rect -28466 33948 -28446 34012
rect -34745 33932 -28446 33948
rect -34745 33868 -28530 33932
rect -28466 33868 -28446 33932
rect -34745 33852 -28446 33868
rect -34745 33788 -28530 33852
rect -28466 33788 -28446 33852
rect -34745 33772 -28446 33788
rect -34745 33708 -28530 33772
rect -28466 33708 -28446 33772
rect -34745 33692 -28446 33708
rect -34745 33628 -28530 33692
rect -28466 33628 -28446 33692
rect -34745 33612 -28446 33628
rect -34745 33548 -28530 33612
rect -28466 33548 -28446 33612
rect -34745 33532 -28446 33548
rect -34745 33468 -28530 33532
rect -28466 33468 -28446 33532
rect -34745 33452 -28446 33468
rect -34745 33388 -28530 33452
rect -28466 33388 -28446 33452
rect -34745 33372 -28446 33388
rect -34745 33308 -28530 33372
rect -28466 33308 -28446 33372
rect -34745 33292 -28446 33308
rect -34745 33228 -28530 33292
rect -28466 33228 -28446 33292
rect -34745 33212 -28446 33228
rect -34745 33148 -28530 33212
rect -28466 33148 -28446 33212
rect -34745 33132 -28446 33148
rect -34745 33068 -28530 33132
rect -28466 33068 -28446 33132
rect -34745 33052 -28446 33068
rect -34745 32988 -28530 33052
rect -28466 32988 -28446 33052
rect -34745 32972 -28446 32988
rect -34745 32908 -28530 32972
rect -28466 32908 -28446 32972
rect -34745 32892 -28446 32908
rect -34745 32828 -28530 32892
rect -28466 32828 -28446 32892
rect -34745 32812 -28446 32828
rect -34745 32748 -28530 32812
rect -28466 32748 -28446 32812
rect -34745 32732 -28446 32748
rect -34745 32668 -28530 32732
rect -28466 32668 -28446 32732
rect -34745 32652 -28446 32668
rect -34745 32588 -28530 32652
rect -28466 32588 -28446 32652
rect -34745 32572 -28446 32588
rect -34745 32508 -28530 32572
rect -28466 32508 -28446 32572
rect -34745 32492 -28446 32508
rect -34745 32428 -28530 32492
rect -28466 32428 -28446 32492
rect -34745 32412 -28446 32428
rect -34745 32348 -28530 32412
rect -28466 32348 -28446 32412
rect -34745 32332 -28446 32348
rect -34745 32268 -28530 32332
rect -28466 32268 -28446 32332
rect -34745 32252 -28446 32268
rect -34745 32188 -28530 32252
rect -28466 32188 -28446 32252
rect -34745 32172 -28446 32188
rect -34745 32108 -28530 32172
rect -28466 32108 -28446 32172
rect -34745 32092 -28446 32108
rect -34745 32028 -28530 32092
rect -28466 32028 -28446 32092
rect -34745 32012 -28446 32028
rect -34745 31948 -28530 32012
rect -28466 31948 -28446 32012
rect -34745 31932 -28446 31948
rect -34745 31868 -28530 31932
rect -28466 31868 -28446 31932
rect -34745 31852 -28446 31868
rect -34745 31788 -28530 31852
rect -28466 31788 -28446 31852
rect -34745 31772 -28446 31788
rect -34745 31708 -28530 31772
rect -28466 31708 -28446 31772
rect -34745 31692 -28446 31708
rect -34745 31628 -28530 31692
rect -28466 31628 -28446 31692
rect -34745 31612 -28446 31628
rect -34745 31548 -28530 31612
rect -28466 31548 -28446 31612
rect -34745 31532 -28446 31548
rect -34745 31468 -28530 31532
rect -28466 31468 -28446 31532
rect -34745 31452 -28446 31468
rect -34745 31388 -28530 31452
rect -28466 31388 -28446 31452
rect -34745 31372 -28446 31388
rect -34745 31308 -28530 31372
rect -28466 31308 -28446 31372
rect -34745 31292 -28446 31308
rect -34745 31228 -28530 31292
rect -28466 31228 -28446 31292
rect -34745 31212 -28446 31228
rect -34745 31148 -28530 31212
rect -28466 31148 -28446 31212
rect -34745 31132 -28446 31148
rect -34745 31068 -28530 31132
rect -28466 31068 -28446 31132
rect -34745 31052 -28446 31068
rect -34745 30988 -28530 31052
rect -28466 30988 -28446 31052
rect -34745 30972 -28446 30988
rect -34745 30908 -28530 30972
rect -28466 30908 -28446 30972
rect -34745 30892 -28446 30908
rect -34745 30828 -28530 30892
rect -28466 30828 -28446 30892
rect -34745 30812 -28446 30828
rect -34745 30748 -28530 30812
rect -28466 30748 -28446 30812
rect -34745 30732 -28446 30748
rect -34745 30668 -28530 30732
rect -28466 30668 -28446 30732
rect -34745 30652 -28446 30668
rect -34745 30588 -28530 30652
rect -28466 30588 -28446 30652
rect -34745 30572 -28446 30588
rect -34745 30508 -28530 30572
rect -28466 30508 -28446 30572
rect -34745 30492 -28446 30508
rect -34745 30428 -28530 30492
rect -28466 30428 -28446 30492
rect -34745 30412 -28446 30428
rect -34745 30348 -28530 30412
rect -28466 30348 -28446 30412
rect -34745 30332 -28446 30348
rect -34745 30268 -28530 30332
rect -28466 30268 -28446 30332
rect -34745 30252 -28446 30268
rect -34745 30188 -28530 30252
rect -28466 30188 -28446 30252
rect -34745 30172 -28446 30188
rect -34745 30108 -28530 30172
rect -28466 30108 -28446 30172
rect -34745 30092 -28446 30108
rect -34745 30028 -28530 30092
rect -28466 30028 -28446 30092
rect -34745 30012 -28446 30028
rect -34745 29948 -28530 30012
rect -28466 29948 -28446 30012
rect -34745 29932 -28446 29948
rect -34745 29868 -28530 29932
rect -28466 29868 -28446 29932
rect -34745 29852 -28446 29868
rect -34745 29788 -28530 29852
rect -28466 29788 -28446 29852
rect -34745 29772 -28446 29788
rect -34745 29708 -28530 29772
rect -28466 29708 -28446 29772
rect -34745 29692 -28446 29708
rect -34745 29628 -28530 29692
rect -28466 29628 -28446 29692
rect -34745 29612 -28446 29628
rect -34745 29548 -28530 29612
rect -28466 29548 -28446 29612
rect -34745 29532 -28446 29548
rect -34745 29468 -28530 29532
rect -28466 29468 -28446 29532
rect -34745 29452 -28446 29468
rect -34745 29388 -28530 29452
rect -28466 29388 -28446 29452
rect -34745 29372 -28446 29388
rect -34745 29308 -28530 29372
rect -28466 29308 -28446 29372
rect -34745 29292 -28446 29308
rect -34745 29228 -28530 29292
rect -28466 29228 -28446 29292
rect -34745 29212 -28446 29228
rect -34745 29148 -28530 29212
rect -28466 29148 -28446 29212
rect -34745 29132 -28446 29148
rect -34745 29068 -28530 29132
rect -28466 29068 -28446 29132
rect -34745 29052 -28446 29068
rect -34745 28988 -28530 29052
rect -28466 28988 -28446 29052
rect -34745 28972 -28446 28988
rect -34745 28908 -28530 28972
rect -28466 28908 -28446 28972
rect -34745 28892 -28446 28908
rect -34745 28828 -28530 28892
rect -28466 28828 -28446 28892
rect -34745 28812 -28446 28828
rect -34745 28748 -28530 28812
rect -28466 28748 -28446 28812
rect -34745 28732 -28446 28748
rect -34745 28668 -28530 28732
rect -28466 28668 -28446 28732
rect -34745 28652 -28446 28668
rect -34745 28588 -28530 28652
rect -28466 28588 -28446 28652
rect -34745 28572 -28446 28588
rect -34745 28508 -28530 28572
rect -28466 28508 -28446 28572
rect -34745 28492 -28446 28508
rect -34745 28428 -28530 28492
rect -28466 28428 -28446 28492
rect -34745 28400 -28446 28428
rect -28426 34572 -22127 34600
rect -28426 34508 -22211 34572
rect -22147 34508 -22127 34572
rect -28426 34492 -22127 34508
rect -28426 34428 -22211 34492
rect -22147 34428 -22127 34492
rect -28426 34412 -22127 34428
rect -28426 34348 -22211 34412
rect -22147 34348 -22127 34412
rect -28426 34332 -22127 34348
rect -28426 34268 -22211 34332
rect -22147 34268 -22127 34332
rect -28426 34252 -22127 34268
rect -28426 34188 -22211 34252
rect -22147 34188 -22127 34252
rect -28426 34172 -22127 34188
rect -28426 34108 -22211 34172
rect -22147 34108 -22127 34172
rect -28426 34092 -22127 34108
rect -28426 34028 -22211 34092
rect -22147 34028 -22127 34092
rect -28426 34012 -22127 34028
rect -28426 33948 -22211 34012
rect -22147 33948 -22127 34012
rect -28426 33932 -22127 33948
rect -28426 33868 -22211 33932
rect -22147 33868 -22127 33932
rect -28426 33852 -22127 33868
rect -28426 33788 -22211 33852
rect -22147 33788 -22127 33852
rect -28426 33772 -22127 33788
rect -28426 33708 -22211 33772
rect -22147 33708 -22127 33772
rect -28426 33692 -22127 33708
rect -28426 33628 -22211 33692
rect -22147 33628 -22127 33692
rect -28426 33612 -22127 33628
rect -28426 33548 -22211 33612
rect -22147 33548 -22127 33612
rect -28426 33532 -22127 33548
rect -28426 33468 -22211 33532
rect -22147 33468 -22127 33532
rect -28426 33452 -22127 33468
rect -28426 33388 -22211 33452
rect -22147 33388 -22127 33452
rect -28426 33372 -22127 33388
rect -28426 33308 -22211 33372
rect -22147 33308 -22127 33372
rect -28426 33292 -22127 33308
rect -28426 33228 -22211 33292
rect -22147 33228 -22127 33292
rect -28426 33212 -22127 33228
rect -28426 33148 -22211 33212
rect -22147 33148 -22127 33212
rect -28426 33132 -22127 33148
rect -28426 33068 -22211 33132
rect -22147 33068 -22127 33132
rect -28426 33052 -22127 33068
rect -28426 32988 -22211 33052
rect -22147 32988 -22127 33052
rect -28426 32972 -22127 32988
rect -28426 32908 -22211 32972
rect -22147 32908 -22127 32972
rect -28426 32892 -22127 32908
rect -28426 32828 -22211 32892
rect -22147 32828 -22127 32892
rect -28426 32812 -22127 32828
rect -28426 32748 -22211 32812
rect -22147 32748 -22127 32812
rect -28426 32732 -22127 32748
rect -28426 32668 -22211 32732
rect -22147 32668 -22127 32732
rect -28426 32652 -22127 32668
rect -28426 32588 -22211 32652
rect -22147 32588 -22127 32652
rect -28426 32572 -22127 32588
rect -28426 32508 -22211 32572
rect -22147 32508 -22127 32572
rect -28426 32492 -22127 32508
rect -28426 32428 -22211 32492
rect -22147 32428 -22127 32492
rect -28426 32412 -22127 32428
rect -28426 32348 -22211 32412
rect -22147 32348 -22127 32412
rect -28426 32332 -22127 32348
rect -28426 32268 -22211 32332
rect -22147 32268 -22127 32332
rect -28426 32252 -22127 32268
rect -28426 32188 -22211 32252
rect -22147 32188 -22127 32252
rect -28426 32172 -22127 32188
rect -28426 32108 -22211 32172
rect -22147 32108 -22127 32172
rect -28426 32092 -22127 32108
rect -28426 32028 -22211 32092
rect -22147 32028 -22127 32092
rect -28426 32012 -22127 32028
rect -28426 31948 -22211 32012
rect -22147 31948 -22127 32012
rect -28426 31932 -22127 31948
rect -28426 31868 -22211 31932
rect -22147 31868 -22127 31932
rect -28426 31852 -22127 31868
rect -28426 31788 -22211 31852
rect -22147 31788 -22127 31852
rect -28426 31772 -22127 31788
rect -28426 31708 -22211 31772
rect -22147 31708 -22127 31772
rect -28426 31692 -22127 31708
rect -28426 31628 -22211 31692
rect -22147 31628 -22127 31692
rect -28426 31612 -22127 31628
rect -28426 31548 -22211 31612
rect -22147 31548 -22127 31612
rect -28426 31532 -22127 31548
rect -28426 31468 -22211 31532
rect -22147 31468 -22127 31532
rect -28426 31452 -22127 31468
rect -28426 31388 -22211 31452
rect -22147 31388 -22127 31452
rect -28426 31372 -22127 31388
rect -28426 31308 -22211 31372
rect -22147 31308 -22127 31372
rect -28426 31292 -22127 31308
rect -28426 31228 -22211 31292
rect -22147 31228 -22127 31292
rect -28426 31212 -22127 31228
rect -28426 31148 -22211 31212
rect -22147 31148 -22127 31212
rect -28426 31132 -22127 31148
rect -28426 31068 -22211 31132
rect -22147 31068 -22127 31132
rect -28426 31052 -22127 31068
rect -28426 30988 -22211 31052
rect -22147 30988 -22127 31052
rect -28426 30972 -22127 30988
rect -28426 30908 -22211 30972
rect -22147 30908 -22127 30972
rect -28426 30892 -22127 30908
rect -28426 30828 -22211 30892
rect -22147 30828 -22127 30892
rect -28426 30812 -22127 30828
rect -28426 30748 -22211 30812
rect -22147 30748 -22127 30812
rect -28426 30732 -22127 30748
rect -28426 30668 -22211 30732
rect -22147 30668 -22127 30732
rect -28426 30652 -22127 30668
rect -28426 30588 -22211 30652
rect -22147 30588 -22127 30652
rect -28426 30572 -22127 30588
rect -28426 30508 -22211 30572
rect -22147 30508 -22127 30572
rect -28426 30492 -22127 30508
rect -28426 30428 -22211 30492
rect -22147 30428 -22127 30492
rect -28426 30412 -22127 30428
rect -28426 30348 -22211 30412
rect -22147 30348 -22127 30412
rect -28426 30332 -22127 30348
rect -28426 30268 -22211 30332
rect -22147 30268 -22127 30332
rect -28426 30252 -22127 30268
rect -28426 30188 -22211 30252
rect -22147 30188 -22127 30252
rect -28426 30172 -22127 30188
rect -28426 30108 -22211 30172
rect -22147 30108 -22127 30172
rect -28426 30092 -22127 30108
rect -28426 30028 -22211 30092
rect -22147 30028 -22127 30092
rect -28426 30012 -22127 30028
rect -28426 29948 -22211 30012
rect -22147 29948 -22127 30012
rect -28426 29932 -22127 29948
rect -28426 29868 -22211 29932
rect -22147 29868 -22127 29932
rect -28426 29852 -22127 29868
rect -28426 29788 -22211 29852
rect -22147 29788 -22127 29852
rect -28426 29772 -22127 29788
rect -28426 29708 -22211 29772
rect -22147 29708 -22127 29772
rect -28426 29692 -22127 29708
rect -28426 29628 -22211 29692
rect -22147 29628 -22127 29692
rect -28426 29612 -22127 29628
rect -28426 29548 -22211 29612
rect -22147 29548 -22127 29612
rect -28426 29532 -22127 29548
rect -28426 29468 -22211 29532
rect -22147 29468 -22127 29532
rect -28426 29452 -22127 29468
rect -28426 29388 -22211 29452
rect -22147 29388 -22127 29452
rect -28426 29372 -22127 29388
rect -28426 29308 -22211 29372
rect -22147 29308 -22127 29372
rect -28426 29292 -22127 29308
rect -28426 29228 -22211 29292
rect -22147 29228 -22127 29292
rect -28426 29212 -22127 29228
rect -28426 29148 -22211 29212
rect -22147 29148 -22127 29212
rect -28426 29132 -22127 29148
rect -28426 29068 -22211 29132
rect -22147 29068 -22127 29132
rect -28426 29052 -22127 29068
rect -28426 28988 -22211 29052
rect -22147 28988 -22127 29052
rect -28426 28972 -22127 28988
rect -28426 28908 -22211 28972
rect -22147 28908 -22127 28972
rect -28426 28892 -22127 28908
rect -28426 28828 -22211 28892
rect -22147 28828 -22127 28892
rect -28426 28812 -22127 28828
rect -28426 28748 -22211 28812
rect -22147 28748 -22127 28812
rect -28426 28732 -22127 28748
rect -28426 28668 -22211 28732
rect -22147 28668 -22127 28732
rect -28426 28652 -22127 28668
rect -28426 28588 -22211 28652
rect -22147 28588 -22127 28652
rect -28426 28572 -22127 28588
rect -28426 28508 -22211 28572
rect -22147 28508 -22127 28572
rect -28426 28492 -22127 28508
rect -28426 28428 -22211 28492
rect -22147 28428 -22127 28492
rect -28426 28400 -22127 28428
rect -22107 34572 -15808 34600
rect -22107 34508 -15892 34572
rect -15828 34508 -15808 34572
rect -22107 34492 -15808 34508
rect -22107 34428 -15892 34492
rect -15828 34428 -15808 34492
rect -22107 34412 -15808 34428
rect -22107 34348 -15892 34412
rect -15828 34348 -15808 34412
rect -22107 34332 -15808 34348
rect -22107 34268 -15892 34332
rect -15828 34268 -15808 34332
rect -22107 34252 -15808 34268
rect -22107 34188 -15892 34252
rect -15828 34188 -15808 34252
rect -22107 34172 -15808 34188
rect -22107 34108 -15892 34172
rect -15828 34108 -15808 34172
rect -22107 34092 -15808 34108
rect -22107 34028 -15892 34092
rect -15828 34028 -15808 34092
rect -22107 34012 -15808 34028
rect -22107 33948 -15892 34012
rect -15828 33948 -15808 34012
rect -22107 33932 -15808 33948
rect -22107 33868 -15892 33932
rect -15828 33868 -15808 33932
rect -22107 33852 -15808 33868
rect -22107 33788 -15892 33852
rect -15828 33788 -15808 33852
rect -22107 33772 -15808 33788
rect -22107 33708 -15892 33772
rect -15828 33708 -15808 33772
rect -22107 33692 -15808 33708
rect -22107 33628 -15892 33692
rect -15828 33628 -15808 33692
rect -22107 33612 -15808 33628
rect -22107 33548 -15892 33612
rect -15828 33548 -15808 33612
rect -22107 33532 -15808 33548
rect -22107 33468 -15892 33532
rect -15828 33468 -15808 33532
rect -22107 33452 -15808 33468
rect -22107 33388 -15892 33452
rect -15828 33388 -15808 33452
rect -22107 33372 -15808 33388
rect -22107 33308 -15892 33372
rect -15828 33308 -15808 33372
rect -22107 33292 -15808 33308
rect -22107 33228 -15892 33292
rect -15828 33228 -15808 33292
rect -22107 33212 -15808 33228
rect -22107 33148 -15892 33212
rect -15828 33148 -15808 33212
rect -22107 33132 -15808 33148
rect -22107 33068 -15892 33132
rect -15828 33068 -15808 33132
rect -22107 33052 -15808 33068
rect -22107 32988 -15892 33052
rect -15828 32988 -15808 33052
rect -22107 32972 -15808 32988
rect -22107 32908 -15892 32972
rect -15828 32908 -15808 32972
rect -22107 32892 -15808 32908
rect -22107 32828 -15892 32892
rect -15828 32828 -15808 32892
rect -22107 32812 -15808 32828
rect -22107 32748 -15892 32812
rect -15828 32748 -15808 32812
rect -22107 32732 -15808 32748
rect -22107 32668 -15892 32732
rect -15828 32668 -15808 32732
rect -22107 32652 -15808 32668
rect -22107 32588 -15892 32652
rect -15828 32588 -15808 32652
rect -22107 32572 -15808 32588
rect -22107 32508 -15892 32572
rect -15828 32508 -15808 32572
rect -22107 32492 -15808 32508
rect -22107 32428 -15892 32492
rect -15828 32428 -15808 32492
rect -22107 32412 -15808 32428
rect -22107 32348 -15892 32412
rect -15828 32348 -15808 32412
rect -22107 32332 -15808 32348
rect -22107 32268 -15892 32332
rect -15828 32268 -15808 32332
rect -22107 32252 -15808 32268
rect -22107 32188 -15892 32252
rect -15828 32188 -15808 32252
rect -22107 32172 -15808 32188
rect -22107 32108 -15892 32172
rect -15828 32108 -15808 32172
rect -22107 32092 -15808 32108
rect -22107 32028 -15892 32092
rect -15828 32028 -15808 32092
rect -22107 32012 -15808 32028
rect -22107 31948 -15892 32012
rect -15828 31948 -15808 32012
rect -22107 31932 -15808 31948
rect -22107 31868 -15892 31932
rect -15828 31868 -15808 31932
rect -22107 31852 -15808 31868
rect -22107 31788 -15892 31852
rect -15828 31788 -15808 31852
rect -22107 31772 -15808 31788
rect -22107 31708 -15892 31772
rect -15828 31708 -15808 31772
rect -22107 31692 -15808 31708
rect -22107 31628 -15892 31692
rect -15828 31628 -15808 31692
rect -22107 31612 -15808 31628
rect -22107 31548 -15892 31612
rect -15828 31548 -15808 31612
rect -22107 31532 -15808 31548
rect -22107 31468 -15892 31532
rect -15828 31468 -15808 31532
rect -22107 31452 -15808 31468
rect -22107 31388 -15892 31452
rect -15828 31388 -15808 31452
rect -22107 31372 -15808 31388
rect -22107 31308 -15892 31372
rect -15828 31308 -15808 31372
rect -22107 31292 -15808 31308
rect -22107 31228 -15892 31292
rect -15828 31228 -15808 31292
rect -22107 31212 -15808 31228
rect -22107 31148 -15892 31212
rect -15828 31148 -15808 31212
rect -22107 31132 -15808 31148
rect -22107 31068 -15892 31132
rect -15828 31068 -15808 31132
rect -22107 31052 -15808 31068
rect -22107 30988 -15892 31052
rect -15828 30988 -15808 31052
rect -22107 30972 -15808 30988
rect -22107 30908 -15892 30972
rect -15828 30908 -15808 30972
rect -22107 30892 -15808 30908
rect -22107 30828 -15892 30892
rect -15828 30828 -15808 30892
rect -22107 30812 -15808 30828
rect -22107 30748 -15892 30812
rect -15828 30748 -15808 30812
rect -22107 30732 -15808 30748
rect -22107 30668 -15892 30732
rect -15828 30668 -15808 30732
rect -22107 30652 -15808 30668
rect -22107 30588 -15892 30652
rect -15828 30588 -15808 30652
rect -22107 30572 -15808 30588
rect -22107 30508 -15892 30572
rect -15828 30508 -15808 30572
rect -22107 30492 -15808 30508
rect -22107 30428 -15892 30492
rect -15828 30428 -15808 30492
rect -22107 30412 -15808 30428
rect -22107 30348 -15892 30412
rect -15828 30348 -15808 30412
rect -22107 30332 -15808 30348
rect -22107 30268 -15892 30332
rect -15828 30268 -15808 30332
rect -22107 30252 -15808 30268
rect -22107 30188 -15892 30252
rect -15828 30188 -15808 30252
rect -22107 30172 -15808 30188
rect -22107 30108 -15892 30172
rect -15828 30108 -15808 30172
rect -22107 30092 -15808 30108
rect -22107 30028 -15892 30092
rect -15828 30028 -15808 30092
rect -22107 30012 -15808 30028
rect -22107 29948 -15892 30012
rect -15828 29948 -15808 30012
rect -22107 29932 -15808 29948
rect -22107 29868 -15892 29932
rect -15828 29868 -15808 29932
rect -22107 29852 -15808 29868
rect -22107 29788 -15892 29852
rect -15828 29788 -15808 29852
rect -22107 29772 -15808 29788
rect -22107 29708 -15892 29772
rect -15828 29708 -15808 29772
rect -22107 29692 -15808 29708
rect -22107 29628 -15892 29692
rect -15828 29628 -15808 29692
rect -22107 29612 -15808 29628
rect -22107 29548 -15892 29612
rect -15828 29548 -15808 29612
rect -22107 29532 -15808 29548
rect -22107 29468 -15892 29532
rect -15828 29468 -15808 29532
rect -22107 29452 -15808 29468
rect -22107 29388 -15892 29452
rect -15828 29388 -15808 29452
rect -22107 29372 -15808 29388
rect -22107 29308 -15892 29372
rect -15828 29308 -15808 29372
rect -22107 29292 -15808 29308
rect -22107 29228 -15892 29292
rect -15828 29228 -15808 29292
rect -22107 29212 -15808 29228
rect -22107 29148 -15892 29212
rect -15828 29148 -15808 29212
rect -22107 29132 -15808 29148
rect -22107 29068 -15892 29132
rect -15828 29068 -15808 29132
rect -22107 29052 -15808 29068
rect -22107 28988 -15892 29052
rect -15828 28988 -15808 29052
rect -22107 28972 -15808 28988
rect -22107 28908 -15892 28972
rect -15828 28908 -15808 28972
rect -22107 28892 -15808 28908
rect -22107 28828 -15892 28892
rect -15828 28828 -15808 28892
rect -22107 28812 -15808 28828
rect -22107 28748 -15892 28812
rect -15828 28748 -15808 28812
rect -22107 28732 -15808 28748
rect -22107 28668 -15892 28732
rect -15828 28668 -15808 28732
rect -22107 28652 -15808 28668
rect -22107 28588 -15892 28652
rect -15828 28588 -15808 28652
rect -22107 28572 -15808 28588
rect -22107 28508 -15892 28572
rect -15828 28508 -15808 28572
rect -22107 28492 -15808 28508
rect -22107 28428 -15892 28492
rect -15828 28428 -15808 28492
rect -22107 28400 -15808 28428
rect -15788 34572 -9489 34600
rect -15788 34508 -9573 34572
rect -9509 34508 -9489 34572
rect -15788 34492 -9489 34508
rect -15788 34428 -9573 34492
rect -9509 34428 -9489 34492
rect -15788 34412 -9489 34428
rect -15788 34348 -9573 34412
rect -9509 34348 -9489 34412
rect -15788 34332 -9489 34348
rect -15788 34268 -9573 34332
rect -9509 34268 -9489 34332
rect -15788 34252 -9489 34268
rect -15788 34188 -9573 34252
rect -9509 34188 -9489 34252
rect -15788 34172 -9489 34188
rect -15788 34108 -9573 34172
rect -9509 34108 -9489 34172
rect -15788 34092 -9489 34108
rect -15788 34028 -9573 34092
rect -9509 34028 -9489 34092
rect -15788 34012 -9489 34028
rect -15788 33948 -9573 34012
rect -9509 33948 -9489 34012
rect -15788 33932 -9489 33948
rect -15788 33868 -9573 33932
rect -9509 33868 -9489 33932
rect -15788 33852 -9489 33868
rect -15788 33788 -9573 33852
rect -9509 33788 -9489 33852
rect -15788 33772 -9489 33788
rect -15788 33708 -9573 33772
rect -9509 33708 -9489 33772
rect -15788 33692 -9489 33708
rect -15788 33628 -9573 33692
rect -9509 33628 -9489 33692
rect -15788 33612 -9489 33628
rect -15788 33548 -9573 33612
rect -9509 33548 -9489 33612
rect -15788 33532 -9489 33548
rect -15788 33468 -9573 33532
rect -9509 33468 -9489 33532
rect -15788 33452 -9489 33468
rect -15788 33388 -9573 33452
rect -9509 33388 -9489 33452
rect -15788 33372 -9489 33388
rect -15788 33308 -9573 33372
rect -9509 33308 -9489 33372
rect -15788 33292 -9489 33308
rect -15788 33228 -9573 33292
rect -9509 33228 -9489 33292
rect -15788 33212 -9489 33228
rect -15788 33148 -9573 33212
rect -9509 33148 -9489 33212
rect -15788 33132 -9489 33148
rect -15788 33068 -9573 33132
rect -9509 33068 -9489 33132
rect -15788 33052 -9489 33068
rect -15788 32988 -9573 33052
rect -9509 32988 -9489 33052
rect -15788 32972 -9489 32988
rect -15788 32908 -9573 32972
rect -9509 32908 -9489 32972
rect -15788 32892 -9489 32908
rect -15788 32828 -9573 32892
rect -9509 32828 -9489 32892
rect -15788 32812 -9489 32828
rect -15788 32748 -9573 32812
rect -9509 32748 -9489 32812
rect -15788 32732 -9489 32748
rect -15788 32668 -9573 32732
rect -9509 32668 -9489 32732
rect -15788 32652 -9489 32668
rect -15788 32588 -9573 32652
rect -9509 32588 -9489 32652
rect -15788 32572 -9489 32588
rect -15788 32508 -9573 32572
rect -9509 32508 -9489 32572
rect -15788 32492 -9489 32508
rect -15788 32428 -9573 32492
rect -9509 32428 -9489 32492
rect -15788 32412 -9489 32428
rect -15788 32348 -9573 32412
rect -9509 32348 -9489 32412
rect -15788 32332 -9489 32348
rect -15788 32268 -9573 32332
rect -9509 32268 -9489 32332
rect -15788 32252 -9489 32268
rect -15788 32188 -9573 32252
rect -9509 32188 -9489 32252
rect -15788 32172 -9489 32188
rect -15788 32108 -9573 32172
rect -9509 32108 -9489 32172
rect -15788 32092 -9489 32108
rect -15788 32028 -9573 32092
rect -9509 32028 -9489 32092
rect -15788 32012 -9489 32028
rect -15788 31948 -9573 32012
rect -9509 31948 -9489 32012
rect -15788 31932 -9489 31948
rect -15788 31868 -9573 31932
rect -9509 31868 -9489 31932
rect -15788 31852 -9489 31868
rect -15788 31788 -9573 31852
rect -9509 31788 -9489 31852
rect -15788 31772 -9489 31788
rect -15788 31708 -9573 31772
rect -9509 31708 -9489 31772
rect -15788 31692 -9489 31708
rect -15788 31628 -9573 31692
rect -9509 31628 -9489 31692
rect -15788 31612 -9489 31628
rect -15788 31548 -9573 31612
rect -9509 31548 -9489 31612
rect -15788 31532 -9489 31548
rect -15788 31468 -9573 31532
rect -9509 31468 -9489 31532
rect -15788 31452 -9489 31468
rect -15788 31388 -9573 31452
rect -9509 31388 -9489 31452
rect -15788 31372 -9489 31388
rect -15788 31308 -9573 31372
rect -9509 31308 -9489 31372
rect -15788 31292 -9489 31308
rect -15788 31228 -9573 31292
rect -9509 31228 -9489 31292
rect -15788 31212 -9489 31228
rect -15788 31148 -9573 31212
rect -9509 31148 -9489 31212
rect -15788 31132 -9489 31148
rect -15788 31068 -9573 31132
rect -9509 31068 -9489 31132
rect -15788 31052 -9489 31068
rect -15788 30988 -9573 31052
rect -9509 30988 -9489 31052
rect -15788 30972 -9489 30988
rect -15788 30908 -9573 30972
rect -9509 30908 -9489 30972
rect -15788 30892 -9489 30908
rect -15788 30828 -9573 30892
rect -9509 30828 -9489 30892
rect -15788 30812 -9489 30828
rect -15788 30748 -9573 30812
rect -9509 30748 -9489 30812
rect -15788 30732 -9489 30748
rect -15788 30668 -9573 30732
rect -9509 30668 -9489 30732
rect -15788 30652 -9489 30668
rect -15788 30588 -9573 30652
rect -9509 30588 -9489 30652
rect -15788 30572 -9489 30588
rect -15788 30508 -9573 30572
rect -9509 30508 -9489 30572
rect -15788 30492 -9489 30508
rect -15788 30428 -9573 30492
rect -9509 30428 -9489 30492
rect -15788 30412 -9489 30428
rect -15788 30348 -9573 30412
rect -9509 30348 -9489 30412
rect -15788 30332 -9489 30348
rect -15788 30268 -9573 30332
rect -9509 30268 -9489 30332
rect -15788 30252 -9489 30268
rect -15788 30188 -9573 30252
rect -9509 30188 -9489 30252
rect -15788 30172 -9489 30188
rect -15788 30108 -9573 30172
rect -9509 30108 -9489 30172
rect -15788 30092 -9489 30108
rect -15788 30028 -9573 30092
rect -9509 30028 -9489 30092
rect -15788 30012 -9489 30028
rect -15788 29948 -9573 30012
rect -9509 29948 -9489 30012
rect -15788 29932 -9489 29948
rect -15788 29868 -9573 29932
rect -9509 29868 -9489 29932
rect -15788 29852 -9489 29868
rect -15788 29788 -9573 29852
rect -9509 29788 -9489 29852
rect -15788 29772 -9489 29788
rect -15788 29708 -9573 29772
rect -9509 29708 -9489 29772
rect -15788 29692 -9489 29708
rect -15788 29628 -9573 29692
rect -9509 29628 -9489 29692
rect -15788 29612 -9489 29628
rect -15788 29548 -9573 29612
rect -9509 29548 -9489 29612
rect -15788 29532 -9489 29548
rect -15788 29468 -9573 29532
rect -9509 29468 -9489 29532
rect -15788 29452 -9489 29468
rect -15788 29388 -9573 29452
rect -9509 29388 -9489 29452
rect -15788 29372 -9489 29388
rect -15788 29308 -9573 29372
rect -9509 29308 -9489 29372
rect -15788 29292 -9489 29308
rect -15788 29228 -9573 29292
rect -9509 29228 -9489 29292
rect -15788 29212 -9489 29228
rect -15788 29148 -9573 29212
rect -9509 29148 -9489 29212
rect -15788 29132 -9489 29148
rect -15788 29068 -9573 29132
rect -9509 29068 -9489 29132
rect -15788 29052 -9489 29068
rect -15788 28988 -9573 29052
rect -9509 28988 -9489 29052
rect -15788 28972 -9489 28988
rect -15788 28908 -9573 28972
rect -9509 28908 -9489 28972
rect -15788 28892 -9489 28908
rect -15788 28828 -9573 28892
rect -9509 28828 -9489 28892
rect -15788 28812 -9489 28828
rect -15788 28748 -9573 28812
rect -9509 28748 -9489 28812
rect -15788 28732 -9489 28748
rect -15788 28668 -9573 28732
rect -9509 28668 -9489 28732
rect -15788 28652 -9489 28668
rect -15788 28588 -9573 28652
rect -9509 28588 -9489 28652
rect -15788 28572 -9489 28588
rect -15788 28508 -9573 28572
rect -9509 28508 -9489 28572
rect -15788 28492 -9489 28508
rect -15788 28428 -9573 28492
rect -9509 28428 -9489 28492
rect -15788 28400 -9489 28428
rect -9469 34572 -3170 34600
rect -9469 34508 -3254 34572
rect -3190 34508 -3170 34572
rect -9469 34492 -3170 34508
rect -9469 34428 -3254 34492
rect -3190 34428 -3170 34492
rect -9469 34412 -3170 34428
rect -9469 34348 -3254 34412
rect -3190 34348 -3170 34412
rect -9469 34332 -3170 34348
rect -9469 34268 -3254 34332
rect -3190 34268 -3170 34332
rect -9469 34252 -3170 34268
rect -9469 34188 -3254 34252
rect -3190 34188 -3170 34252
rect -9469 34172 -3170 34188
rect -9469 34108 -3254 34172
rect -3190 34108 -3170 34172
rect -9469 34092 -3170 34108
rect -9469 34028 -3254 34092
rect -3190 34028 -3170 34092
rect -9469 34012 -3170 34028
rect -9469 33948 -3254 34012
rect -3190 33948 -3170 34012
rect -9469 33932 -3170 33948
rect -9469 33868 -3254 33932
rect -3190 33868 -3170 33932
rect -9469 33852 -3170 33868
rect -9469 33788 -3254 33852
rect -3190 33788 -3170 33852
rect -9469 33772 -3170 33788
rect -9469 33708 -3254 33772
rect -3190 33708 -3170 33772
rect -9469 33692 -3170 33708
rect -9469 33628 -3254 33692
rect -3190 33628 -3170 33692
rect -9469 33612 -3170 33628
rect -9469 33548 -3254 33612
rect -3190 33548 -3170 33612
rect -9469 33532 -3170 33548
rect -9469 33468 -3254 33532
rect -3190 33468 -3170 33532
rect -9469 33452 -3170 33468
rect -9469 33388 -3254 33452
rect -3190 33388 -3170 33452
rect -9469 33372 -3170 33388
rect -9469 33308 -3254 33372
rect -3190 33308 -3170 33372
rect -9469 33292 -3170 33308
rect -9469 33228 -3254 33292
rect -3190 33228 -3170 33292
rect -9469 33212 -3170 33228
rect -9469 33148 -3254 33212
rect -3190 33148 -3170 33212
rect -9469 33132 -3170 33148
rect -9469 33068 -3254 33132
rect -3190 33068 -3170 33132
rect -9469 33052 -3170 33068
rect -9469 32988 -3254 33052
rect -3190 32988 -3170 33052
rect -9469 32972 -3170 32988
rect -9469 32908 -3254 32972
rect -3190 32908 -3170 32972
rect -9469 32892 -3170 32908
rect -9469 32828 -3254 32892
rect -3190 32828 -3170 32892
rect -9469 32812 -3170 32828
rect -9469 32748 -3254 32812
rect -3190 32748 -3170 32812
rect -9469 32732 -3170 32748
rect -9469 32668 -3254 32732
rect -3190 32668 -3170 32732
rect -9469 32652 -3170 32668
rect -9469 32588 -3254 32652
rect -3190 32588 -3170 32652
rect -9469 32572 -3170 32588
rect -9469 32508 -3254 32572
rect -3190 32508 -3170 32572
rect -9469 32492 -3170 32508
rect -9469 32428 -3254 32492
rect -3190 32428 -3170 32492
rect -9469 32412 -3170 32428
rect -9469 32348 -3254 32412
rect -3190 32348 -3170 32412
rect -9469 32332 -3170 32348
rect -9469 32268 -3254 32332
rect -3190 32268 -3170 32332
rect -9469 32252 -3170 32268
rect -9469 32188 -3254 32252
rect -3190 32188 -3170 32252
rect -9469 32172 -3170 32188
rect -9469 32108 -3254 32172
rect -3190 32108 -3170 32172
rect -9469 32092 -3170 32108
rect -9469 32028 -3254 32092
rect -3190 32028 -3170 32092
rect -9469 32012 -3170 32028
rect -9469 31948 -3254 32012
rect -3190 31948 -3170 32012
rect -9469 31932 -3170 31948
rect -9469 31868 -3254 31932
rect -3190 31868 -3170 31932
rect -9469 31852 -3170 31868
rect -9469 31788 -3254 31852
rect -3190 31788 -3170 31852
rect -9469 31772 -3170 31788
rect -9469 31708 -3254 31772
rect -3190 31708 -3170 31772
rect -9469 31692 -3170 31708
rect -9469 31628 -3254 31692
rect -3190 31628 -3170 31692
rect -9469 31612 -3170 31628
rect -9469 31548 -3254 31612
rect -3190 31548 -3170 31612
rect -9469 31532 -3170 31548
rect -9469 31468 -3254 31532
rect -3190 31468 -3170 31532
rect -9469 31452 -3170 31468
rect -9469 31388 -3254 31452
rect -3190 31388 -3170 31452
rect -9469 31372 -3170 31388
rect -9469 31308 -3254 31372
rect -3190 31308 -3170 31372
rect -9469 31292 -3170 31308
rect -9469 31228 -3254 31292
rect -3190 31228 -3170 31292
rect -9469 31212 -3170 31228
rect -9469 31148 -3254 31212
rect -3190 31148 -3170 31212
rect -9469 31132 -3170 31148
rect -9469 31068 -3254 31132
rect -3190 31068 -3170 31132
rect -9469 31052 -3170 31068
rect -9469 30988 -3254 31052
rect -3190 30988 -3170 31052
rect -9469 30972 -3170 30988
rect -9469 30908 -3254 30972
rect -3190 30908 -3170 30972
rect -9469 30892 -3170 30908
rect -9469 30828 -3254 30892
rect -3190 30828 -3170 30892
rect -9469 30812 -3170 30828
rect -9469 30748 -3254 30812
rect -3190 30748 -3170 30812
rect -9469 30732 -3170 30748
rect -9469 30668 -3254 30732
rect -3190 30668 -3170 30732
rect -9469 30652 -3170 30668
rect -9469 30588 -3254 30652
rect -3190 30588 -3170 30652
rect -9469 30572 -3170 30588
rect -9469 30508 -3254 30572
rect -3190 30508 -3170 30572
rect -9469 30492 -3170 30508
rect -9469 30428 -3254 30492
rect -3190 30428 -3170 30492
rect -9469 30412 -3170 30428
rect -9469 30348 -3254 30412
rect -3190 30348 -3170 30412
rect -9469 30332 -3170 30348
rect -9469 30268 -3254 30332
rect -3190 30268 -3170 30332
rect -9469 30252 -3170 30268
rect -9469 30188 -3254 30252
rect -3190 30188 -3170 30252
rect -9469 30172 -3170 30188
rect -9469 30108 -3254 30172
rect -3190 30108 -3170 30172
rect -9469 30092 -3170 30108
rect -9469 30028 -3254 30092
rect -3190 30028 -3170 30092
rect -9469 30012 -3170 30028
rect -9469 29948 -3254 30012
rect -3190 29948 -3170 30012
rect -9469 29932 -3170 29948
rect -9469 29868 -3254 29932
rect -3190 29868 -3170 29932
rect -9469 29852 -3170 29868
rect -9469 29788 -3254 29852
rect -3190 29788 -3170 29852
rect -9469 29772 -3170 29788
rect -9469 29708 -3254 29772
rect -3190 29708 -3170 29772
rect -9469 29692 -3170 29708
rect -9469 29628 -3254 29692
rect -3190 29628 -3170 29692
rect -9469 29612 -3170 29628
rect -9469 29548 -3254 29612
rect -3190 29548 -3170 29612
rect -9469 29532 -3170 29548
rect -9469 29468 -3254 29532
rect -3190 29468 -3170 29532
rect -9469 29452 -3170 29468
rect -9469 29388 -3254 29452
rect -3190 29388 -3170 29452
rect -9469 29372 -3170 29388
rect -9469 29308 -3254 29372
rect -3190 29308 -3170 29372
rect -9469 29292 -3170 29308
rect -9469 29228 -3254 29292
rect -3190 29228 -3170 29292
rect -9469 29212 -3170 29228
rect -9469 29148 -3254 29212
rect -3190 29148 -3170 29212
rect -9469 29132 -3170 29148
rect -9469 29068 -3254 29132
rect -3190 29068 -3170 29132
rect -9469 29052 -3170 29068
rect -9469 28988 -3254 29052
rect -3190 28988 -3170 29052
rect -9469 28972 -3170 28988
rect -9469 28908 -3254 28972
rect -3190 28908 -3170 28972
rect -9469 28892 -3170 28908
rect -9469 28828 -3254 28892
rect -3190 28828 -3170 28892
rect -9469 28812 -3170 28828
rect -9469 28748 -3254 28812
rect -3190 28748 -3170 28812
rect -9469 28732 -3170 28748
rect -9469 28668 -3254 28732
rect -3190 28668 -3170 28732
rect -9469 28652 -3170 28668
rect -9469 28588 -3254 28652
rect -3190 28588 -3170 28652
rect -9469 28572 -3170 28588
rect -9469 28508 -3254 28572
rect -3190 28508 -3170 28572
rect -9469 28492 -3170 28508
rect -9469 28428 -3254 28492
rect -3190 28428 -3170 28492
rect -9469 28400 -3170 28428
rect -3150 34572 3149 34600
rect -3150 34508 3065 34572
rect 3129 34508 3149 34572
rect -3150 34492 3149 34508
rect -3150 34428 3065 34492
rect 3129 34428 3149 34492
rect -3150 34412 3149 34428
rect -3150 34348 3065 34412
rect 3129 34348 3149 34412
rect -3150 34332 3149 34348
rect -3150 34268 3065 34332
rect 3129 34268 3149 34332
rect -3150 34252 3149 34268
rect -3150 34188 3065 34252
rect 3129 34188 3149 34252
rect -3150 34172 3149 34188
rect -3150 34108 3065 34172
rect 3129 34108 3149 34172
rect -3150 34092 3149 34108
rect -3150 34028 3065 34092
rect 3129 34028 3149 34092
rect -3150 34012 3149 34028
rect -3150 33948 3065 34012
rect 3129 33948 3149 34012
rect -3150 33932 3149 33948
rect -3150 33868 3065 33932
rect 3129 33868 3149 33932
rect -3150 33852 3149 33868
rect -3150 33788 3065 33852
rect 3129 33788 3149 33852
rect -3150 33772 3149 33788
rect -3150 33708 3065 33772
rect 3129 33708 3149 33772
rect -3150 33692 3149 33708
rect -3150 33628 3065 33692
rect 3129 33628 3149 33692
rect -3150 33612 3149 33628
rect -3150 33548 3065 33612
rect 3129 33548 3149 33612
rect -3150 33532 3149 33548
rect -3150 33468 3065 33532
rect 3129 33468 3149 33532
rect -3150 33452 3149 33468
rect -3150 33388 3065 33452
rect 3129 33388 3149 33452
rect -3150 33372 3149 33388
rect -3150 33308 3065 33372
rect 3129 33308 3149 33372
rect -3150 33292 3149 33308
rect -3150 33228 3065 33292
rect 3129 33228 3149 33292
rect -3150 33212 3149 33228
rect -3150 33148 3065 33212
rect 3129 33148 3149 33212
rect -3150 33132 3149 33148
rect -3150 33068 3065 33132
rect 3129 33068 3149 33132
rect -3150 33052 3149 33068
rect -3150 32988 3065 33052
rect 3129 32988 3149 33052
rect -3150 32972 3149 32988
rect -3150 32908 3065 32972
rect 3129 32908 3149 32972
rect -3150 32892 3149 32908
rect -3150 32828 3065 32892
rect 3129 32828 3149 32892
rect -3150 32812 3149 32828
rect -3150 32748 3065 32812
rect 3129 32748 3149 32812
rect -3150 32732 3149 32748
rect -3150 32668 3065 32732
rect 3129 32668 3149 32732
rect -3150 32652 3149 32668
rect -3150 32588 3065 32652
rect 3129 32588 3149 32652
rect -3150 32572 3149 32588
rect -3150 32508 3065 32572
rect 3129 32508 3149 32572
rect -3150 32492 3149 32508
rect -3150 32428 3065 32492
rect 3129 32428 3149 32492
rect -3150 32412 3149 32428
rect -3150 32348 3065 32412
rect 3129 32348 3149 32412
rect -3150 32332 3149 32348
rect -3150 32268 3065 32332
rect 3129 32268 3149 32332
rect -3150 32252 3149 32268
rect -3150 32188 3065 32252
rect 3129 32188 3149 32252
rect -3150 32172 3149 32188
rect -3150 32108 3065 32172
rect 3129 32108 3149 32172
rect -3150 32092 3149 32108
rect -3150 32028 3065 32092
rect 3129 32028 3149 32092
rect -3150 32012 3149 32028
rect -3150 31948 3065 32012
rect 3129 31948 3149 32012
rect -3150 31932 3149 31948
rect -3150 31868 3065 31932
rect 3129 31868 3149 31932
rect -3150 31852 3149 31868
rect -3150 31788 3065 31852
rect 3129 31788 3149 31852
rect -3150 31772 3149 31788
rect -3150 31708 3065 31772
rect 3129 31708 3149 31772
rect -3150 31692 3149 31708
rect -3150 31628 3065 31692
rect 3129 31628 3149 31692
rect -3150 31612 3149 31628
rect -3150 31548 3065 31612
rect 3129 31548 3149 31612
rect -3150 31532 3149 31548
rect -3150 31468 3065 31532
rect 3129 31468 3149 31532
rect -3150 31452 3149 31468
rect -3150 31388 3065 31452
rect 3129 31388 3149 31452
rect -3150 31372 3149 31388
rect -3150 31308 3065 31372
rect 3129 31308 3149 31372
rect -3150 31292 3149 31308
rect -3150 31228 3065 31292
rect 3129 31228 3149 31292
rect -3150 31212 3149 31228
rect -3150 31148 3065 31212
rect 3129 31148 3149 31212
rect -3150 31132 3149 31148
rect -3150 31068 3065 31132
rect 3129 31068 3149 31132
rect -3150 31052 3149 31068
rect -3150 30988 3065 31052
rect 3129 30988 3149 31052
rect -3150 30972 3149 30988
rect -3150 30908 3065 30972
rect 3129 30908 3149 30972
rect -3150 30892 3149 30908
rect -3150 30828 3065 30892
rect 3129 30828 3149 30892
rect -3150 30812 3149 30828
rect -3150 30748 3065 30812
rect 3129 30748 3149 30812
rect -3150 30732 3149 30748
rect -3150 30668 3065 30732
rect 3129 30668 3149 30732
rect -3150 30652 3149 30668
rect -3150 30588 3065 30652
rect 3129 30588 3149 30652
rect -3150 30572 3149 30588
rect -3150 30508 3065 30572
rect 3129 30508 3149 30572
rect -3150 30492 3149 30508
rect -3150 30428 3065 30492
rect 3129 30428 3149 30492
rect -3150 30412 3149 30428
rect -3150 30348 3065 30412
rect 3129 30348 3149 30412
rect -3150 30332 3149 30348
rect -3150 30268 3065 30332
rect 3129 30268 3149 30332
rect -3150 30252 3149 30268
rect -3150 30188 3065 30252
rect 3129 30188 3149 30252
rect -3150 30172 3149 30188
rect -3150 30108 3065 30172
rect 3129 30108 3149 30172
rect -3150 30092 3149 30108
rect -3150 30028 3065 30092
rect 3129 30028 3149 30092
rect -3150 30012 3149 30028
rect -3150 29948 3065 30012
rect 3129 29948 3149 30012
rect -3150 29932 3149 29948
rect -3150 29868 3065 29932
rect 3129 29868 3149 29932
rect -3150 29852 3149 29868
rect -3150 29788 3065 29852
rect 3129 29788 3149 29852
rect -3150 29772 3149 29788
rect -3150 29708 3065 29772
rect 3129 29708 3149 29772
rect -3150 29692 3149 29708
rect -3150 29628 3065 29692
rect 3129 29628 3149 29692
rect -3150 29612 3149 29628
rect -3150 29548 3065 29612
rect 3129 29548 3149 29612
rect -3150 29532 3149 29548
rect -3150 29468 3065 29532
rect 3129 29468 3149 29532
rect -3150 29452 3149 29468
rect -3150 29388 3065 29452
rect 3129 29388 3149 29452
rect -3150 29372 3149 29388
rect -3150 29308 3065 29372
rect 3129 29308 3149 29372
rect -3150 29292 3149 29308
rect -3150 29228 3065 29292
rect 3129 29228 3149 29292
rect -3150 29212 3149 29228
rect -3150 29148 3065 29212
rect 3129 29148 3149 29212
rect -3150 29132 3149 29148
rect -3150 29068 3065 29132
rect 3129 29068 3149 29132
rect -3150 29052 3149 29068
rect -3150 28988 3065 29052
rect 3129 28988 3149 29052
rect -3150 28972 3149 28988
rect -3150 28908 3065 28972
rect 3129 28908 3149 28972
rect -3150 28892 3149 28908
rect -3150 28828 3065 28892
rect 3129 28828 3149 28892
rect -3150 28812 3149 28828
rect -3150 28748 3065 28812
rect 3129 28748 3149 28812
rect -3150 28732 3149 28748
rect -3150 28668 3065 28732
rect 3129 28668 3149 28732
rect -3150 28652 3149 28668
rect -3150 28588 3065 28652
rect 3129 28588 3149 28652
rect -3150 28572 3149 28588
rect -3150 28508 3065 28572
rect 3129 28508 3149 28572
rect -3150 28492 3149 28508
rect -3150 28428 3065 28492
rect 3129 28428 3149 28492
rect -3150 28400 3149 28428
rect 3169 34572 9468 34600
rect 3169 34508 9384 34572
rect 9448 34508 9468 34572
rect 3169 34492 9468 34508
rect 3169 34428 9384 34492
rect 9448 34428 9468 34492
rect 3169 34412 9468 34428
rect 3169 34348 9384 34412
rect 9448 34348 9468 34412
rect 3169 34332 9468 34348
rect 3169 34268 9384 34332
rect 9448 34268 9468 34332
rect 3169 34252 9468 34268
rect 3169 34188 9384 34252
rect 9448 34188 9468 34252
rect 3169 34172 9468 34188
rect 3169 34108 9384 34172
rect 9448 34108 9468 34172
rect 3169 34092 9468 34108
rect 3169 34028 9384 34092
rect 9448 34028 9468 34092
rect 3169 34012 9468 34028
rect 3169 33948 9384 34012
rect 9448 33948 9468 34012
rect 3169 33932 9468 33948
rect 3169 33868 9384 33932
rect 9448 33868 9468 33932
rect 3169 33852 9468 33868
rect 3169 33788 9384 33852
rect 9448 33788 9468 33852
rect 3169 33772 9468 33788
rect 3169 33708 9384 33772
rect 9448 33708 9468 33772
rect 3169 33692 9468 33708
rect 3169 33628 9384 33692
rect 9448 33628 9468 33692
rect 3169 33612 9468 33628
rect 3169 33548 9384 33612
rect 9448 33548 9468 33612
rect 3169 33532 9468 33548
rect 3169 33468 9384 33532
rect 9448 33468 9468 33532
rect 3169 33452 9468 33468
rect 3169 33388 9384 33452
rect 9448 33388 9468 33452
rect 3169 33372 9468 33388
rect 3169 33308 9384 33372
rect 9448 33308 9468 33372
rect 3169 33292 9468 33308
rect 3169 33228 9384 33292
rect 9448 33228 9468 33292
rect 3169 33212 9468 33228
rect 3169 33148 9384 33212
rect 9448 33148 9468 33212
rect 3169 33132 9468 33148
rect 3169 33068 9384 33132
rect 9448 33068 9468 33132
rect 3169 33052 9468 33068
rect 3169 32988 9384 33052
rect 9448 32988 9468 33052
rect 3169 32972 9468 32988
rect 3169 32908 9384 32972
rect 9448 32908 9468 32972
rect 3169 32892 9468 32908
rect 3169 32828 9384 32892
rect 9448 32828 9468 32892
rect 3169 32812 9468 32828
rect 3169 32748 9384 32812
rect 9448 32748 9468 32812
rect 3169 32732 9468 32748
rect 3169 32668 9384 32732
rect 9448 32668 9468 32732
rect 3169 32652 9468 32668
rect 3169 32588 9384 32652
rect 9448 32588 9468 32652
rect 3169 32572 9468 32588
rect 3169 32508 9384 32572
rect 9448 32508 9468 32572
rect 3169 32492 9468 32508
rect 3169 32428 9384 32492
rect 9448 32428 9468 32492
rect 3169 32412 9468 32428
rect 3169 32348 9384 32412
rect 9448 32348 9468 32412
rect 3169 32332 9468 32348
rect 3169 32268 9384 32332
rect 9448 32268 9468 32332
rect 3169 32252 9468 32268
rect 3169 32188 9384 32252
rect 9448 32188 9468 32252
rect 3169 32172 9468 32188
rect 3169 32108 9384 32172
rect 9448 32108 9468 32172
rect 3169 32092 9468 32108
rect 3169 32028 9384 32092
rect 9448 32028 9468 32092
rect 3169 32012 9468 32028
rect 3169 31948 9384 32012
rect 9448 31948 9468 32012
rect 3169 31932 9468 31948
rect 3169 31868 9384 31932
rect 9448 31868 9468 31932
rect 3169 31852 9468 31868
rect 3169 31788 9384 31852
rect 9448 31788 9468 31852
rect 3169 31772 9468 31788
rect 3169 31708 9384 31772
rect 9448 31708 9468 31772
rect 3169 31692 9468 31708
rect 3169 31628 9384 31692
rect 9448 31628 9468 31692
rect 3169 31612 9468 31628
rect 3169 31548 9384 31612
rect 9448 31548 9468 31612
rect 3169 31532 9468 31548
rect 3169 31468 9384 31532
rect 9448 31468 9468 31532
rect 3169 31452 9468 31468
rect 3169 31388 9384 31452
rect 9448 31388 9468 31452
rect 3169 31372 9468 31388
rect 3169 31308 9384 31372
rect 9448 31308 9468 31372
rect 3169 31292 9468 31308
rect 3169 31228 9384 31292
rect 9448 31228 9468 31292
rect 3169 31212 9468 31228
rect 3169 31148 9384 31212
rect 9448 31148 9468 31212
rect 3169 31132 9468 31148
rect 3169 31068 9384 31132
rect 9448 31068 9468 31132
rect 3169 31052 9468 31068
rect 3169 30988 9384 31052
rect 9448 30988 9468 31052
rect 3169 30972 9468 30988
rect 3169 30908 9384 30972
rect 9448 30908 9468 30972
rect 3169 30892 9468 30908
rect 3169 30828 9384 30892
rect 9448 30828 9468 30892
rect 3169 30812 9468 30828
rect 3169 30748 9384 30812
rect 9448 30748 9468 30812
rect 3169 30732 9468 30748
rect 3169 30668 9384 30732
rect 9448 30668 9468 30732
rect 3169 30652 9468 30668
rect 3169 30588 9384 30652
rect 9448 30588 9468 30652
rect 3169 30572 9468 30588
rect 3169 30508 9384 30572
rect 9448 30508 9468 30572
rect 3169 30492 9468 30508
rect 3169 30428 9384 30492
rect 9448 30428 9468 30492
rect 3169 30412 9468 30428
rect 3169 30348 9384 30412
rect 9448 30348 9468 30412
rect 3169 30332 9468 30348
rect 3169 30268 9384 30332
rect 9448 30268 9468 30332
rect 3169 30252 9468 30268
rect 3169 30188 9384 30252
rect 9448 30188 9468 30252
rect 3169 30172 9468 30188
rect 3169 30108 9384 30172
rect 9448 30108 9468 30172
rect 3169 30092 9468 30108
rect 3169 30028 9384 30092
rect 9448 30028 9468 30092
rect 3169 30012 9468 30028
rect 3169 29948 9384 30012
rect 9448 29948 9468 30012
rect 3169 29932 9468 29948
rect 3169 29868 9384 29932
rect 9448 29868 9468 29932
rect 3169 29852 9468 29868
rect 3169 29788 9384 29852
rect 9448 29788 9468 29852
rect 3169 29772 9468 29788
rect 3169 29708 9384 29772
rect 9448 29708 9468 29772
rect 3169 29692 9468 29708
rect 3169 29628 9384 29692
rect 9448 29628 9468 29692
rect 3169 29612 9468 29628
rect 3169 29548 9384 29612
rect 9448 29548 9468 29612
rect 3169 29532 9468 29548
rect 3169 29468 9384 29532
rect 9448 29468 9468 29532
rect 3169 29452 9468 29468
rect 3169 29388 9384 29452
rect 9448 29388 9468 29452
rect 3169 29372 9468 29388
rect 3169 29308 9384 29372
rect 9448 29308 9468 29372
rect 3169 29292 9468 29308
rect 3169 29228 9384 29292
rect 9448 29228 9468 29292
rect 3169 29212 9468 29228
rect 3169 29148 9384 29212
rect 9448 29148 9468 29212
rect 3169 29132 9468 29148
rect 3169 29068 9384 29132
rect 9448 29068 9468 29132
rect 3169 29052 9468 29068
rect 3169 28988 9384 29052
rect 9448 28988 9468 29052
rect 3169 28972 9468 28988
rect 3169 28908 9384 28972
rect 9448 28908 9468 28972
rect 3169 28892 9468 28908
rect 3169 28828 9384 28892
rect 9448 28828 9468 28892
rect 3169 28812 9468 28828
rect 3169 28748 9384 28812
rect 9448 28748 9468 28812
rect 3169 28732 9468 28748
rect 3169 28668 9384 28732
rect 9448 28668 9468 28732
rect 3169 28652 9468 28668
rect 3169 28588 9384 28652
rect 9448 28588 9468 28652
rect 3169 28572 9468 28588
rect 3169 28508 9384 28572
rect 9448 28508 9468 28572
rect 3169 28492 9468 28508
rect 3169 28428 9384 28492
rect 9448 28428 9468 28492
rect 3169 28400 9468 28428
rect 9488 34572 15787 34600
rect 9488 34508 15703 34572
rect 15767 34508 15787 34572
rect 9488 34492 15787 34508
rect 9488 34428 15703 34492
rect 15767 34428 15787 34492
rect 9488 34412 15787 34428
rect 9488 34348 15703 34412
rect 15767 34348 15787 34412
rect 9488 34332 15787 34348
rect 9488 34268 15703 34332
rect 15767 34268 15787 34332
rect 9488 34252 15787 34268
rect 9488 34188 15703 34252
rect 15767 34188 15787 34252
rect 9488 34172 15787 34188
rect 9488 34108 15703 34172
rect 15767 34108 15787 34172
rect 9488 34092 15787 34108
rect 9488 34028 15703 34092
rect 15767 34028 15787 34092
rect 9488 34012 15787 34028
rect 9488 33948 15703 34012
rect 15767 33948 15787 34012
rect 9488 33932 15787 33948
rect 9488 33868 15703 33932
rect 15767 33868 15787 33932
rect 9488 33852 15787 33868
rect 9488 33788 15703 33852
rect 15767 33788 15787 33852
rect 9488 33772 15787 33788
rect 9488 33708 15703 33772
rect 15767 33708 15787 33772
rect 9488 33692 15787 33708
rect 9488 33628 15703 33692
rect 15767 33628 15787 33692
rect 9488 33612 15787 33628
rect 9488 33548 15703 33612
rect 15767 33548 15787 33612
rect 9488 33532 15787 33548
rect 9488 33468 15703 33532
rect 15767 33468 15787 33532
rect 9488 33452 15787 33468
rect 9488 33388 15703 33452
rect 15767 33388 15787 33452
rect 9488 33372 15787 33388
rect 9488 33308 15703 33372
rect 15767 33308 15787 33372
rect 9488 33292 15787 33308
rect 9488 33228 15703 33292
rect 15767 33228 15787 33292
rect 9488 33212 15787 33228
rect 9488 33148 15703 33212
rect 15767 33148 15787 33212
rect 9488 33132 15787 33148
rect 9488 33068 15703 33132
rect 15767 33068 15787 33132
rect 9488 33052 15787 33068
rect 9488 32988 15703 33052
rect 15767 32988 15787 33052
rect 9488 32972 15787 32988
rect 9488 32908 15703 32972
rect 15767 32908 15787 32972
rect 9488 32892 15787 32908
rect 9488 32828 15703 32892
rect 15767 32828 15787 32892
rect 9488 32812 15787 32828
rect 9488 32748 15703 32812
rect 15767 32748 15787 32812
rect 9488 32732 15787 32748
rect 9488 32668 15703 32732
rect 15767 32668 15787 32732
rect 9488 32652 15787 32668
rect 9488 32588 15703 32652
rect 15767 32588 15787 32652
rect 9488 32572 15787 32588
rect 9488 32508 15703 32572
rect 15767 32508 15787 32572
rect 9488 32492 15787 32508
rect 9488 32428 15703 32492
rect 15767 32428 15787 32492
rect 9488 32412 15787 32428
rect 9488 32348 15703 32412
rect 15767 32348 15787 32412
rect 9488 32332 15787 32348
rect 9488 32268 15703 32332
rect 15767 32268 15787 32332
rect 9488 32252 15787 32268
rect 9488 32188 15703 32252
rect 15767 32188 15787 32252
rect 9488 32172 15787 32188
rect 9488 32108 15703 32172
rect 15767 32108 15787 32172
rect 9488 32092 15787 32108
rect 9488 32028 15703 32092
rect 15767 32028 15787 32092
rect 9488 32012 15787 32028
rect 9488 31948 15703 32012
rect 15767 31948 15787 32012
rect 9488 31932 15787 31948
rect 9488 31868 15703 31932
rect 15767 31868 15787 31932
rect 9488 31852 15787 31868
rect 9488 31788 15703 31852
rect 15767 31788 15787 31852
rect 9488 31772 15787 31788
rect 9488 31708 15703 31772
rect 15767 31708 15787 31772
rect 9488 31692 15787 31708
rect 9488 31628 15703 31692
rect 15767 31628 15787 31692
rect 9488 31612 15787 31628
rect 9488 31548 15703 31612
rect 15767 31548 15787 31612
rect 9488 31532 15787 31548
rect 9488 31468 15703 31532
rect 15767 31468 15787 31532
rect 9488 31452 15787 31468
rect 9488 31388 15703 31452
rect 15767 31388 15787 31452
rect 9488 31372 15787 31388
rect 9488 31308 15703 31372
rect 15767 31308 15787 31372
rect 9488 31292 15787 31308
rect 9488 31228 15703 31292
rect 15767 31228 15787 31292
rect 9488 31212 15787 31228
rect 9488 31148 15703 31212
rect 15767 31148 15787 31212
rect 9488 31132 15787 31148
rect 9488 31068 15703 31132
rect 15767 31068 15787 31132
rect 9488 31052 15787 31068
rect 9488 30988 15703 31052
rect 15767 30988 15787 31052
rect 9488 30972 15787 30988
rect 9488 30908 15703 30972
rect 15767 30908 15787 30972
rect 9488 30892 15787 30908
rect 9488 30828 15703 30892
rect 15767 30828 15787 30892
rect 9488 30812 15787 30828
rect 9488 30748 15703 30812
rect 15767 30748 15787 30812
rect 9488 30732 15787 30748
rect 9488 30668 15703 30732
rect 15767 30668 15787 30732
rect 9488 30652 15787 30668
rect 9488 30588 15703 30652
rect 15767 30588 15787 30652
rect 9488 30572 15787 30588
rect 9488 30508 15703 30572
rect 15767 30508 15787 30572
rect 9488 30492 15787 30508
rect 9488 30428 15703 30492
rect 15767 30428 15787 30492
rect 9488 30412 15787 30428
rect 9488 30348 15703 30412
rect 15767 30348 15787 30412
rect 9488 30332 15787 30348
rect 9488 30268 15703 30332
rect 15767 30268 15787 30332
rect 9488 30252 15787 30268
rect 9488 30188 15703 30252
rect 15767 30188 15787 30252
rect 9488 30172 15787 30188
rect 9488 30108 15703 30172
rect 15767 30108 15787 30172
rect 9488 30092 15787 30108
rect 9488 30028 15703 30092
rect 15767 30028 15787 30092
rect 9488 30012 15787 30028
rect 9488 29948 15703 30012
rect 15767 29948 15787 30012
rect 9488 29932 15787 29948
rect 9488 29868 15703 29932
rect 15767 29868 15787 29932
rect 9488 29852 15787 29868
rect 9488 29788 15703 29852
rect 15767 29788 15787 29852
rect 9488 29772 15787 29788
rect 9488 29708 15703 29772
rect 15767 29708 15787 29772
rect 9488 29692 15787 29708
rect 9488 29628 15703 29692
rect 15767 29628 15787 29692
rect 9488 29612 15787 29628
rect 9488 29548 15703 29612
rect 15767 29548 15787 29612
rect 9488 29532 15787 29548
rect 9488 29468 15703 29532
rect 15767 29468 15787 29532
rect 9488 29452 15787 29468
rect 9488 29388 15703 29452
rect 15767 29388 15787 29452
rect 9488 29372 15787 29388
rect 9488 29308 15703 29372
rect 15767 29308 15787 29372
rect 9488 29292 15787 29308
rect 9488 29228 15703 29292
rect 15767 29228 15787 29292
rect 9488 29212 15787 29228
rect 9488 29148 15703 29212
rect 15767 29148 15787 29212
rect 9488 29132 15787 29148
rect 9488 29068 15703 29132
rect 15767 29068 15787 29132
rect 9488 29052 15787 29068
rect 9488 28988 15703 29052
rect 15767 28988 15787 29052
rect 9488 28972 15787 28988
rect 9488 28908 15703 28972
rect 15767 28908 15787 28972
rect 9488 28892 15787 28908
rect 9488 28828 15703 28892
rect 15767 28828 15787 28892
rect 9488 28812 15787 28828
rect 9488 28748 15703 28812
rect 15767 28748 15787 28812
rect 9488 28732 15787 28748
rect 9488 28668 15703 28732
rect 15767 28668 15787 28732
rect 9488 28652 15787 28668
rect 9488 28588 15703 28652
rect 15767 28588 15787 28652
rect 9488 28572 15787 28588
rect 9488 28508 15703 28572
rect 15767 28508 15787 28572
rect 9488 28492 15787 28508
rect 9488 28428 15703 28492
rect 15767 28428 15787 28492
rect 9488 28400 15787 28428
rect 15807 34572 22106 34600
rect 15807 34508 22022 34572
rect 22086 34508 22106 34572
rect 15807 34492 22106 34508
rect 15807 34428 22022 34492
rect 22086 34428 22106 34492
rect 15807 34412 22106 34428
rect 15807 34348 22022 34412
rect 22086 34348 22106 34412
rect 15807 34332 22106 34348
rect 15807 34268 22022 34332
rect 22086 34268 22106 34332
rect 15807 34252 22106 34268
rect 15807 34188 22022 34252
rect 22086 34188 22106 34252
rect 15807 34172 22106 34188
rect 15807 34108 22022 34172
rect 22086 34108 22106 34172
rect 15807 34092 22106 34108
rect 15807 34028 22022 34092
rect 22086 34028 22106 34092
rect 15807 34012 22106 34028
rect 15807 33948 22022 34012
rect 22086 33948 22106 34012
rect 15807 33932 22106 33948
rect 15807 33868 22022 33932
rect 22086 33868 22106 33932
rect 15807 33852 22106 33868
rect 15807 33788 22022 33852
rect 22086 33788 22106 33852
rect 15807 33772 22106 33788
rect 15807 33708 22022 33772
rect 22086 33708 22106 33772
rect 15807 33692 22106 33708
rect 15807 33628 22022 33692
rect 22086 33628 22106 33692
rect 15807 33612 22106 33628
rect 15807 33548 22022 33612
rect 22086 33548 22106 33612
rect 15807 33532 22106 33548
rect 15807 33468 22022 33532
rect 22086 33468 22106 33532
rect 15807 33452 22106 33468
rect 15807 33388 22022 33452
rect 22086 33388 22106 33452
rect 15807 33372 22106 33388
rect 15807 33308 22022 33372
rect 22086 33308 22106 33372
rect 15807 33292 22106 33308
rect 15807 33228 22022 33292
rect 22086 33228 22106 33292
rect 15807 33212 22106 33228
rect 15807 33148 22022 33212
rect 22086 33148 22106 33212
rect 15807 33132 22106 33148
rect 15807 33068 22022 33132
rect 22086 33068 22106 33132
rect 15807 33052 22106 33068
rect 15807 32988 22022 33052
rect 22086 32988 22106 33052
rect 15807 32972 22106 32988
rect 15807 32908 22022 32972
rect 22086 32908 22106 32972
rect 15807 32892 22106 32908
rect 15807 32828 22022 32892
rect 22086 32828 22106 32892
rect 15807 32812 22106 32828
rect 15807 32748 22022 32812
rect 22086 32748 22106 32812
rect 15807 32732 22106 32748
rect 15807 32668 22022 32732
rect 22086 32668 22106 32732
rect 15807 32652 22106 32668
rect 15807 32588 22022 32652
rect 22086 32588 22106 32652
rect 15807 32572 22106 32588
rect 15807 32508 22022 32572
rect 22086 32508 22106 32572
rect 15807 32492 22106 32508
rect 15807 32428 22022 32492
rect 22086 32428 22106 32492
rect 15807 32412 22106 32428
rect 15807 32348 22022 32412
rect 22086 32348 22106 32412
rect 15807 32332 22106 32348
rect 15807 32268 22022 32332
rect 22086 32268 22106 32332
rect 15807 32252 22106 32268
rect 15807 32188 22022 32252
rect 22086 32188 22106 32252
rect 15807 32172 22106 32188
rect 15807 32108 22022 32172
rect 22086 32108 22106 32172
rect 15807 32092 22106 32108
rect 15807 32028 22022 32092
rect 22086 32028 22106 32092
rect 15807 32012 22106 32028
rect 15807 31948 22022 32012
rect 22086 31948 22106 32012
rect 15807 31932 22106 31948
rect 15807 31868 22022 31932
rect 22086 31868 22106 31932
rect 15807 31852 22106 31868
rect 15807 31788 22022 31852
rect 22086 31788 22106 31852
rect 15807 31772 22106 31788
rect 15807 31708 22022 31772
rect 22086 31708 22106 31772
rect 15807 31692 22106 31708
rect 15807 31628 22022 31692
rect 22086 31628 22106 31692
rect 15807 31612 22106 31628
rect 15807 31548 22022 31612
rect 22086 31548 22106 31612
rect 15807 31532 22106 31548
rect 15807 31468 22022 31532
rect 22086 31468 22106 31532
rect 15807 31452 22106 31468
rect 15807 31388 22022 31452
rect 22086 31388 22106 31452
rect 15807 31372 22106 31388
rect 15807 31308 22022 31372
rect 22086 31308 22106 31372
rect 15807 31292 22106 31308
rect 15807 31228 22022 31292
rect 22086 31228 22106 31292
rect 15807 31212 22106 31228
rect 15807 31148 22022 31212
rect 22086 31148 22106 31212
rect 15807 31132 22106 31148
rect 15807 31068 22022 31132
rect 22086 31068 22106 31132
rect 15807 31052 22106 31068
rect 15807 30988 22022 31052
rect 22086 30988 22106 31052
rect 15807 30972 22106 30988
rect 15807 30908 22022 30972
rect 22086 30908 22106 30972
rect 15807 30892 22106 30908
rect 15807 30828 22022 30892
rect 22086 30828 22106 30892
rect 15807 30812 22106 30828
rect 15807 30748 22022 30812
rect 22086 30748 22106 30812
rect 15807 30732 22106 30748
rect 15807 30668 22022 30732
rect 22086 30668 22106 30732
rect 15807 30652 22106 30668
rect 15807 30588 22022 30652
rect 22086 30588 22106 30652
rect 15807 30572 22106 30588
rect 15807 30508 22022 30572
rect 22086 30508 22106 30572
rect 15807 30492 22106 30508
rect 15807 30428 22022 30492
rect 22086 30428 22106 30492
rect 15807 30412 22106 30428
rect 15807 30348 22022 30412
rect 22086 30348 22106 30412
rect 15807 30332 22106 30348
rect 15807 30268 22022 30332
rect 22086 30268 22106 30332
rect 15807 30252 22106 30268
rect 15807 30188 22022 30252
rect 22086 30188 22106 30252
rect 15807 30172 22106 30188
rect 15807 30108 22022 30172
rect 22086 30108 22106 30172
rect 15807 30092 22106 30108
rect 15807 30028 22022 30092
rect 22086 30028 22106 30092
rect 15807 30012 22106 30028
rect 15807 29948 22022 30012
rect 22086 29948 22106 30012
rect 15807 29932 22106 29948
rect 15807 29868 22022 29932
rect 22086 29868 22106 29932
rect 15807 29852 22106 29868
rect 15807 29788 22022 29852
rect 22086 29788 22106 29852
rect 15807 29772 22106 29788
rect 15807 29708 22022 29772
rect 22086 29708 22106 29772
rect 15807 29692 22106 29708
rect 15807 29628 22022 29692
rect 22086 29628 22106 29692
rect 15807 29612 22106 29628
rect 15807 29548 22022 29612
rect 22086 29548 22106 29612
rect 15807 29532 22106 29548
rect 15807 29468 22022 29532
rect 22086 29468 22106 29532
rect 15807 29452 22106 29468
rect 15807 29388 22022 29452
rect 22086 29388 22106 29452
rect 15807 29372 22106 29388
rect 15807 29308 22022 29372
rect 22086 29308 22106 29372
rect 15807 29292 22106 29308
rect 15807 29228 22022 29292
rect 22086 29228 22106 29292
rect 15807 29212 22106 29228
rect 15807 29148 22022 29212
rect 22086 29148 22106 29212
rect 15807 29132 22106 29148
rect 15807 29068 22022 29132
rect 22086 29068 22106 29132
rect 15807 29052 22106 29068
rect 15807 28988 22022 29052
rect 22086 28988 22106 29052
rect 15807 28972 22106 28988
rect 15807 28908 22022 28972
rect 22086 28908 22106 28972
rect 15807 28892 22106 28908
rect 15807 28828 22022 28892
rect 22086 28828 22106 28892
rect 15807 28812 22106 28828
rect 15807 28748 22022 28812
rect 22086 28748 22106 28812
rect 15807 28732 22106 28748
rect 15807 28668 22022 28732
rect 22086 28668 22106 28732
rect 15807 28652 22106 28668
rect 15807 28588 22022 28652
rect 22086 28588 22106 28652
rect 15807 28572 22106 28588
rect 15807 28508 22022 28572
rect 22086 28508 22106 28572
rect 15807 28492 22106 28508
rect 15807 28428 22022 28492
rect 22086 28428 22106 28492
rect 15807 28400 22106 28428
rect 22126 34572 28425 34600
rect 22126 34508 28341 34572
rect 28405 34508 28425 34572
rect 22126 34492 28425 34508
rect 22126 34428 28341 34492
rect 28405 34428 28425 34492
rect 22126 34412 28425 34428
rect 22126 34348 28341 34412
rect 28405 34348 28425 34412
rect 22126 34332 28425 34348
rect 22126 34268 28341 34332
rect 28405 34268 28425 34332
rect 22126 34252 28425 34268
rect 22126 34188 28341 34252
rect 28405 34188 28425 34252
rect 22126 34172 28425 34188
rect 22126 34108 28341 34172
rect 28405 34108 28425 34172
rect 22126 34092 28425 34108
rect 22126 34028 28341 34092
rect 28405 34028 28425 34092
rect 22126 34012 28425 34028
rect 22126 33948 28341 34012
rect 28405 33948 28425 34012
rect 22126 33932 28425 33948
rect 22126 33868 28341 33932
rect 28405 33868 28425 33932
rect 22126 33852 28425 33868
rect 22126 33788 28341 33852
rect 28405 33788 28425 33852
rect 22126 33772 28425 33788
rect 22126 33708 28341 33772
rect 28405 33708 28425 33772
rect 22126 33692 28425 33708
rect 22126 33628 28341 33692
rect 28405 33628 28425 33692
rect 22126 33612 28425 33628
rect 22126 33548 28341 33612
rect 28405 33548 28425 33612
rect 22126 33532 28425 33548
rect 22126 33468 28341 33532
rect 28405 33468 28425 33532
rect 22126 33452 28425 33468
rect 22126 33388 28341 33452
rect 28405 33388 28425 33452
rect 22126 33372 28425 33388
rect 22126 33308 28341 33372
rect 28405 33308 28425 33372
rect 22126 33292 28425 33308
rect 22126 33228 28341 33292
rect 28405 33228 28425 33292
rect 22126 33212 28425 33228
rect 22126 33148 28341 33212
rect 28405 33148 28425 33212
rect 22126 33132 28425 33148
rect 22126 33068 28341 33132
rect 28405 33068 28425 33132
rect 22126 33052 28425 33068
rect 22126 32988 28341 33052
rect 28405 32988 28425 33052
rect 22126 32972 28425 32988
rect 22126 32908 28341 32972
rect 28405 32908 28425 32972
rect 22126 32892 28425 32908
rect 22126 32828 28341 32892
rect 28405 32828 28425 32892
rect 22126 32812 28425 32828
rect 22126 32748 28341 32812
rect 28405 32748 28425 32812
rect 22126 32732 28425 32748
rect 22126 32668 28341 32732
rect 28405 32668 28425 32732
rect 22126 32652 28425 32668
rect 22126 32588 28341 32652
rect 28405 32588 28425 32652
rect 22126 32572 28425 32588
rect 22126 32508 28341 32572
rect 28405 32508 28425 32572
rect 22126 32492 28425 32508
rect 22126 32428 28341 32492
rect 28405 32428 28425 32492
rect 22126 32412 28425 32428
rect 22126 32348 28341 32412
rect 28405 32348 28425 32412
rect 22126 32332 28425 32348
rect 22126 32268 28341 32332
rect 28405 32268 28425 32332
rect 22126 32252 28425 32268
rect 22126 32188 28341 32252
rect 28405 32188 28425 32252
rect 22126 32172 28425 32188
rect 22126 32108 28341 32172
rect 28405 32108 28425 32172
rect 22126 32092 28425 32108
rect 22126 32028 28341 32092
rect 28405 32028 28425 32092
rect 22126 32012 28425 32028
rect 22126 31948 28341 32012
rect 28405 31948 28425 32012
rect 22126 31932 28425 31948
rect 22126 31868 28341 31932
rect 28405 31868 28425 31932
rect 22126 31852 28425 31868
rect 22126 31788 28341 31852
rect 28405 31788 28425 31852
rect 22126 31772 28425 31788
rect 22126 31708 28341 31772
rect 28405 31708 28425 31772
rect 22126 31692 28425 31708
rect 22126 31628 28341 31692
rect 28405 31628 28425 31692
rect 22126 31612 28425 31628
rect 22126 31548 28341 31612
rect 28405 31548 28425 31612
rect 22126 31532 28425 31548
rect 22126 31468 28341 31532
rect 28405 31468 28425 31532
rect 22126 31452 28425 31468
rect 22126 31388 28341 31452
rect 28405 31388 28425 31452
rect 22126 31372 28425 31388
rect 22126 31308 28341 31372
rect 28405 31308 28425 31372
rect 22126 31292 28425 31308
rect 22126 31228 28341 31292
rect 28405 31228 28425 31292
rect 22126 31212 28425 31228
rect 22126 31148 28341 31212
rect 28405 31148 28425 31212
rect 22126 31132 28425 31148
rect 22126 31068 28341 31132
rect 28405 31068 28425 31132
rect 22126 31052 28425 31068
rect 22126 30988 28341 31052
rect 28405 30988 28425 31052
rect 22126 30972 28425 30988
rect 22126 30908 28341 30972
rect 28405 30908 28425 30972
rect 22126 30892 28425 30908
rect 22126 30828 28341 30892
rect 28405 30828 28425 30892
rect 22126 30812 28425 30828
rect 22126 30748 28341 30812
rect 28405 30748 28425 30812
rect 22126 30732 28425 30748
rect 22126 30668 28341 30732
rect 28405 30668 28425 30732
rect 22126 30652 28425 30668
rect 22126 30588 28341 30652
rect 28405 30588 28425 30652
rect 22126 30572 28425 30588
rect 22126 30508 28341 30572
rect 28405 30508 28425 30572
rect 22126 30492 28425 30508
rect 22126 30428 28341 30492
rect 28405 30428 28425 30492
rect 22126 30412 28425 30428
rect 22126 30348 28341 30412
rect 28405 30348 28425 30412
rect 22126 30332 28425 30348
rect 22126 30268 28341 30332
rect 28405 30268 28425 30332
rect 22126 30252 28425 30268
rect 22126 30188 28341 30252
rect 28405 30188 28425 30252
rect 22126 30172 28425 30188
rect 22126 30108 28341 30172
rect 28405 30108 28425 30172
rect 22126 30092 28425 30108
rect 22126 30028 28341 30092
rect 28405 30028 28425 30092
rect 22126 30012 28425 30028
rect 22126 29948 28341 30012
rect 28405 29948 28425 30012
rect 22126 29932 28425 29948
rect 22126 29868 28341 29932
rect 28405 29868 28425 29932
rect 22126 29852 28425 29868
rect 22126 29788 28341 29852
rect 28405 29788 28425 29852
rect 22126 29772 28425 29788
rect 22126 29708 28341 29772
rect 28405 29708 28425 29772
rect 22126 29692 28425 29708
rect 22126 29628 28341 29692
rect 28405 29628 28425 29692
rect 22126 29612 28425 29628
rect 22126 29548 28341 29612
rect 28405 29548 28425 29612
rect 22126 29532 28425 29548
rect 22126 29468 28341 29532
rect 28405 29468 28425 29532
rect 22126 29452 28425 29468
rect 22126 29388 28341 29452
rect 28405 29388 28425 29452
rect 22126 29372 28425 29388
rect 22126 29308 28341 29372
rect 28405 29308 28425 29372
rect 22126 29292 28425 29308
rect 22126 29228 28341 29292
rect 28405 29228 28425 29292
rect 22126 29212 28425 29228
rect 22126 29148 28341 29212
rect 28405 29148 28425 29212
rect 22126 29132 28425 29148
rect 22126 29068 28341 29132
rect 28405 29068 28425 29132
rect 22126 29052 28425 29068
rect 22126 28988 28341 29052
rect 28405 28988 28425 29052
rect 22126 28972 28425 28988
rect 22126 28908 28341 28972
rect 28405 28908 28425 28972
rect 22126 28892 28425 28908
rect 22126 28828 28341 28892
rect 28405 28828 28425 28892
rect 22126 28812 28425 28828
rect 22126 28748 28341 28812
rect 28405 28748 28425 28812
rect 22126 28732 28425 28748
rect 22126 28668 28341 28732
rect 28405 28668 28425 28732
rect 22126 28652 28425 28668
rect 22126 28588 28341 28652
rect 28405 28588 28425 28652
rect 22126 28572 28425 28588
rect 22126 28508 28341 28572
rect 28405 28508 28425 28572
rect 22126 28492 28425 28508
rect 22126 28428 28341 28492
rect 28405 28428 28425 28492
rect 22126 28400 28425 28428
rect 28445 34572 34744 34600
rect 28445 34508 34660 34572
rect 34724 34508 34744 34572
rect 28445 34492 34744 34508
rect 28445 34428 34660 34492
rect 34724 34428 34744 34492
rect 28445 34412 34744 34428
rect 28445 34348 34660 34412
rect 34724 34348 34744 34412
rect 28445 34332 34744 34348
rect 28445 34268 34660 34332
rect 34724 34268 34744 34332
rect 28445 34252 34744 34268
rect 28445 34188 34660 34252
rect 34724 34188 34744 34252
rect 28445 34172 34744 34188
rect 28445 34108 34660 34172
rect 34724 34108 34744 34172
rect 28445 34092 34744 34108
rect 28445 34028 34660 34092
rect 34724 34028 34744 34092
rect 28445 34012 34744 34028
rect 28445 33948 34660 34012
rect 34724 33948 34744 34012
rect 28445 33932 34744 33948
rect 28445 33868 34660 33932
rect 34724 33868 34744 33932
rect 28445 33852 34744 33868
rect 28445 33788 34660 33852
rect 34724 33788 34744 33852
rect 28445 33772 34744 33788
rect 28445 33708 34660 33772
rect 34724 33708 34744 33772
rect 28445 33692 34744 33708
rect 28445 33628 34660 33692
rect 34724 33628 34744 33692
rect 28445 33612 34744 33628
rect 28445 33548 34660 33612
rect 34724 33548 34744 33612
rect 28445 33532 34744 33548
rect 28445 33468 34660 33532
rect 34724 33468 34744 33532
rect 28445 33452 34744 33468
rect 28445 33388 34660 33452
rect 34724 33388 34744 33452
rect 28445 33372 34744 33388
rect 28445 33308 34660 33372
rect 34724 33308 34744 33372
rect 28445 33292 34744 33308
rect 28445 33228 34660 33292
rect 34724 33228 34744 33292
rect 28445 33212 34744 33228
rect 28445 33148 34660 33212
rect 34724 33148 34744 33212
rect 28445 33132 34744 33148
rect 28445 33068 34660 33132
rect 34724 33068 34744 33132
rect 28445 33052 34744 33068
rect 28445 32988 34660 33052
rect 34724 32988 34744 33052
rect 28445 32972 34744 32988
rect 28445 32908 34660 32972
rect 34724 32908 34744 32972
rect 28445 32892 34744 32908
rect 28445 32828 34660 32892
rect 34724 32828 34744 32892
rect 28445 32812 34744 32828
rect 28445 32748 34660 32812
rect 34724 32748 34744 32812
rect 28445 32732 34744 32748
rect 28445 32668 34660 32732
rect 34724 32668 34744 32732
rect 28445 32652 34744 32668
rect 28445 32588 34660 32652
rect 34724 32588 34744 32652
rect 28445 32572 34744 32588
rect 28445 32508 34660 32572
rect 34724 32508 34744 32572
rect 28445 32492 34744 32508
rect 28445 32428 34660 32492
rect 34724 32428 34744 32492
rect 28445 32412 34744 32428
rect 28445 32348 34660 32412
rect 34724 32348 34744 32412
rect 28445 32332 34744 32348
rect 28445 32268 34660 32332
rect 34724 32268 34744 32332
rect 28445 32252 34744 32268
rect 28445 32188 34660 32252
rect 34724 32188 34744 32252
rect 28445 32172 34744 32188
rect 28445 32108 34660 32172
rect 34724 32108 34744 32172
rect 28445 32092 34744 32108
rect 28445 32028 34660 32092
rect 34724 32028 34744 32092
rect 28445 32012 34744 32028
rect 28445 31948 34660 32012
rect 34724 31948 34744 32012
rect 28445 31932 34744 31948
rect 28445 31868 34660 31932
rect 34724 31868 34744 31932
rect 28445 31852 34744 31868
rect 28445 31788 34660 31852
rect 34724 31788 34744 31852
rect 28445 31772 34744 31788
rect 28445 31708 34660 31772
rect 34724 31708 34744 31772
rect 28445 31692 34744 31708
rect 28445 31628 34660 31692
rect 34724 31628 34744 31692
rect 28445 31612 34744 31628
rect 28445 31548 34660 31612
rect 34724 31548 34744 31612
rect 28445 31532 34744 31548
rect 28445 31468 34660 31532
rect 34724 31468 34744 31532
rect 28445 31452 34744 31468
rect 28445 31388 34660 31452
rect 34724 31388 34744 31452
rect 28445 31372 34744 31388
rect 28445 31308 34660 31372
rect 34724 31308 34744 31372
rect 28445 31292 34744 31308
rect 28445 31228 34660 31292
rect 34724 31228 34744 31292
rect 28445 31212 34744 31228
rect 28445 31148 34660 31212
rect 34724 31148 34744 31212
rect 28445 31132 34744 31148
rect 28445 31068 34660 31132
rect 34724 31068 34744 31132
rect 28445 31052 34744 31068
rect 28445 30988 34660 31052
rect 34724 30988 34744 31052
rect 28445 30972 34744 30988
rect 28445 30908 34660 30972
rect 34724 30908 34744 30972
rect 28445 30892 34744 30908
rect 28445 30828 34660 30892
rect 34724 30828 34744 30892
rect 28445 30812 34744 30828
rect 28445 30748 34660 30812
rect 34724 30748 34744 30812
rect 28445 30732 34744 30748
rect 28445 30668 34660 30732
rect 34724 30668 34744 30732
rect 28445 30652 34744 30668
rect 28445 30588 34660 30652
rect 34724 30588 34744 30652
rect 28445 30572 34744 30588
rect 28445 30508 34660 30572
rect 34724 30508 34744 30572
rect 28445 30492 34744 30508
rect 28445 30428 34660 30492
rect 34724 30428 34744 30492
rect 28445 30412 34744 30428
rect 28445 30348 34660 30412
rect 34724 30348 34744 30412
rect 28445 30332 34744 30348
rect 28445 30268 34660 30332
rect 34724 30268 34744 30332
rect 28445 30252 34744 30268
rect 28445 30188 34660 30252
rect 34724 30188 34744 30252
rect 28445 30172 34744 30188
rect 28445 30108 34660 30172
rect 34724 30108 34744 30172
rect 28445 30092 34744 30108
rect 28445 30028 34660 30092
rect 34724 30028 34744 30092
rect 28445 30012 34744 30028
rect 28445 29948 34660 30012
rect 34724 29948 34744 30012
rect 28445 29932 34744 29948
rect 28445 29868 34660 29932
rect 34724 29868 34744 29932
rect 28445 29852 34744 29868
rect 28445 29788 34660 29852
rect 34724 29788 34744 29852
rect 28445 29772 34744 29788
rect 28445 29708 34660 29772
rect 34724 29708 34744 29772
rect 28445 29692 34744 29708
rect 28445 29628 34660 29692
rect 34724 29628 34744 29692
rect 28445 29612 34744 29628
rect 28445 29548 34660 29612
rect 34724 29548 34744 29612
rect 28445 29532 34744 29548
rect 28445 29468 34660 29532
rect 34724 29468 34744 29532
rect 28445 29452 34744 29468
rect 28445 29388 34660 29452
rect 34724 29388 34744 29452
rect 28445 29372 34744 29388
rect 28445 29308 34660 29372
rect 34724 29308 34744 29372
rect 28445 29292 34744 29308
rect 28445 29228 34660 29292
rect 34724 29228 34744 29292
rect 28445 29212 34744 29228
rect 28445 29148 34660 29212
rect 34724 29148 34744 29212
rect 28445 29132 34744 29148
rect 28445 29068 34660 29132
rect 34724 29068 34744 29132
rect 28445 29052 34744 29068
rect 28445 28988 34660 29052
rect 34724 28988 34744 29052
rect 28445 28972 34744 28988
rect 28445 28908 34660 28972
rect 34724 28908 34744 28972
rect 28445 28892 34744 28908
rect 28445 28828 34660 28892
rect 34724 28828 34744 28892
rect 28445 28812 34744 28828
rect 28445 28748 34660 28812
rect 34724 28748 34744 28812
rect 28445 28732 34744 28748
rect 28445 28668 34660 28732
rect 34724 28668 34744 28732
rect 28445 28652 34744 28668
rect 28445 28588 34660 28652
rect 34724 28588 34744 28652
rect 28445 28572 34744 28588
rect 28445 28508 34660 28572
rect 34724 28508 34744 28572
rect 28445 28492 34744 28508
rect 28445 28428 34660 28492
rect 34724 28428 34744 28492
rect 28445 28400 34744 28428
rect 34764 34572 41063 34600
rect 34764 34508 40979 34572
rect 41043 34508 41063 34572
rect 34764 34492 41063 34508
rect 34764 34428 40979 34492
rect 41043 34428 41063 34492
rect 34764 34412 41063 34428
rect 34764 34348 40979 34412
rect 41043 34348 41063 34412
rect 34764 34332 41063 34348
rect 34764 34268 40979 34332
rect 41043 34268 41063 34332
rect 34764 34252 41063 34268
rect 34764 34188 40979 34252
rect 41043 34188 41063 34252
rect 34764 34172 41063 34188
rect 34764 34108 40979 34172
rect 41043 34108 41063 34172
rect 34764 34092 41063 34108
rect 34764 34028 40979 34092
rect 41043 34028 41063 34092
rect 34764 34012 41063 34028
rect 34764 33948 40979 34012
rect 41043 33948 41063 34012
rect 34764 33932 41063 33948
rect 34764 33868 40979 33932
rect 41043 33868 41063 33932
rect 34764 33852 41063 33868
rect 34764 33788 40979 33852
rect 41043 33788 41063 33852
rect 34764 33772 41063 33788
rect 34764 33708 40979 33772
rect 41043 33708 41063 33772
rect 34764 33692 41063 33708
rect 34764 33628 40979 33692
rect 41043 33628 41063 33692
rect 34764 33612 41063 33628
rect 34764 33548 40979 33612
rect 41043 33548 41063 33612
rect 34764 33532 41063 33548
rect 34764 33468 40979 33532
rect 41043 33468 41063 33532
rect 34764 33452 41063 33468
rect 34764 33388 40979 33452
rect 41043 33388 41063 33452
rect 34764 33372 41063 33388
rect 34764 33308 40979 33372
rect 41043 33308 41063 33372
rect 34764 33292 41063 33308
rect 34764 33228 40979 33292
rect 41043 33228 41063 33292
rect 34764 33212 41063 33228
rect 34764 33148 40979 33212
rect 41043 33148 41063 33212
rect 34764 33132 41063 33148
rect 34764 33068 40979 33132
rect 41043 33068 41063 33132
rect 34764 33052 41063 33068
rect 34764 32988 40979 33052
rect 41043 32988 41063 33052
rect 34764 32972 41063 32988
rect 34764 32908 40979 32972
rect 41043 32908 41063 32972
rect 34764 32892 41063 32908
rect 34764 32828 40979 32892
rect 41043 32828 41063 32892
rect 34764 32812 41063 32828
rect 34764 32748 40979 32812
rect 41043 32748 41063 32812
rect 34764 32732 41063 32748
rect 34764 32668 40979 32732
rect 41043 32668 41063 32732
rect 34764 32652 41063 32668
rect 34764 32588 40979 32652
rect 41043 32588 41063 32652
rect 34764 32572 41063 32588
rect 34764 32508 40979 32572
rect 41043 32508 41063 32572
rect 34764 32492 41063 32508
rect 34764 32428 40979 32492
rect 41043 32428 41063 32492
rect 34764 32412 41063 32428
rect 34764 32348 40979 32412
rect 41043 32348 41063 32412
rect 34764 32332 41063 32348
rect 34764 32268 40979 32332
rect 41043 32268 41063 32332
rect 34764 32252 41063 32268
rect 34764 32188 40979 32252
rect 41043 32188 41063 32252
rect 34764 32172 41063 32188
rect 34764 32108 40979 32172
rect 41043 32108 41063 32172
rect 34764 32092 41063 32108
rect 34764 32028 40979 32092
rect 41043 32028 41063 32092
rect 34764 32012 41063 32028
rect 34764 31948 40979 32012
rect 41043 31948 41063 32012
rect 34764 31932 41063 31948
rect 34764 31868 40979 31932
rect 41043 31868 41063 31932
rect 34764 31852 41063 31868
rect 34764 31788 40979 31852
rect 41043 31788 41063 31852
rect 34764 31772 41063 31788
rect 34764 31708 40979 31772
rect 41043 31708 41063 31772
rect 34764 31692 41063 31708
rect 34764 31628 40979 31692
rect 41043 31628 41063 31692
rect 34764 31612 41063 31628
rect 34764 31548 40979 31612
rect 41043 31548 41063 31612
rect 34764 31532 41063 31548
rect 34764 31468 40979 31532
rect 41043 31468 41063 31532
rect 34764 31452 41063 31468
rect 34764 31388 40979 31452
rect 41043 31388 41063 31452
rect 34764 31372 41063 31388
rect 34764 31308 40979 31372
rect 41043 31308 41063 31372
rect 34764 31292 41063 31308
rect 34764 31228 40979 31292
rect 41043 31228 41063 31292
rect 34764 31212 41063 31228
rect 34764 31148 40979 31212
rect 41043 31148 41063 31212
rect 34764 31132 41063 31148
rect 34764 31068 40979 31132
rect 41043 31068 41063 31132
rect 34764 31052 41063 31068
rect 34764 30988 40979 31052
rect 41043 30988 41063 31052
rect 34764 30972 41063 30988
rect 34764 30908 40979 30972
rect 41043 30908 41063 30972
rect 34764 30892 41063 30908
rect 34764 30828 40979 30892
rect 41043 30828 41063 30892
rect 34764 30812 41063 30828
rect 34764 30748 40979 30812
rect 41043 30748 41063 30812
rect 34764 30732 41063 30748
rect 34764 30668 40979 30732
rect 41043 30668 41063 30732
rect 34764 30652 41063 30668
rect 34764 30588 40979 30652
rect 41043 30588 41063 30652
rect 34764 30572 41063 30588
rect 34764 30508 40979 30572
rect 41043 30508 41063 30572
rect 34764 30492 41063 30508
rect 34764 30428 40979 30492
rect 41043 30428 41063 30492
rect 34764 30412 41063 30428
rect 34764 30348 40979 30412
rect 41043 30348 41063 30412
rect 34764 30332 41063 30348
rect 34764 30268 40979 30332
rect 41043 30268 41063 30332
rect 34764 30252 41063 30268
rect 34764 30188 40979 30252
rect 41043 30188 41063 30252
rect 34764 30172 41063 30188
rect 34764 30108 40979 30172
rect 41043 30108 41063 30172
rect 34764 30092 41063 30108
rect 34764 30028 40979 30092
rect 41043 30028 41063 30092
rect 34764 30012 41063 30028
rect 34764 29948 40979 30012
rect 41043 29948 41063 30012
rect 34764 29932 41063 29948
rect 34764 29868 40979 29932
rect 41043 29868 41063 29932
rect 34764 29852 41063 29868
rect 34764 29788 40979 29852
rect 41043 29788 41063 29852
rect 34764 29772 41063 29788
rect 34764 29708 40979 29772
rect 41043 29708 41063 29772
rect 34764 29692 41063 29708
rect 34764 29628 40979 29692
rect 41043 29628 41063 29692
rect 34764 29612 41063 29628
rect 34764 29548 40979 29612
rect 41043 29548 41063 29612
rect 34764 29532 41063 29548
rect 34764 29468 40979 29532
rect 41043 29468 41063 29532
rect 34764 29452 41063 29468
rect 34764 29388 40979 29452
rect 41043 29388 41063 29452
rect 34764 29372 41063 29388
rect 34764 29308 40979 29372
rect 41043 29308 41063 29372
rect 34764 29292 41063 29308
rect 34764 29228 40979 29292
rect 41043 29228 41063 29292
rect 34764 29212 41063 29228
rect 34764 29148 40979 29212
rect 41043 29148 41063 29212
rect 34764 29132 41063 29148
rect 34764 29068 40979 29132
rect 41043 29068 41063 29132
rect 34764 29052 41063 29068
rect 34764 28988 40979 29052
rect 41043 28988 41063 29052
rect 34764 28972 41063 28988
rect 34764 28908 40979 28972
rect 41043 28908 41063 28972
rect 34764 28892 41063 28908
rect 34764 28828 40979 28892
rect 41043 28828 41063 28892
rect 34764 28812 41063 28828
rect 34764 28748 40979 28812
rect 41043 28748 41063 28812
rect 34764 28732 41063 28748
rect 34764 28668 40979 28732
rect 41043 28668 41063 28732
rect 34764 28652 41063 28668
rect 34764 28588 40979 28652
rect 41043 28588 41063 28652
rect 34764 28572 41063 28588
rect 34764 28508 40979 28572
rect 41043 28508 41063 28572
rect 34764 28492 41063 28508
rect 34764 28428 40979 28492
rect 41043 28428 41063 28492
rect 34764 28400 41063 28428
rect 41083 34572 47382 34600
rect 41083 34508 47298 34572
rect 47362 34508 47382 34572
rect 41083 34492 47382 34508
rect 41083 34428 47298 34492
rect 47362 34428 47382 34492
rect 41083 34412 47382 34428
rect 41083 34348 47298 34412
rect 47362 34348 47382 34412
rect 41083 34332 47382 34348
rect 41083 34268 47298 34332
rect 47362 34268 47382 34332
rect 41083 34252 47382 34268
rect 41083 34188 47298 34252
rect 47362 34188 47382 34252
rect 41083 34172 47382 34188
rect 41083 34108 47298 34172
rect 47362 34108 47382 34172
rect 41083 34092 47382 34108
rect 41083 34028 47298 34092
rect 47362 34028 47382 34092
rect 41083 34012 47382 34028
rect 41083 33948 47298 34012
rect 47362 33948 47382 34012
rect 41083 33932 47382 33948
rect 41083 33868 47298 33932
rect 47362 33868 47382 33932
rect 41083 33852 47382 33868
rect 41083 33788 47298 33852
rect 47362 33788 47382 33852
rect 41083 33772 47382 33788
rect 41083 33708 47298 33772
rect 47362 33708 47382 33772
rect 41083 33692 47382 33708
rect 41083 33628 47298 33692
rect 47362 33628 47382 33692
rect 41083 33612 47382 33628
rect 41083 33548 47298 33612
rect 47362 33548 47382 33612
rect 41083 33532 47382 33548
rect 41083 33468 47298 33532
rect 47362 33468 47382 33532
rect 41083 33452 47382 33468
rect 41083 33388 47298 33452
rect 47362 33388 47382 33452
rect 41083 33372 47382 33388
rect 41083 33308 47298 33372
rect 47362 33308 47382 33372
rect 41083 33292 47382 33308
rect 41083 33228 47298 33292
rect 47362 33228 47382 33292
rect 41083 33212 47382 33228
rect 41083 33148 47298 33212
rect 47362 33148 47382 33212
rect 41083 33132 47382 33148
rect 41083 33068 47298 33132
rect 47362 33068 47382 33132
rect 41083 33052 47382 33068
rect 41083 32988 47298 33052
rect 47362 32988 47382 33052
rect 41083 32972 47382 32988
rect 41083 32908 47298 32972
rect 47362 32908 47382 32972
rect 41083 32892 47382 32908
rect 41083 32828 47298 32892
rect 47362 32828 47382 32892
rect 41083 32812 47382 32828
rect 41083 32748 47298 32812
rect 47362 32748 47382 32812
rect 41083 32732 47382 32748
rect 41083 32668 47298 32732
rect 47362 32668 47382 32732
rect 41083 32652 47382 32668
rect 41083 32588 47298 32652
rect 47362 32588 47382 32652
rect 41083 32572 47382 32588
rect 41083 32508 47298 32572
rect 47362 32508 47382 32572
rect 41083 32492 47382 32508
rect 41083 32428 47298 32492
rect 47362 32428 47382 32492
rect 41083 32412 47382 32428
rect 41083 32348 47298 32412
rect 47362 32348 47382 32412
rect 41083 32332 47382 32348
rect 41083 32268 47298 32332
rect 47362 32268 47382 32332
rect 41083 32252 47382 32268
rect 41083 32188 47298 32252
rect 47362 32188 47382 32252
rect 41083 32172 47382 32188
rect 41083 32108 47298 32172
rect 47362 32108 47382 32172
rect 41083 32092 47382 32108
rect 41083 32028 47298 32092
rect 47362 32028 47382 32092
rect 41083 32012 47382 32028
rect 41083 31948 47298 32012
rect 47362 31948 47382 32012
rect 41083 31932 47382 31948
rect 41083 31868 47298 31932
rect 47362 31868 47382 31932
rect 41083 31852 47382 31868
rect 41083 31788 47298 31852
rect 47362 31788 47382 31852
rect 41083 31772 47382 31788
rect 41083 31708 47298 31772
rect 47362 31708 47382 31772
rect 41083 31692 47382 31708
rect 41083 31628 47298 31692
rect 47362 31628 47382 31692
rect 41083 31612 47382 31628
rect 41083 31548 47298 31612
rect 47362 31548 47382 31612
rect 41083 31532 47382 31548
rect 41083 31468 47298 31532
rect 47362 31468 47382 31532
rect 41083 31452 47382 31468
rect 41083 31388 47298 31452
rect 47362 31388 47382 31452
rect 41083 31372 47382 31388
rect 41083 31308 47298 31372
rect 47362 31308 47382 31372
rect 41083 31292 47382 31308
rect 41083 31228 47298 31292
rect 47362 31228 47382 31292
rect 41083 31212 47382 31228
rect 41083 31148 47298 31212
rect 47362 31148 47382 31212
rect 41083 31132 47382 31148
rect 41083 31068 47298 31132
rect 47362 31068 47382 31132
rect 41083 31052 47382 31068
rect 41083 30988 47298 31052
rect 47362 30988 47382 31052
rect 41083 30972 47382 30988
rect 41083 30908 47298 30972
rect 47362 30908 47382 30972
rect 41083 30892 47382 30908
rect 41083 30828 47298 30892
rect 47362 30828 47382 30892
rect 41083 30812 47382 30828
rect 41083 30748 47298 30812
rect 47362 30748 47382 30812
rect 41083 30732 47382 30748
rect 41083 30668 47298 30732
rect 47362 30668 47382 30732
rect 41083 30652 47382 30668
rect 41083 30588 47298 30652
rect 47362 30588 47382 30652
rect 41083 30572 47382 30588
rect 41083 30508 47298 30572
rect 47362 30508 47382 30572
rect 41083 30492 47382 30508
rect 41083 30428 47298 30492
rect 47362 30428 47382 30492
rect 41083 30412 47382 30428
rect 41083 30348 47298 30412
rect 47362 30348 47382 30412
rect 41083 30332 47382 30348
rect 41083 30268 47298 30332
rect 47362 30268 47382 30332
rect 41083 30252 47382 30268
rect 41083 30188 47298 30252
rect 47362 30188 47382 30252
rect 41083 30172 47382 30188
rect 41083 30108 47298 30172
rect 47362 30108 47382 30172
rect 41083 30092 47382 30108
rect 41083 30028 47298 30092
rect 47362 30028 47382 30092
rect 41083 30012 47382 30028
rect 41083 29948 47298 30012
rect 47362 29948 47382 30012
rect 41083 29932 47382 29948
rect 41083 29868 47298 29932
rect 47362 29868 47382 29932
rect 41083 29852 47382 29868
rect 41083 29788 47298 29852
rect 47362 29788 47382 29852
rect 41083 29772 47382 29788
rect 41083 29708 47298 29772
rect 47362 29708 47382 29772
rect 41083 29692 47382 29708
rect 41083 29628 47298 29692
rect 47362 29628 47382 29692
rect 41083 29612 47382 29628
rect 41083 29548 47298 29612
rect 47362 29548 47382 29612
rect 41083 29532 47382 29548
rect 41083 29468 47298 29532
rect 47362 29468 47382 29532
rect 41083 29452 47382 29468
rect 41083 29388 47298 29452
rect 47362 29388 47382 29452
rect 41083 29372 47382 29388
rect 41083 29308 47298 29372
rect 47362 29308 47382 29372
rect 41083 29292 47382 29308
rect 41083 29228 47298 29292
rect 47362 29228 47382 29292
rect 41083 29212 47382 29228
rect 41083 29148 47298 29212
rect 47362 29148 47382 29212
rect 41083 29132 47382 29148
rect 41083 29068 47298 29132
rect 47362 29068 47382 29132
rect 41083 29052 47382 29068
rect 41083 28988 47298 29052
rect 47362 28988 47382 29052
rect 41083 28972 47382 28988
rect 41083 28908 47298 28972
rect 47362 28908 47382 28972
rect 41083 28892 47382 28908
rect 41083 28828 47298 28892
rect 47362 28828 47382 28892
rect 41083 28812 47382 28828
rect 41083 28748 47298 28812
rect 47362 28748 47382 28812
rect 41083 28732 47382 28748
rect 41083 28668 47298 28732
rect 47362 28668 47382 28732
rect 41083 28652 47382 28668
rect 41083 28588 47298 28652
rect 47362 28588 47382 28652
rect 41083 28572 47382 28588
rect 41083 28508 47298 28572
rect 47362 28508 47382 28572
rect 41083 28492 47382 28508
rect 41083 28428 47298 28492
rect 47362 28428 47382 28492
rect 41083 28400 47382 28428
rect -47383 28272 -41084 28300
rect -47383 28208 -41168 28272
rect -41104 28208 -41084 28272
rect -47383 28192 -41084 28208
rect -47383 28128 -41168 28192
rect -41104 28128 -41084 28192
rect -47383 28112 -41084 28128
rect -47383 28048 -41168 28112
rect -41104 28048 -41084 28112
rect -47383 28032 -41084 28048
rect -47383 27968 -41168 28032
rect -41104 27968 -41084 28032
rect -47383 27952 -41084 27968
rect -47383 27888 -41168 27952
rect -41104 27888 -41084 27952
rect -47383 27872 -41084 27888
rect -47383 27808 -41168 27872
rect -41104 27808 -41084 27872
rect -47383 27792 -41084 27808
rect -47383 27728 -41168 27792
rect -41104 27728 -41084 27792
rect -47383 27712 -41084 27728
rect -47383 27648 -41168 27712
rect -41104 27648 -41084 27712
rect -47383 27632 -41084 27648
rect -47383 27568 -41168 27632
rect -41104 27568 -41084 27632
rect -47383 27552 -41084 27568
rect -47383 27488 -41168 27552
rect -41104 27488 -41084 27552
rect -47383 27472 -41084 27488
rect -47383 27408 -41168 27472
rect -41104 27408 -41084 27472
rect -47383 27392 -41084 27408
rect -47383 27328 -41168 27392
rect -41104 27328 -41084 27392
rect -47383 27312 -41084 27328
rect -47383 27248 -41168 27312
rect -41104 27248 -41084 27312
rect -47383 27232 -41084 27248
rect -47383 27168 -41168 27232
rect -41104 27168 -41084 27232
rect -47383 27152 -41084 27168
rect -47383 27088 -41168 27152
rect -41104 27088 -41084 27152
rect -47383 27072 -41084 27088
rect -47383 27008 -41168 27072
rect -41104 27008 -41084 27072
rect -47383 26992 -41084 27008
rect -47383 26928 -41168 26992
rect -41104 26928 -41084 26992
rect -47383 26912 -41084 26928
rect -47383 26848 -41168 26912
rect -41104 26848 -41084 26912
rect -47383 26832 -41084 26848
rect -47383 26768 -41168 26832
rect -41104 26768 -41084 26832
rect -47383 26752 -41084 26768
rect -47383 26688 -41168 26752
rect -41104 26688 -41084 26752
rect -47383 26672 -41084 26688
rect -47383 26608 -41168 26672
rect -41104 26608 -41084 26672
rect -47383 26592 -41084 26608
rect -47383 26528 -41168 26592
rect -41104 26528 -41084 26592
rect -47383 26512 -41084 26528
rect -47383 26448 -41168 26512
rect -41104 26448 -41084 26512
rect -47383 26432 -41084 26448
rect -47383 26368 -41168 26432
rect -41104 26368 -41084 26432
rect -47383 26352 -41084 26368
rect -47383 26288 -41168 26352
rect -41104 26288 -41084 26352
rect -47383 26272 -41084 26288
rect -47383 26208 -41168 26272
rect -41104 26208 -41084 26272
rect -47383 26192 -41084 26208
rect -47383 26128 -41168 26192
rect -41104 26128 -41084 26192
rect -47383 26112 -41084 26128
rect -47383 26048 -41168 26112
rect -41104 26048 -41084 26112
rect -47383 26032 -41084 26048
rect -47383 25968 -41168 26032
rect -41104 25968 -41084 26032
rect -47383 25952 -41084 25968
rect -47383 25888 -41168 25952
rect -41104 25888 -41084 25952
rect -47383 25872 -41084 25888
rect -47383 25808 -41168 25872
rect -41104 25808 -41084 25872
rect -47383 25792 -41084 25808
rect -47383 25728 -41168 25792
rect -41104 25728 -41084 25792
rect -47383 25712 -41084 25728
rect -47383 25648 -41168 25712
rect -41104 25648 -41084 25712
rect -47383 25632 -41084 25648
rect -47383 25568 -41168 25632
rect -41104 25568 -41084 25632
rect -47383 25552 -41084 25568
rect -47383 25488 -41168 25552
rect -41104 25488 -41084 25552
rect -47383 25472 -41084 25488
rect -47383 25408 -41168 25472
rect -41104 25408 -41084 25472
rect -47383 25392 -41084 25408
rect -47383 25328 -41168 25392
rect -41104 25328 -41084 25392
rect -47383 25312 -41084 25328
rect -47383 25248 -41168 25312
rect -41104 25248 -41084 25312
rect -47383 25232 -41084 25248
rect -47383 25168 -41168 25232
rect -41104 25168 -41084 25232
rect -47383 25152 -41084 25168
rect -47383 25088 -41168 25152
rect -41104 25088 -41084 25152
rect -47383 25072 -41084 25088
rect -47383 25008 -41168 25072
rect -41104 25008 -41084 25072
rect -47383 24992 -41084 25008
rect -47383 24928 -41168 24992
rect -41104 24928 -41084 24992
rect -47383 24912 -41084 24928
rect -47383 24848 -41168 24912
rect -41104 24848 -41084 24912
rect -47383 24832 -41084 24848
rect -47383 24768 -41168 24832
rect -41104 24768 -41084 24832
rect -47383 24752 -41084 24768
rect -47383 24688 -41168 24752
rect -41104 24688 -41084 24752
rect -47383 24672 -41084 24688
rect -47383 24608 -41168 24672
rect -41104 24608 -41084 24672
rect -47383 24592 -41084 24608
rect -47383 24528 -41168 24592
rect -41104 24528 -41084 24592
rect -47383 24512 -41084 24528
rect -47383 24448 -41168 24512
rect -41104 24448 -41084 24512
rect -47383 24432 -41084 24448
rect -47383 24368 -41168 24432
rect -41104 24368 -41084 24432
rect -47383 24352 -41084 24368
rect -47383 24288 -41168 24352
rect -41104 24288 -41084 24352
rect -47383 24272 -41084 24288
rect -47383 24208 -41168 24272
rect -41104 24208 -41084 24272
rect -47383 24192 -41084 24208
rect -47383 24128 -41168 24192
rect -41104 24128 -41084 24192
rect -47383 24112 -41084 24128
rect -47383 24048 -41168 24112
rect -41104 24048 -41084 24112
rect -47383 24032 -41084 24048
rect -47383 23968 -41168 24032
rect -41104 23968 -41084 24032
rect -47383 23952 -41084 23968
rect -47383 23888 -41168 23952
rect -41104 23888 -41084 23952
rect -47383 23872 -41084 23888
rect -47383 23808 -41168 23872
rect -41104 23808 -41084 23872
rect -47383 23792 -41084 23808
rect -47383 23728 -41168 23792
rect -41104 23728 -41084 23792
rect -47383 23712 -41084 23728
rect -47383 23648 -41168 23712
rect -41104 23648 -41084 23712
rect -47383 23632 -41084 23648
rect -47383 23568 -41168 23632
rect -41104 23568 -41084 23632
rect -47383 23552 -41084 23568
rect -47383 23488 -41168 23552
rect -41104 23488 -41084 23552
rect -47383 23472 -41084 23488
rect -47383 23408 -41168 23472
rect -41104 23408 -41084 23472
rect -47383 23392 -41084 23408
rect -47383 23328 -41168 23392
rect -41104 23328 -41084 23392
rect -47383 23312 -41084 23328
rect -47383 23248 -41168 23312
rect -41104 23248 -41084 23312
rect -47383 23232 -41084 23248
rect -47383 23168 -41168 23232
rect -41104 23168 -41084 23232
rect -47383 23152 -41084 23168
rect -47383 23088 -41168 23152
rect -41104 23088 -41084 23152
rect -47383 23072 -41084 23088
rect -47383 23008 -41168 23072
rect -41104 23008 -41084 23072
rect -47383 22992 -41084 23008
rect -47383 22928 -41168 22992
rect -41104 22928 -41084 22992
rect -47383 22912 -41084 22928
rect -47383 22848 -41168 22912
rect -41104 22848 -41084 22912
rect -47383 22832 -41084 22848
rect -47383 22768 -41168 22832
rect -41104 22768 -41084 22832
rect -47383 22752 -41084 22768
rect -47383 22688 -41168 22752
rect -41104 22688 -41084 22752
rect -47383 22672 -41084 22688
rect -47383 22608 -41168 22672
rect -41104 22608 -41084 22672
rect -47383 22592 -41084 22608
rect -47383 22528 -41168 22592
rect -41104 22528 -41084 22592
rect -47383 22512 -41084 22528
rect -47383 22448 -41168 22512
rect -41104 22448 -41084 22512
rect -47383 22432 -41084 22448
rect -47383 22368 -41168 22432
rect -41104 22368 -41084 22432
rect -47383 22352 -41084 22368
rect -47383 22288 -41168 22352
rect -41104 22288 -41084 22352
rect -47383 22272 -41084 22288
rect -47383 22208 -41168 22272
rect -41104 22208 -41084 22272
rect -47383 22192 -41084 22208
rect -47383 22128 -41168 22192
rect -41104 22128 -41084 22192
rect -47383 22100 -41084 22128
rect -41064 28272 -34765 28300
rect -41064 28208 -34849 28272
rect -34785 28208 -34765 28272
rect -41064 28192 -34765 28208
rect -41064 28128 -34849 28192
rect -34785 28128 -34765 28192
rect -41064 28112 -34765 28128
rect -41064 28048 -34849 28112
rect -34785 28048 -34765 28112
rect -41064 28032 -34765 28048
rect -41064 27968 -34849 28032
rect -34785 27968 -34765 28032
rect -41064 27952 -34765 27968
rect -41064 27888 -34849 27952
rect -34785 27888 -34765 27952
rect -41064 27872 -34765 27888
rect -41064 27808 -34849 27872
rect -34785 27808 -34765 27872
rect -41064 27792 -34765 27808
rect -41064 27728 -34849 27792
rect -34785 27728 -34765 27792
rect -41064 27712 -34765 27728
rect -41064 27648 -34849 27712
rect -34785 27648 -34765 27712
rect -41064 27632 -34765 27648
rect -41064 27568 -34849 27632
rect -34785 27568 -34765 27632
rect -41064 27552 -34765 27568
rect -41064 27488 -34849 27552
rect -34785 27488 -34765 27552
rect -41064 27472 -34765 27488
rect -41064 27408 -34849 27472
rect -34785 27408 -34765 27472
rect -41064 27392 -34765 27408
rect -41064 27328 -34849 27392
rect -34785 27328 -34765 27392
rect -41064 27312 -34765 27328
rect -41064 27248 -34849 27312
rect -34785 27248 -34765 27312
rect -41064 27232 -34765 27248
rect -41064 27168 -34849 27232
rect -34785 27168 -34765 27232
rect -41064 27152 -34765 27168
rect -41064 27088 -34849 27152
rect -34785 27088 -34765 27152
rect -41064 27072 -34765 27088
rect -41064 27008 -34849 27072
rect -34785 27008 -34765 27072
rect -41064 26992 -34765 27008
rect -41064 26928 -34849 26992
rect -34785 26928 -34765 26992
rect -41064 26912 -34765 26928
rect -41064 26848 -34849 26912
rect -34785 26848 -34765 26912
rect -41064 26832 -34765 26848
rect -41064 26768 -34849 26832
rect -34785 26768 -34765 26832
rect -41064 26752 -34765 26768
rect -41064 26688 -34849 26752
rect -34785 26688 -34765 26752
rect -41064 26672 -34765 26688
rect -41064 26608 -34849 26672
rect -34785 26608 -34765 26672
rect -41064 26592 -34765 26608
rect -41064 26528 -34849 26592
rect -34785 26528 -34765 26592
rect -41064 26512 -34765 26528
rect -41064 26448 -34849 26512
rect -34785 26448 -34765 26512
rect -41064 26432 -34765 26448
rect -41064 26368 -34849 26432
rect -34785 26368 -34765 26432
rect -41064 26352 -34765 26368
rect -41064 26288 -34849 26352
rect -34785 26288 -34765 26352
rect -41064 26272 -34765 26288
rect -41064 26208 -34849 26272
rect -34785 26208 -34765 26272
rect -41064 26192 -34765 26208
rect -41064 26128 -34849 26192
rect -34785 26128 -34765 26192
rect -41064 26112 -34765 26128
rect -41064 26048 -34849 26112
rect -34785 26048 -34765 26112
rect -41064 26032 -34765 26048
rect -41064 25968 -34849 26032
rect -34785 25968 -34765 26032
rect -41064 25952 -34765 25968
rect -41064 25888 -34849 25952
rect -34785 25888 -34765 25952
rect -41064 25872 -34765 25888
rect -41064 25808 -34849 25872
rect -34785 25808 -34765 25872
rect -41064 25792 -34765 25808
rect -41064 25728 -34849 25792
rect -34785 25728 -34765 25792
rect -41064 25712 -34765 25728
rect -41064 25648 -34849 25712
rect -34785 25648 -34765 25712
rect -41064 25632 -34765 25648
rect -41064 25568 -34849 25632
rect -34785 25568 -34765 25632
rect -41064 25552 -34765 25568
rect -41064 25488 -34849 25552
rect -34785 25488 -34765 25552
rect -41064 25472 -34765 25488
rect -41064 25408 -34849 25472
rect -34785 25408 -34765 25472
rect -41064 25392 -34765 25408
rect -41064 25328 -34849 25392
rect -34785 25328 -34765 25392
rect -41064 25312 -34765 25328
rect -41064 25248 -34849 25312
rect -34785 25248 -34765 25312
rect -41064 25232 -34765 25248
rect -41064 25168 -34849 25232
rect -34785 25168 -34765 25232
rect -41064 25152 -34765 25168
rect -41064 25088 -34849 25152
rect -34785 25088 -34765 25152
rect -41064 25072 -34765 25088
rect -41064 25008 -34849 25072
rect -34785 25008 -34765 25072
rect -41064 24992 -34765 25008
rect -41064 24928 -34849 24992
rect -34785 24928 -34765 24992
rect -41064 24912 -34765 24928
rect -41064 24848 -34849 24912
rect -34785 24848 -34765 24912
rect -41064 24832 -34765 24848
rect -41064 24768 -34849 24832
rect -34785 24768 -34765 24832
rect -41064 24752 -34765 24768
rect -41064 24688 -34849 24752
rect -34785 24688 -34765 24752
rect -41064 24672 -34765 24688
rect -41064 24608 -34849 24672
rect -34785 24608 -34765 24672
rect -41064 24592 -34765 24608
rect -41064 24528 -34849 24592
rect -34785 24528 -34765 24592
rect -41064 24512 -34765 24528
rect -41064 24448 -34849 24512
rect -34785 24448 -34765 24512
rect -41064 24432 -34765 24448
rect -41064 24368 -34849 24432
rect -34785 24368 -34765 24432
rect -41064 24352 -34765 24368
rect -41064 24288 -34849 24352
rect -34785 24288 -34765 24352
rect -41064 24272 -34765 24288
rect -41064 24208 -34849 24272
rect -34785 24208 -34765 24272
rect -41064 24192 -34765 24208
rect -41064 24128 -34849 24192
rect -34785 24128 -34765 24192
rect -41064 24112 -34765 24128
rect -41064 24048 -34849 24112
rect -34785 24048 -34765 24112
rect -41064 24032 -34765 24048
rect -41064 23968 -34849 24032
rect -34785 23968 -34765 24032
rect -41064 23952 -34765 23968
rect -41064 23888 -34849 23952
rect -34785 23888 -34765 23952
rect -41064 23872 -34765 23888
rect -41064 23808 -34849 23872
rect -34785 23808 -34765 23872
rect -41064 23792 -34765 23808
rect -41064 23728 -34849 23792
rect -34785 23728 -34765 23792
rect -41064 23712 -34765 23728
rect -41064 23648 -34849 23712
rect -34785 23648 -34765 23712
rect -41064 23632 -34765 23648
rect -41064 23568 -34849 23632
rect -34785 23568 -34765 23632
rect -41064 23552 -34765 23568
rect -41064 23488 -34849 23552
rect -34785 23488 -34765 23552
rect -41064 23472 -34765 23488
rect -41064 23408 -34849 23472
rect -34785 23408 -34765 23472
rect -41064 23392 -34765 23408
rect -41064 23328 -34849 23392
rect -34785 23328 -34765 23392
rect -41064 23312 -34765 23328
rect -41064 23248 -34849 23312
rect -34785 23248 -34765 23312
rect -41064 23232 -34765 23248
rect -41064 23168 -34849 23232
rect -34785 23168 -34765 23232
rect -41064 23152 -34765 23168
rect -41064 23088 -34849 23152
rect -34785 23088 -34765 23152
rect -41064 23072 -34765 23088
rect -41064 23008 -34849 23072
rect -34785 23008 -34765 23072
rect -41064 22992 -34765 23008
rect -41064 22928 -34849 22992
rect -34785 22928 -34765 22992
rect -41064 22912 -34765 22928
rect -41064 22848 -34849 22912
rect -34785 22848 -34765 22912
rect -41064 22832 -34765 22848
rect -41064 22768 -34849 22832
rect -34785 22768 -34765 22832
rect -41064 22752 -34765 22768
rect -41064 22688 -34849 22752
rect -34785 22688 -34765 22752
rect -41064 22672 -34765 22688
rect -41064 22608 -34849 22672
rect -34785 22608 -34765 22672
rect -41064 22592 -34765 22608
rect -41064 22528 -34849 22592
rect -34785 22528 -34765 22592
rect -41064 22512 -34765 22528
rect -41064 22448 -34849 22512
rect -34785 22448 -34765 22512
rect -41064 22432 -34765 22448
rect -41064 22368 -34849 22432
rect -34785 22368 -34765 22432
rect -41064 22352 -34765 22368
rect -41064 22288 -34849 22352
rect -34785 22288 -34765 22352
rect -41064 22272 -34765 22288
rect -41064 22208 -34849 22272
rect -34785 22208 -34765 22272
rect -41064 22192 -34765 22208
rect -41064 22128 -34849 22192
rect -34785 22128 -34765 22192
rect -41064 22100 -34765 22128
rect -34745 28272 -28446 28300
rect -34745 28208 -28530 28272
rect -28466 28208 -28446 28272
rect -34745 28192 -28446 28208
rect -34745 28128 -28530 28192
rect -28466 28128 -28446 28192
rect -34745 28112 -28446 28128
rect -34745 28048 -28530 28112
rect -28466 28048 -28446 28112
rect -34745 28032 -28446 28048
rect -34745 27968 -28530 28032
rect -28466 27968 -28446 28032
rect -34745 27952 -28446 27968
rect -34745 27888 -28530 27952
rect -28466 27888 -28446 27952
rect -34745 27872 -28446 27888
rect -34745 27808 -28530 27872
rect -28466 27808 -28446 27872
rect -34745 27792 -28446 27808
rect -34745 27728 -28530 27792
rect -28466 27728 -28446 27792
rect -34745 27712 -28446 27728
rect -34745 27648 -28530 27712
rect -28466 27648 -28446 27712
rect -34745 27632 -28446 27648
rect -34745 27568 -28530 27632
rect -28466 27568 -28446 27632
rect -34745 27552 -28446 27568
rect -34745 27488 -28530 27552
rect -28466 27488 -28446 27552
rect -34745 27472 -28446 27488
rect -34745 27408 -28530 27472
rect -28466 27408 -28446 27472
rect -34745 27392 -28446 27408
rect -34745 27328 -28530 27392
rect -28466 27328 -28446 27392
rect -34745 27312 -28446 27328
rect -34745 27248 -28530 27312
rect -28466 27248 -28446 27312
rect -34745 27232 -28446 27248
rect -34745 27168 -28530 27232
rect -28466 27168 -28446 27232
rect -34745 27152 -28446 27168
rect -34745 27088 -28530 27152
rect -28466 27088 -28446 27152
rect -34745 27072 -28446 27088
rect -34745 27008 -28530 27072
rect -28466 27008 -28446 27072
rect -34745 26992 -28446 27008
rect -34745 26928 -28530 26992
rect -28466 26928 -28446 26992
rect -34745 26912 -28446 26928
rect -34745 26848 -28530 26912
rect -28466 26848 -28446 26912
rect -34745 26832 -28446 26848
rect -34745 26768 -28530 26832
rect -28466 26768 -28446 26832
rect -34745 26752 -28446 26768
rect -34745 26688 -28530 26752
rect -28466 26688 -28446 26752
rect -34745 26672 -28446 26688
rect -34745 26608 -28530 26672
rect -28466 26608 -28446 26672
rect -34745 26592 -28446 26608
rect -34745 26528 -28530 26592
rect -28466 26528 -28446 26592
rect -34745 26512 -28446 26528
rect -34745 26448 -28530 26512
rect -28466 26448 -28446 26512
rect -34745 26432 -28446 26448
rect -34745 26368 -28530 26432
rect -28466 26368 -28446 26432
rect -34745 26352 -28446 26368
rect -34745 26288 -28530 26352
rect -28466 26288 -28446 26352
rect -34745 26272 -28446 26288
rect -34745 26208 -28530 26272
rect -28466 26208 -28446 26272
rect -34745 26192 -28446 26208
rect -34745 26128 -28530 26192
rect -28466 26128 -28446 26192
rect -34745 26112 -28446 26128
rect -34745 26048 -28530 26112
rect -28466 26048 -28446 26112
rect -34745 26032 -28446 26048
rect -34745 25968 -28530 26032
rect -28466 25968 -28446 26032
rect -34745 25952 -28446 25968
rect -34745 25888 -28530 25952
rect -28466 25888 -28446 25952
rect -34745 25872 -28446 25888
rect -34745 25808 -28530 25872
rect -28466 25808 -28446 25872
rect -34745 25792 -28446 25808
rect -34745 25728 -28530 25792
rect -28466 25728 -28446 25792
rect -34745 25712 -28446 25728
rect -34745 25648 -28530 25712
rect -28466 25648 -28446 25712
rect -34745 25632 -28446 25648
rect -34745 25568 -28530 25632
rect -28466 25568 -28446 25632
rect -34745 25552 -28446 25568
rect -34745 25488 -28530 25552
rect -28466 25488 -28446 25552
rect -34745 25472 -28446 25488
rect -34745 25408 -28530 25472
rect -28466 25408 -28446 25472
rect -34745 25392 -28446 25408
rect -34745 25328 -28530 25392
rect -28466 25328 -28446 25392
rect -34745 25312 -28446 25328
rect -34745 25248 -28530 25312
rect -28466 25248 -28446 25312
rect -34745 25232 -28446 25248
rect -34745 25168 -28530 25232
rect -28466 25168 -28446 25232
rect -34745 25152 -28446 25168
rect -34745 25088 -28530 25152
rect -28466 25088 -28446 25152
rect -34745 25072 -28446 25088
rect -34745 25008 -28530 25072
rect -28466 25008 -28446 25072
rect -34745 24992 -28446 25008
rect -34745 24928 -28530 24992
rect -28466 24928 -28446 24992
rect -34745 24912 -28446 24928
rect -34745 24848 -28530 24912
rect -28466 24848 -28446 24912
rect -34745 24832 -28446 24848
rect -34745 24768 -28530 24832
rect -28466 24768 -28446 24832
rect -34745 24752 -28446 24768
rect -34745 24688 -28530 24752
rect -28466 24688 -28446 24752
rect -34745 24672 -28446 24688
rect -34745 24608 -28530 24672
rect -28466 24608 -28446 24672
rect -34745 24592 -28446 24608
rect -34745 24528 -28530 24592
rect -28466 24528 -28446 24592
rect -34745 24512 -28446 24528
rect -34745 24448 -28530 24512
rect -28466 24448 -28446 24512
rect -34745 24432 -28446 24448
rect -34745 24368 -28530 24432
rect -28466 24368 -28446 24432
rect -34745 24352 -28446 24368
rect -34745 24288 -28530 24352
rect -28466 24288 -28446 24352
rect -34745 24272 -28446 24288
rect -34745 24208 -28530 24272
rect -28466 24208 -28446 24272
rect -34745 24192 -28446 24208
rect -34745 24128 -28530 24192
rect -28466 24128 -28446 24192
rect -34745 24112 -28446 24128
rect -34745 24048 -28530 24112
rect -28466 24048 -28446 24112
rect -34745 24032 -28446 24048
rect -34745 23968 -28530 24032
rect -28466 23968 -28446 24032
rect -34745 23952 -28446 23968
rect -34745 23888 -28530 23952
rect -28466 23888 -28446 23952
rect -34745 23872 -28446 23888
rect -34745 23808 -28530 23872
rect -28466 23808 -28446 23872
rect -34745 23792 -28446 23808
rect -34745 23728 -28530 23792
rect -28466 23728 -28446 23792
rect -34745 23712 -28446 23728
rect -34745 23648 -28530 23712
rect -28466 23648 -28446 23712
rect -34745 23632 -28446 23648
rect -34745 23568 -28530 23632
rect -28466 23568 -28446 23632
rect -34745 23552 -28446 23568
rect -34745 23488 -28530 23552
rect -28466 23488 -28446 23552
rect -34745 23472 -28446 23488
rect -34745 23408 -28530 23472
rect -28466 23408 -28446 23472
rect -34745 23392 -28446 23408
rect -34745 23328 -28530 23392
rect -28466 23328 -28446 23392
rect -34745 23312 -28446 23328
rect -34745 23248 -28530 23312
rect -28466 23248 -28446 23312
rect -34745 23232 -28446 23248
rect -34745 23168 -28530 23232
rect -28466 23168 -28446 23232
rect -34745 23152 -28446 23168
rect -34745 23088 -28530 23152
rect -28466 23088 -28446 23152
rect -34745 23072 -28446 23088
rect -34745 23008 -28530 23072
rect -28466 23008 -28446 23072
rect -34745 22992 -28446 23008
rect -34745 22928 -28530 22992
rect -28466 22928 -28446 22992
rect -34745 22912 -28446 22928
rect -34745 22848 -28530 22912
rect -28466 22848 -28446 22912
rect -34745 22832 -28446 22848
rect -34745 22768 -28530 22832
rect -28466 22768 -28446 22832
rect -34745 22752 -28446 22768
rect -34745 22688 -28530 22752
rect -28466 22688 -28446 22752
rect -34745 22672 -28446 22688
rect -34745 22608 -28530 22672
rect -28466 22608 -28446 22672
rect -34745 22592 -28446 22608
rect -34745 22528 -28530 22592
rect -28466 22528 -28446 22592
rect -34745 22512 -28446 22528
rect -34745 22448 -28530 22512
rect -28466 22448 -28446 22512
rect -34745 22432 -28446 22448
rect -34745 22368 -28530 22432
rect -28466 22368 -28446 22432
rect -34745 22352 -28446 22368
rect -34745 22288 -28530 22352
rect -28466 22288 -28446 22352
rect -34745 22272 -28446 22288
rect -34745 22208 -28530 22272
rect -28466 22208 -28446 22272
rect -34745 22192 -28446 22208
rect -34745 22128 -28530 22192
rect -28466 22128 -28446 22192
rect -34745 22100 -28446 22128
rect -28426 28272 -22127 28300
rect -28426 28208 -22211 28272
rect -22147 28208 -22127 28272
rect -28426 28192 -22127 28208
rect -28426 28128 -22211 28192
rect -22147 28128 -22127 28192
rect -28426 28112 -22127 28128
rect -28426 28048 -22211 28112
rect -22147 28048 -22127 28112
rect -28426 28032 -22127 28048
rect -28426 27968 -22211 28032
rect -22147 27968 -22127 28032
rect -28426 27952 -22127 27968
rect -28426 27888 -22211 27952
rect -22147 27888 -22127 27952
rect -28426 27872 -22127 27888
rect -28426 27808 -22211 27872
rect -22147 27808 -22127 27872
rect -28426 27792 -22127 27808
rect -28426 27728 -22211 27792
rect -22147 27728 -22127 27792
rect -28426 27712 -22127 27728
rect -28426 27648 -22211 27712
rect -22147 27648 -22127 27712
rect -28426 27632 -22127 27648
rect -28426 27568 -22211 27632
rect -22147 27568 -22127 27632
rect -28426 27552 -22127 27568
rect -28426 27488 -22211 27552
rect -22147 27488 -22127 27552
rect -28426 27472 -22127 27488
rect -28426 27408 -22211 27472
rect -22147 27408 -22127 27472
rect -28426 27392 -22127 27408
rect -28426 27328 -22211 27392
rect -22147 27328 -22127 27392
rect -28426 27312 -22127 27328
rect -28426 27248 -22211 27312
rect -22147 27248 -22127 27312
rect -28426 27232 -22127 27248
rect -28426 27168 -22211 27232
rect -22147 27168 -22127 27232
rect -28426 27152 -22127 27168
rect -28426 27088 -22211 27152
rect -22147 27088 -22127 27152
rect -28426 27072 -22127 27088
rect -28426 27008 -22211 27072
rect -22147 27008 -22127 27072
rect -28426 26992 -22127 27008
rect -28426 26928 -22211 26992
rect -22147 26928 -22127 26992
rect -28426 26912 -22127 26928
rect -28426 26848 -22211 26912
rect -22147 26848 -22127 26912
rect -28426 26832 -22127 26848
rect -28426 26768 -22211 26832
rect -22147 26768 -22127 26832
rect -28426 26752 -22127 26768
rect -28426 26688 -22211 26752
rect -22147 26688 -22127 26752
rect -28426 26672 -22127 26688
rect -28426 26608 -22211 26672
rect -22147 26608 -22127 26672
rect -28426 26592 -22127 26608
rect -28426 26528 -22211 26592
rect -22147 26528 -22127 26592
rect -28426 26512 -22127 26528
rect -28426 26448 -22211 26512
rect -22147 26448 -22127 26512
rect -28426 26432 -22127 26448
rect -28426 26368 -22211 26432
rect -22147 26368 -22127 26432
rect -28426 26352 -22127 26368
rect -28426 26288 -22211 26352
rect -22147 26288 -22127 26352
rect -28426 26272 -22127 26288
rect -28426 26208 -22211 26272
rect -22147 26208 -22127 26272
rect -28426 26192 -22127 26208
rect -28426 26128 -22211 26192
rect -22147 26128 -22127 26192
rect -28426 26112 -22127 26128
rect -28426 26048 -22211 26112
rect -22147 26048 -22127 26112
rect -28426 26032 -22127 26048
rect -28426 25968 -22211 26032
rect -22147 25968 -22127 26032
rect -28426 25952 -22127 25968
rect -28426 25888 -22211 25952
rect -22147 25888 -22127 25952
rect -28426 25872 -22127 25888
rect -28426 25808 -22211 25872
rect -22147 25808 -22127 25872
rect -28426 25792 -22127 25808
rect -28426 25728 -22211 25792
rect -22147 25728 -22127 25792
rect -28426 25712 -22127 25728
rect -28426 25648 -22211 25712
rect -22147 25648 -22127 25712
rect -28426 25632 -22127 25648
rect -28426 25568 -22211 25632
rect -22147 25568 -22127 25632
rect -28426 25552 -22127 25568
rect -28426 25488 -22211 25552
rect -22147 25488 -22127 25552
rect -28426 25472 -22127 25488
rect -28426 25408 -22211 25472
rect -22147 25408 -22127 25472
rect -28426 25392 -22127 25408
rect -28426 25328 -22211 25392
rect -22147 25328 -22127 25392
rect -28426 25312 -22127 25328
rect -28426 25248 -22211 25312
rect -22147 25248 -22127 25312
rect -28426 25232 -22127 25248
rect -28426 25168 -22211 25232
rect -22147 25168 -22127 25232
rect -28426 25152 -22127 25168
rect -28426 25088 -22211 25152
rect -22147 25088 -22127 25152
rect -28426 25072 -22127 25088
rect -28426 25008 -22211 25072
rect -22147 25008 -22127 25072
rect -28426 24992 -22127 25008
rect -28426 24928 -22211 24992
rect -22147 24928 -22127 24992
rect -28426 24912 -22127 24928
rect -28426 24848 -22211 24912
rect -22147 24848 -22127 24912
rect -28426 24832 -22127 24848
rect -28426 24768 -22211 24832
rect -22147 24768 -22127 24832
rect -28426 24752 -22127 24768
rect -28426 24688 -22211 24752
rect -22147 24688 -22127 24752
rect -28426 24672 -22127 24688
rect -28426 24608 -22211 24672
rect -22147 24608 -22127 24672
rect -28426 24592 -22127 24608
rect -28426 24528 -22211 24592
rect -22147 24528 -22127 24592
rect -28426 24512 -22127 24528
rect -28426 24448 -22211 24512
rect -22147 24448 -22127 24512
rect -28426 24432 -22127 24448
rect -28426 24368 -22211 24432
rect -22147 24368 -22127 24432
rect -28426 24352 -22127 24368
rect -28426 24288 -22211 24352
rect -22147 24288 -22127 24352
rect -28426 24272 -22127 24288
rect -28426 24208 -22211 24272
rect -22147 24208 -22127 24272
rect -28426 24192 -22127 24208
rect -28426 24128 -22211 24192
rect -22147 24128 -22127 24192
rect -28426 24112 -22127 24128
rect -28426 24048 -22211 24112
rect -22147 24048 -22127 24112
rect -28426 24032 -22127 24048
rect -28426 23968 -22211 24032
rect -22147 23968 -22127 24032
rect -28426 23952 -22127 23968
rect -28426 23888 -22211 23952
rect -22147 23888 -22127 23952
rect -28426 23872 -22127 23888
rect -28426 23808 -22211 23872
rect -22147 23808 -22127 23872
rect -28426 23792 -22127 23808
rect -28426 23728 -22211 23792
rect -22147 23728 -22127 23792
rect -28426 23712 -22127 23728
rect -28426 23648 -22211 23712
rect -22147 23648 -22127 23712
rect -28426 23632 -22127 23648
rect -28426 23568 -22211 23632
rect -22147 23568 -22127 23632
rect -28426 23552 -22127 23568
rect -28426 23488 -22211 23552
rect -22147 23488 -22127 23552
rect -28426 23472 -22127 23488
rect -28426 23408 -22211 23472
rect -22147 23408 -22127 23472
rect -28426 23392 -22127 23408
rect -28426 23328 -22211 23392
rect -22147 23328 -22127 23392
rect -28426 23312 -22127 23328
rect -28426 23248 -22211 23312
rect -22147 23248 -22127 23312
rect -28426 23232 -22127 23248
rect -28426 23168 -22211 23232
rect -22147 23168 -22127 23232
rect -28426 23152 -22127 23168
rect -28426 23088 -22211 23152
rect -22147 23088 -22127 23152
rect -28426 23072 -22127 23088
rect -28426 23008 -22211 23072
rect -22147 23008 -22127 23072
rect -28426 22992 -22127 23008
rect -28426 22928 -22211 22992
rect -22147 22928 -22127 22992
rect -28426 22912 -22127 22928
rect -28426 22848 -22211 22912
rect -22147 22848 -22127 22912
rect -28426 22832 -22127 22848
rect -28426 22768 -22211 22832
rect -22147 22768 -22127 22832
rect -28426 22752 -22127 22768
rect -28426 22688 -22211 22752
rect -22147 22688 -22127 22752
rect -28426 22672 -22127 22688
rect -28426 22608 -22211 22672
rect -22147 22608 -22127 22672
rect -28426 22592 -22127 22608
rect -28426 22528 -22211 22592
rect -22147 22528 -22127 22592
rect -28426 22512 -22127 22528
rect -28426 22448 -22211 22512
rect -22147 22448 -22127 22512
rect -28426 22432 -22127 22448
rect -28426 22368 -22211 22432
rect -22147 22368 -22127 22432
rect -28426 22352 -22127 22368
rect -28426 22288 -22211 22352
rect -22147 22288 -22127 22352
rect -28426 22272 -22127 22288
rect -28426 22208 -22211 22272
rect -22147 22208 -22127 22272
rect -28426 22192 -22127 22208
rect -28426 22128 -22211 22192
rect -22147 22128 -22127 22192
rect -28426 22100 -22127 22128
rect -22107 28272 -15808 28300
rect -22107 28208 -15892 28272
rect -15828 28208 -15808 28272
rect -22107 28192 -15808 28208
rect -22107 28128 -15892 28192
rect -15828 28128 -15808 28192
rect -22107 28112 -15808 28128
rect -22107 28048 -15892 28112
rect -15828 28048 -15808 28112
rect -22107 28032 -15808 28048
rect -22107 27968 -15892 28032
rect -15828 27968 -15808 28032
rect -22107 27952 -15808 27968
rect -22107 27888 -15892 27952
rect -15828 27888 -15808 27952
rect -22107 27872 -15808 27888
rect -22107 27808 -15892 27872
rect -15828 27808 -15808 27872
rect -22107 27792 -15808 27808
rect -22107 27728 -15892 27792
rect -15828 27728 -15808 27792
rect -22107 27712 -15808 27728
rect -22107 27648 -15892 27712
rect -15828 27648 -15808 27712
rect -22107 27632 -15808 27648
rect -22107 27568 -15892 27632
rect -15828 27568 -15808 27632
rect -22107 27552 -15808 27568
rect -22107 27488 -15892 27552
rect -15828 27488 -15808 27552
rect -22107 27472 -15808 27488
rect -22107 27408 -15892 27472
rect -15828 27408 -15808 27472
rect -22107 27392 -15808 27408
rect -22107 27328 -15892 27392
rect -15828 27328 -15808 27392
rect -22107 27312 -15808 27328
rect -22107 27248 -15892 27312
rect -15828 27248 -15808 27312
rect -22107 27232 -15808 27248
rect -22107 27168 -15892 27232
rect -15828 27168 -15808 27232
rect -22107 27152 -15808 27168
rect -22107 27088 -15892 27152
rect -15828 27088 -15808 27152
rect -22107 27072 -15808 27088
rect -22107 27008 -15892 27072
rect -15828 27008 -15808 27072
rect -22107 26992 -15808 27008
rect -22107 26928 -15892 26992
rect -15828 26928 -15808 26992
rect -22107 26912 -15808 26928
rect -22107 26848 -15892 26912
rect -15828 26848 -15808 26912
rect -22107 26832 -15808 26848
rect -22107 26768 -15892 26832
rect -15828 26768 -15808 26832
rect -22107 26752 -15808 26768
rect -22107 26688 -15892 26752
rect -15828 26688 -15808 26752
rect -22107 26672 -15808 26688
rect -22107 26608 -15892 26672
rect -15828 26608 -15808 26672
rect -22107 26592 -15808 26608
rect -22107 26528 -15892 26592
rect -15828 26528 -15808 26592
rect -22107 26512 -15808 26528
rect -22107 26448 -15892 26512
rect -15828 26448 -15808 26512
rect -22107 26432 -15808 26448
rect -22107 26368 -15892 26432
rect -15828 26368 -15808 26432
rect -22107 26352 -15808 26368
rect -22107 26288 -15892 26352
rect -15828 26288 -15808 26352
rect -22107 26272 -15808 26288
rect -22107 26208 -15892 26272
rect -15828 26208 -15808 26272
rect -22107 26192 -15808 26208
rect -22107 26128 -15892 26192
rect -15828 26128 -15808 26192
rect -22107 26112 -15808 26128
rect -22107 26048 -15892 26112
rect -15828 26048 -15808 26112
rect -22107 26032 -15808 26048
rect -22107 25968 -15892 26032
rect -15828 25968 -15808 26032
rect -22107 25952 -15808 25968
rect -22107 25888 -15892 25952
rect -15828 25888 -15808 25952
rect -22107 25872 -15808 25888
rect -22107 25808 -15892 25872
rect -15828 25808 -15808 25872
rect -22107 25792 -15808 25808
rect -22107 25728 -15892 25792
rect -15828 25728 -15808 25792
rect -22107 25712 -15808 25728
rect -22107 25648 -15892 25712
rect -15828 25648 -15808 25712
rect -22107 25632 -15808 25648
rect -22107 25568 -15892 25632
rect -15828 25568 -15808 25632
rect -22107 25552 -15808 25568
rect -22107 25488 -15892 25552
rect -15828 25488 -15808 25552
rect -22107 25472 -15808 25488
rect -22107 25408 -15892 25472
rect -15828 25408 -15808 25472
rect -22107 25392 -15808 25408
rect -22107 25328 -15892 25392
rect -15828 25328 -15808 25392
rect -22107 25312 -15808 25328
rect -22107 25248 -15892 25312
rect -15828 25248 -15808 25312
rect -22107 25232 -15808 25248
rect -22107 25168 -15892 25232
rect -15828 25168 -15808 25232
rect -22107 25152 -15808 25168
rect -22107 25088 -15892 25152
rect -15828 25088 -15808 25152
rect -22107 25072 -15808 25088
rect -22107 25008 -15892 25072
rect -15828 25008 -15808 25072
rect -22107 24992 -15808 25008
rect -22107 24928 -15892 24992
rect -15828 24928 -15808 24992
rect -22107 24912 -15808 24928
rect -22107 24848 -15892 24912
rect -15828 24848 -15808 24912
rect -22107 24832 -15808 24848
rect -22107 24768 -15892 24832
rect -15828 24768 -15808 24832
rect -22107 24752 -15808 24768
rect -22107 24688 -15892 24752
rect -15828 24688 -15808 24752
rect -22107 24672 -15808 24688
rect -22107 24608 -15892 24672
rect -15828 24608 -15808 24672
rect -22107 24592 -15808 24608
rect -22107 24528 -15892 24592
rect -15828 24528 -15808 24592
rect -22107 24512 -15808 24528
rect -22107 24448 -15892 24512
rect -15828 24448 -15808 24512
rect -22107 24432 -15808 24448
rect -22107 24368 -15892 24432
rect -15828 24368 -15808 24432
rect -22107 24352 -15808 24368
rect -22107 24288 -15892 24352
rect -15828 24288 -15808 24352
rect -22107 24272 -15808 24288
rect -22107 24208 -15892 24272
rect -15828 24208 -15808 24272
rect -22107 24192 -15808 24208
rect -22107 24128 -15892 24192
rect -15828 24128 -15808 24192
rect -22107 24112 -15808 24128
rect -22107 24048 -15892 24112
rect -15828 24048 -15808 24112
rect -22107 24032 -15808 24048
rect -22107 23968 -15892 24032
rect -15828 23968 -15808 24032
rect -22107 23952 -15808 23968
rect -22107 23888 -15892 23952
rect -15828 23888 -15808 23952
rect -22107 23872 -15808 23888
rect -22107 23808 -15892 23872
rect -15828 23808 -15808 23872
rect -22107 23792 -15808 23808
rect -22107 23728 -15892 23792
rect -15828 23728 -15808 23792
rect -22107 23712 -15808 23728
rect -22107 23648 -15892 23712
rect -15828 23648 -15808 23712
rect -22107 23632 -15808 23648
rect -22107 23568 -15892 23632
rect -15828 23568 -15808 23632
rect -22107 23552 -15808 23568
rect -22107 23488 -15892 23552
rect -15828 23488 -15808 23552
rect -22107 23472 -15808 23488
rect -22107 23408 -15892 23472
rect -15828 23408 -15808 23472
rect -22107 23392 -15808 23408
rect -22107 23328 -15892 23392
rect -15828 23328 -15808 23392
rect -22107 23312 -15808 23328
rect -22107 23248 -15892 23312
rect -15828 23248 -15808 23312
rect -22107 23232 -15808 23248
rect -22107 23168 -15892 23232
rect -15828 23168 -15808 23232
rect -22107 23152 -15808 23168
rect -22107 23088 -15892 23152
rect -15828 23088 -15808 23152
rect -22107 23072 -15808 23088
rect -22107 23008 -15892 23072
rect -15828 23008 -15808 23072
rect -22107 22992 -15808 23008
rect -22107 22928 -15892 22992
rect -15828 22928 -15808 22992
rect -22107 22912 -15808 22928
rect -22107 22848 -15892 22912
rect -15828 22848 -15808 22912
rect -22107 22832 -15808 22848
rect -22107 22768 -15892 22832
rect -15828 22768 -15808 22832
rect -22107 22752 -15808 22768
rect -22107 22688 -15892 22752
rect -15828 22688 -15808 22752
rect -22107 22672 -15808 22688
rect -22107 22608 -15892 22672
rect -15828 22608 -15808 22672
rect -22107 22592 -15808 22608
rect -22107 22528 -15892 22592
rect -15828 22528 -15808 22592
rect -22107 22512 -15808 22528
rect -22107 22448 -15892 22512
rect -15828 22448 -15808 22512
rect -22107 22432 -15808 22448
rect -22107 22368 -15892 22432
rect -15828 22368 -15808 22432
rect -22107 22352 -15808 22368
rect -22107 22288 -15892 22352
rect -15828 22288 -15808 22352
rect -22107 22272 -15808 22288
rect -22107 22208 -15892 22272
rect -15828 22208 -15808 22272
rect -22107 22192 -15808 22208
rect -22107 22128 -15892 22192
rect -15828 22128 -15808 22192
rect -22107 22100 -15808 22128
rect -15788 28272 -9489 28300
rect -15788 28208 -9573 28272
rect -9509 28208 -9489 28272
rect -15788 28192 -9489 28208
rect -15788 28128 -9573 28192
rect -9509 28128 -9489 28192
rect -15788 28112 -9489 28128
rect -15788 28048 -9573 28112
rect -9509 28048 -9489 28112
rect -15788 28032 -9489 28048
rect -15788 27968 -9573 28032
rect -9509 27968 -9489 28032
rect -15788 27952 -9489 27968
rect -15788 27888 -9573 27952
rect -9509 27888 -9489 27952
rect -15788 27872 -9489 27888
rect -15788 27808 -9573 27872
rect -9509 27808 -9489 27872
rect -15788 27792 -9489 27808
rect -15788 27728 -9573 27792
rect -9509 27728 -9489 27792
rect -15788 27712 -9489 27728
rect -15788 27648 -9573 27712
rect -9509 27648 -9489 27712
rect -15788 27632 -9489 27648
rect -15788 27568 -9573 27632
rect -9509 27568 -9489 27632
rect -15788 27552 -9489 27568
rect -15788 27488 -9573 27552
rect -9509 27488 -9489 27552
rect -15788 27472 -9489 27488
rect -15788 27408 -9573 27472
rect -9509 27408 -9489 27472
rect -15788 27392 -9489 27408
rect -15788 27328 -9573 27392
rect -9509 27328 -9489 27392
rect -15788 27312 -9489 27328
rect -15788 27248 -9573 27312
rect -9509 27248 -9489 27312
rect -15788 27232 -9489 27248
rect -15788 27168 -9573 27232
rect -9509 27168 -9489 27232
rect -15788 27152 -9489 27168
rect -15788 27088 -9573 27152
rect -9509 27088 -9489 27152
rect -15788 27072 -9489 27088
rect -15788 27008 -9573 27072
rect -9509 27008 -9489 27072
rect -15788 26992 -9489 27008
rect -15788 26928 -9573 26992
rect -9509 26928 -9489 26992
rect -15788 26912 -9489 26928
rect -15788 26848 -9573 26912
rect -9509 26848 -9489 26912
rect -15788 26832 -9489 26848
rect -15788 26768 -9573 26832
rect -9509 26768 -9489 26832
rect -15788 26752 -9489 26768
rect -15788 26688 -9573 26752
rect -9509 26688 -9489 26752
rect -15788 26672 -9489 26688
rect -15788 26608 -9573 26672
rect -9509 26608 -9489 26672
rect -15788 26592 -9489 26608
rect -15788 26528 -9573 26592
rect -9509 26528 -9489 26592
rect -15788 26512 -9489 26528
rect -15788 26448 -9573 26512
rect -9509 26448 -9489 26512
rect -15788 26432 -9489 26448
rect -15788 26368 -9573 26432
rect -9509 26368 -9489 26432
rect -15788 26352 -9489 26368
rect -15788 26288 -9573 26352
rect -9509 26288 -9489 26352
rect -15788 26272 -9489 26288
rect -15788 26208 -9573 26272
rect -9509 26208 -9489 26272
rect -15788 26192 -9489 26208
rect -15788 26128 -9573 26192
rect -9509 26128 -9489 26192
rect -15788 26112 -9489 26128
rect -15788 26048 -9573 26112
rect -9509 26048 -9489 26112
rect -15788 26032 -9489 26048
rect -15788 25968 -9573 26032
rect -9509 25968 -9489 26032
rect -15788 25952 -9489 25968
rect -15788 25888 -9573 25952
rect -9509 25888 -9489 25952
rect -15788 25872 -9489 25888
rect -15788 25808 -9573 25872
rect -9509 25808 -9489 25872
rect -15788 25792 -9489 25808
rect -15788 25728 -9573 25792
rect -9509 25728 -9489 25792
rect -15788 25712 -9489 25728
rect -15788 25648 -9573 25712
rect -9509 25648 -9489 25712
rect -15788 25632 -9489 25648
rect -15788 25568 -9573 25632
rect -9509 25568 -9489 25632
rect -15788 25552 -9489 25568
rect -15788 25488 -9573 25552
rect -9509 25488 -9489 25552
rect -15788 25472 -9489 25488
rect -15788 25408 -9573 25472
rect -9509 25408 -9489 25472
rect -15788 25392 -9489 25408
rect -15788 25328 -9573 25392
rect -9509 25328 -9489 25392
rect -15788 25312 -9489 25328
rect -15788 25248 -9573 25312
rect -9509 25248 -9489 25312
rect -15788 25232 -9489 25248
rect -15788 25168 -9573 25232
rect -9509 25168 -9489 25232
rect -15788 25152 -9489 25168
rect -15788 25088 -9573 25152
rect -9509 25088 -9489 25152
rect -15788 25072 -9489 25088
rect -15788 25008 -9573 25072
rect -9509 25008 -9489 25072
rect -15788 24992 -9489 25008
rect -15788 24928 -9573 24992
rect -9509 24928 -9489 24992
rect -15788 24912 -9489 24928
rect -15788 24848 -9573 24912
rect -9509 24848 -9489 24912
rect -15788 24832 -9489 24848
rect -15788 24768 -9573 24832
rect -9509 24768 -9489 24832
rect -15788 24752 -9489 24768
rect -15788 24688 -9573 24752
rect -9509 24688 -9489 24752
rect -15788 24672 -9489 24688
rect -15788 24608 -9573 24672
rect -9509 24608 -9489 24672
rect -15788 24592 -9489 24608
rect -15788 24528 -9573 24592
rect -9509 24528 -9489 24592
rect -15788 24512 -9489 24528
rect -15788 24448 -9573 24512
rect -9509 24448 -9489 24512
rect -15788 24432 -9489 24448
rect -15788 24368 -9573 24432
rect -9509 24368 -9489 24432
rect -15788 24352 -9489 24368
rect -15788 24288 -9573 24352
rect -9509 24288 -9489 24352
rect -15788 24272 -9489 24288
rect -15788 24208 -9573 24272
rect -9509 24208 -9489 24272
rect -15788 24192 -9489 24208
rect -15788 24128 -9573 24192
rect -9509 24128 -9489 24192
rect -15788 24112 -9489 24128
rect -15788 24048 -9573 24112
rect -9509 24048 -9489 24112
rect -15788 24032 -9489 24048
rect -15788 23968 -9573 24032
rect -9509 23968 -9489 24032
rect -15788 23952 -9489 23968
rect -15788 23888 -9573 23952
rect -9509 23888 -9489 23952
rect -15788 23872 -9489 23888
rect -15788 23808 -9573 23872
rect -9509 23808 -9489 23872
rect -15788 23792 -9489 23808
rect -15788 23728 -9573 23792
rect -9509 23728 -9489 23792
rect -15788 23712 -9489 23728
rect -15788 23648 -9573 23712
rect -9509 23648 -9489 23712
rect -15788 23632 -9489 23648
rect -15788 23568 -9573 23632
rect -9509 23568 -9489 23632
rect -15788 23552 -9489 23568
rect -15788 23488 -9573 23552
rect -9509 23488 -9489 23552
rect -15788 23472 -9489 23488
rect -15788 23408 -9573 23472
rect -9509 23408 -9489 23472
rect -15788 23392 -9489 23408
rect -15788 23328 -9573 23392
rect -9509 23328 -9489 23392
rect -15788 23312 -9489 23328
rect -15788 23248 -9573 23312
rect -9509 23248 -9489 23312
rect -15788 23232 -9489 23248
rect -15788 23168 -9573 23232
rect -9509 23168 -9489 23232
rect -15788 23152 -9489 23168
rect -15788 23088 -9573 23152
rect -9509 23088 -9489 23152
rect -15788 23072 -9489 23088
rect -15788 23008 -9573 23072
rect -9509 23008 -9489 23072
rect -15788 22992 -9489 23008
rect -15788 22928 -9573 22992
rect -9509 22928 -9489 22992
rect -15788 22912 -9489 22928
rect -15788 22848 -9573 22912
rect -9509 22848 -9489 22912
rect -15788 22832 -9489 22848
rect -15788 22768 -9573 22832
rect -9509 22768 -9489 22832
rect -15788 22752 -9489 22768
rect -15788 22688 -9573 22752
rect -9509 22688 -9489 22752
rect -15788 22672 -9489 22688
rect -15788 22608 -9573 22672
rect -9509 22608 -9489 22672
rect -15788 22592 -9489 22608
rect -15788 22528 -9573 22592
rect -9509 22528 -9489 22592
rect -15788 22512 -9489 22528
rect -15788 22448 -9573 22512
rect -9509 22448 -9489 22512
rect -15788 22432 -9489 22448
rect -15788 22368 -9573 22432
rect -9509 22368 -9489 22432
rect -15788 22352 -9489 22368
rect -15788 22288 -9573 22352
rect -9509 22288 -9489 22352
rect -15788 22272 -9489 22288
rect -15788 22208 -9573 22272
rect -9509 22208 -9489 22272
rect -15788 22192 -9489 22208
rect -15788 22128 -9573 22192
rect -9509 22128 -9489 22192
rect -15788 22100 -9489 22128
rect -9469 28272 -3170 28300
rect -9469 28208 -3254 28272
rect -3190 28208 -3170 28272
rect -9469 28192 -3170 28208
rect -9469 28128 -3254 28192
rect -3190 28128 -3170 28192
rect -9469 28112 -3170 28128
rect -9469 28048 -3254 28112
rect -3190 28048 -3170 28112
rect -9469 28032 -3170 28048
rect -9469 27968 -3254 28032
rect -3190 27968 -3170 28032
rect -9469 27952 -3170 27968
rect -9469 27888 -3254 27952
rect -3190 27888 -3170 27952
rect -9469 27872 -3170 27888
rect -9469 27808 -3254 27872
rect -3190 27808 -3170 27872
rect -9469 27792 -3170 27808
rect -9469 27728 -3254 27792
rect -3190 27728 -3170 27792
rect -9469 27712 -3170 27728
rect -9469 27648 -3254 27712
rect -3190 27648 -3170 27712
rect -9469 27632 -3170 27648
rect -9469 27568 -3254 27632
rect -3190 27568 -3170 27632
rect -9469 27552 -3170 27568
rect -9469 27488 -3254 27552
rect -3190 27488 -3170 27552
rect -9469 27472 -3170 27488
rect -9469 27408 -3254 27472
rect -3190 27408 -3170 27472
rect -9469 27392 -3170 27408
rect -9469 27328 -3254 27392
rect -3190 27328 -3170 27392
rect -9469 27312 -3170 27328
rect -9469 27248 -3254 27312
rect -3190 27248 -3170 27312
rect -9469 27232 -3170 27248
rect -9469 27168 -3254 27232
rect -3190 27168 -3170 27232
rect -9469 27152 -3170 27168
rect -9469 27088 -3254 27152
rect -3190 27088 -3170 27152
rect -9469 27072 -3170 27088
rect -9469 27008 -3254 27072
rect -3190 27008 -3170 27072
rect -9469 26992 -3170 27008
rect -9469 26928 -3254 26992
rect -3190 26928 -3170 26992
rect -9469 26912 -3170 26928
rect -9469 26848 -3254 26912
rect -3190 26848 -3170 26912
rect -9469 26832 -3170 26848
rect -9469 26768 -3254 26832
rect -3190 26768 -3170 26832
rect -9469 26752 -3170 26768
rect -9469 26688 -3254 26752
rect -3190 26688 -3170 26752
rect -9469 26672 -3170 26688
rect -9469 26608 -3254 26672
rect -3190 26608 -3170 26672
rect -9469 26592 -3170 26608
rect -9469 26528 -3254 26592
rect -3190 26528 -3170 26592
rect -9469 26512 -3170 26528
rect -9469 26448 -3254 26512
rect -3190 26448 -3170 26512
rect -9469 26432 -3170 26448
rect -9469 26368 -3254 26432
rect -3190 26368 -3170 26432
rect -9469 26352 -3170 26368
rect -9469 26288 -3254 26352
rect -3190 26288 -3170 26352
rect -9469 26272 -3170 26288
rect -9469 26208 -3254 26272
rect -3190 26208 -3170 26272
rect -9469 26192 -3170 26208
rect -9469 26128 -3254 26192
rect -3190 26128 -3170 26192
rect -9469 26112 -3170 26128
rect -9469 26048 -3254 26112
rect -3190 26048 -3170 26112
rect -9469 26032 -3170 26048
rect -9469 25968 -3254 26032
rect -3190 25968 -3170 26032
rect -9469 25952 -3170 25968
rect -9469 25888 -3254 25952
rect -3190 25888 -3170 25952
rect -9469 25872 -3170 25888
rect -9469 25808 -3254 25872
rect -3190 25808 -3170 25872
rect -9469 25792 -3170 25808
rect -9469 25728 -3254 25792
rect -3190 25728 -3170 25792
rect -9469 25712 -3170 25728
rect -9469 25648 -3254 25712
rect -3190 25648 -3170 25712
rect -9469 25632 -3170 25648
rect -9469 25568 -3254 25632
rect -3190 25568 -3170 25632
rect -9469 25552 -3170 25568
rect -9469 25488 -3254 25552
rect -3190 25488 -3170 25552
rect -9469 25472 -3170 25488
rect -9469 25408 -3254 25472
rect -3190 25408 -3170 25472
rect -9469 25392 -3170 25408
rect -9469 25328 -3254 25392
rect -3190 25328 -3170 25392
rect -9469 25312 -3170 25328
rect -9469 25248 -3254 25312
rect -3190 25248 -3170 25312
rect -9469 25232 -3170 25248
rect -9469 25168 -3254 25232
rect -3190 25168 -3170 25232
rect -9469 25152 -3170 25168
rect -9469 25088 -3254 25152
rect -3190 25088 -3170 25152
rect -9469 25072 -3170 25088
rect -9469 25008 -3254 25072
rect -3190 25008 -3170 25072
rect -9469 24992 -3170 25008
rect -9469 24928 -3254 24992
rect -3190 24928 -3170 24992
rect -9469 24912 -3170 24928
rect -9469 24848 -3254 24912
rect -3190 24848 -3170 24912
rect -9469 24832 -3170 24848
rect -9469 24768 -3254 24832
rect -3190 24768 -3170 24832
rect -9469 24752 -3170 24768
rect -9469 24688 -3254 24752
rect -3190 24688 -3170 24752
rect -9469 24672 -3170 24688
rect -9469 24608 -3254 24672
rect -3190 24608 -3170 24672
rect -9469 24592 -3170 24608
rect -9469 24528 -3254 24592
rect -3190 24528 -3170 24592
rect -9469 24512 -3170 24528
rect -9469 24448 -3254 24512
rect -3190 24448 -3170 24512
rect -9469 24432 -3170 24448
rect -9469 24368 -3254 24432
rect -3190 24368 -3170 24432
rect -9469 24352 -3170 24368
rect -9469 24288 -3254 24352
rect -3190 24288 -3170 24352
rect -9469 24272 -3170 24288
rect -9469 24208 -3254 24272
rect -3190 24208 -3170 24272
rect -9469 24192 -3170 24208
rect -9469 24128 -3254 24192
rect -3190 24128 -3170 24192
rect -9469 24112 -3170 24128
rect -9469 24048 -3254 24112
rect -3190 24048 -3170 24112
rect -9469 24032 -3170 24048
rect -9469 23968 -3254 24032
rect -3190 23968 -3170 24032
rect -9469 23952 -3170 23968
rect -9469 23888 -3254 23952
rect -3190 23888 -3170 23952
rect -9469 23872 -3170 23888
rect -9469 23808 -3254 23872
rect -3190 23808 -3170 23872
rect -9469 23792 -3170 23808
rect -9469 23728 -3254 23792
rect -3190 23728 -3170 23792
rect -9469 23712 -3170 23728
rect -9469 23648 -3254 23712
rect -3190 23648 -3170 23712
rect -9469 23632 -3170 23648
rect -9469 23568 -3254 23632
rect -3190 23568 -3170 23632
rect -9469 23552 -3170 23568
rect -9469 23488 -3254 23552
rect -3190 23488 -3170 23552
rect -9469 23472 -3170 23488
rect -9469 23408 -3254 23472
rect -3190 23408 -3170 23472
rect -9469 23392 -3170 23408
rect -9469 23328 -3254 23392
rect -3190 23328 -3170 23392
rect -9469 23312 -3170 23328
rect -9469 23248 -3254 23312
rect -3190 23248 -3170 23312
rect -9469 23232 -3170 23248
rect -9469 23168 -3254 23232
rect -3190 23168 -3170 23232
rect -9469 23152 -3170 23168
rect -9469 23088 -3254 23152
rect -3190 23088 -3170 23152
rect -9469 23072 -3170 23088
rect -9469 23008 -3254 23072
rect -3190 23008 -3170 23072
rect -9469 22992 -3170 23008
rect -9469 22928 -3254 22992
rect -3190 22928 -3170 22992
rect -9469 22912 -3170 22928
rect -9469 22848 -3254 22912
rect -3190 22848 -3170 22912
rect -9469 22832 -3170 22848
rect -9469 22768 -3254 22832
rect -3190 22768 -3170 22832
rect -9469 22752 -3170 22768
rect -9469 22688 -3254 22752
rect -3190 22688 -3170 22752
rect -9469 22672 -3170 22688
rect -9469 22608 -3254 22672
rect -3190 22608 -3170 22672
rect -9469 22592 -3170 22608
rect -9469 22528 -3254 22592
rect -3190 22528 -3170 22592
rect -9469 22512 -3170 22528
rect -9469 22448 -3254 22512
rect -3190 22448 -3170 22512
rect -9469 22432 -3170 22448
rect -9469 22368 -3254 22432
rect -3190 22368 -3170 22432
rect -9469 22352 -3170 22368
rect -9469 22288 -3254 22352
rect -3190 22288 -3170 22352
rect -9469 22272 -3170 22288
rect -9469 22208 -3254 22272
rect -3190 22208 -3170 22272
rect -9469 22192 -3170 22208
rect -9469 22128 -3254 22192
rect -3190 22128 -3170 22192
rect -9469 22100 -3170 22128
rect -3150 28272 3149 28300
rect -3150 28208 3065 28272
rect 3129 28208 3149 28272
rect -3150 28192 3149 28208
rect -3150 28128 3065 28192
rect 3129 28128 3149 28192
rect -3150 28112 3149 28128
rect -3150 28048 3065 28112
rect 3129 28048 3149 28112
rect -3150 28032 3149 28048
rect -3150 27968 3065 28032
rect 3129 27968 3149 28032
rect -3150 27952 3149 27968
rect -3150 27888 3065 27952
rect 3129 27888 3149 27952
rect -3150 27872 3149 27888
rect -3150 27808 3065 27872
rect 3129 27808 3149 27872
rect -3150 27792 3149 27808
rect -3150 27728 3065 27792
rect 3129 27728 3149 27792
rect -3150 27712 3149 27728
rect -3150 27648 3065 27712
rect 3129 27648 3149 27712
rect -3150 27632 3149 27648
rect -3150 27568 3065 27632
rect 3129 27568 3149 27632
rect -3150 27552 3149 27568
rect -3150 27488 3065 27552
rect 3129 27488 3149 27552
rect -3150 27472 3149 27488
rect -3150 27408 3065 27472
rect 3129 27408 3149 27472
rect -3150 27392 3149 27408
rect -3150 27328 3065 27392
rect 3129 27328 3149 27392
rect -3150 27312 3149 27328
rect -3150 27248 3065 27312
rect 3129 27248 3149 27312
rect -3150 27232 3149 27248
rect -3150 27168 3065 27232
rect 3129 27168 3149 27232
rect -3150 27152 3149 27168
rect -3150 27088 3065 27152
rect 3129 27088 3149 27152
rect -3150 27072 3149 27088
rect -3150 27008 3065 27072
rect 3129 27008 3149 27072
rect -3150 26992 3149 27008
rect -3150 26928 3065 26992
rect 3129 26928 3149 26992
rect -3150 26912 3149 26928
rect -3150 26848 3065 26912
rect 3129 26848 3149 26912
rect -3150 26832 3149 26848
rect -3150 26768 3065 26832
rect 3129 26768 3149 26832
rect -3150 26752 3149 26768
rect -3150 26688 3065 26752
rect 3129 26688 3149 26752
rect -3150 26672 3149 26688
rect -3150 26608 3065 26672
rect 3129 26608 3149 26672
rect -3150 26592 3149 26608
rect -3150 26528 3065 26592
rect 3129 26528 3149 26592
rect -3150 26512 3149 26528
rect -3150 26448 3065 26512
rect 3129 26448 3149 26512
rect -3150 26432 3149 26448
rect -3150 26368 3065 26432
rect 3129 26368 3149 26432
rect -3150 26352 3149 26368
rect -3150 26288 3065 26352
rect 3129 26288 3149 26352
rect -3150 26272 3149 26288
rect -3150 26208 3065 26272
rect 3129 26208 3149 26272
rect -3150 26192 3149 26208
rect -3150 26128 3065 26192
rect 3129 26128 3149 26192
rect -3150 26112 3149 26128
rect -3150 26048 3065 26112
rect 3129 26048 3149 26112
rect -3150 26032 3149 26048
rect -3150 25968 3065 26032
rect 3129 25968 3149 26032
rect -3150 25952 3149 25968
rect -3150 25888 3065 25952
rect 3129 25888 3149 25952
rect -3150 25872 3149 25888
rect -3150 25808 3065 25872
rect 3129 25808 3149 25872
rect -3150 25792 3149 25808
rect -3150 25728 3065 25792
rect 3129 25728 3149 25792
rect -3150 25712 3149 25728
rect -3150 25648 3065 25712
rect 3129 25648 3149 25712
rect -3150 25632 3149 25648
rect -3150 25568 3065 25632
rect 3129 25568 3149 25632
rect -3150 25552 3149 25568
rect -3150 25488 3065 25552
rect 3129 25488 3149 25552
rect -3150 25472 3149 25488
rect -3150 25408 3065 25472
rect 3129 25408 3149 25472
rect -3150 25392 3149 25408
rect -3150 25328 3065 25392
rect 3129 25328 3149 25392
rect -3150 25312 3149 25328
rect -3150 25248 3065 25312
rect 3129 25248 3149 25312
rect -3150 25232 3149 25248
rect -3150 25168 3065 25232
rect 3129 25168 3149 25232
rect -3150 25152 3149 25168
rect -3150 25088 3065 25152
rect 3129 25088 3149 25152
rect -3150 25072 3149 25088
rect -3150 25008 3065 25072
rect 3129 25008 3149 25072
rect -3150 24992 3149 25008
rect -3150 24928 3065 24992
rect 3129 24928 3149 24992
rect -3150 24912 3149 24928
rect -3150 24848 3065 24912
rect 3129 24848 3149 24912
rect -3150 24832 3149 24848
rect -3150 24768 3065 24832
rect 3129 24768 3149 24832
rect -3150 24752 3149 24768
rect -3150 24688 3065 24752
rect 3129 24688 3149 24752
rect -3150 24672 3149 24688
rect -3150 24608 3065 24672
rect 3129 24608 3149 24672
rect -3150 24592 3149 24608
rect -3150 24528 3065 24592
rect 3129 24528 3149 24592
rect -3150 24512 3149 24528
rect -3150 24448 3065 24512
rect 3129 24448 3149 24512
rect -3150 24432 3149 24448
rect -3150 24368 3065 24432
rect 3129 24368 3149 24432
rect -3150 24352 3149 24368
rect -3150 24288 3065 24352
rect 3129 24288 3149 24352
rect -3150 24272 3149 24288
rect -3150 24208 3065 24272
rect 3129 24208 3149 24272
rect -3150 24192 3149 24208
rect -3150 24128 3065 24192
rect 3129 24128 3149 24192
rect -3150 24112 3149 24128
rect -3150 24048 3065 24112
rect 3129 24048 3149 24112
rect -3150 24032 3149 24048
rect -3150 23968 3065 24032
rect 3129 23968 3149 24032
rect -3150 23952 3149 23968
rect -3150 23888 3065 23952
rect 3129 23888 3149 23952
rect -3150 23872 3149 23888
rect -3150 23808 3065 23872
rect 3129 23808 3149 23872
rect -3150 23792 3149 23808
rect -3150 23728 3065 23792
rect 3129 23728 3149 23792
rect -3150 23712 3149 23728
rect -3150 23648 3065 23712
rect 3129 23648 3149 23712
rect -3150 23632 3149 23648
rect -3150 23568 3065 23632
rect 3129 23568 3149 23632
rect -3150 23552 3149 23568
rect -3150 23488 3065 23552
rect 3129 23488 3149 23552
rect -3150 23472 3149 23488
rect -3150 23408 3065 23472
rect 3129 23408 3149 23472
rect -3150 23392 3149 23408
rect -3150 23328 3065 23392
rect 3129 23328 3149 23392
rect -3150 23312 3149 23328
rect -3150 23248 3065 23312
rect 3129 23248 3149 23312
rect -3150 23232 3149 23248
rect -3150 23168 3065 23232
rect 3129 23168 3149 23232
rect -3150 23152 3149 23168
rect -3150 23088 3065 23152
rect 3129 23088 3149 23152
rect -3150 23072 3149 23088
rect -3150 23008 3065 23072
rect 3129 23008 3149 23072
rect -3150 22992 3149 23008
rect -3150 22928 3065 22992
rect 3129 22928 3149 22992
rect -3150 22912 3149 22928
rect -3150 22848 3065 22912
rect 3129 22848 3149 22912
rect -3150 22832 3149 22848
rect -3150 22768 3065 22832
rect 3129 22768 3149 22832
rect -3150 22752 3149 22768
rect -3150 22688 3065 22752
rect 3129 22688 3149 22752
rect -3150 22672 3149 22688
rect -3150 22608 3065 22672
rect 3129 22608 3149 22672
rect -3150 22592 3149 22608
rect -3150 22528 3065 22592
rect 3129 22528 3149 22592
rect -3150 22512 3149 22528
rect -3150 22448 3065 22512
rect 3129 22448 3149 22512
rect -3150 22432 3149 22448
rect -3150 22368 3065 22432
rect 3129 22368 3149 22432
rect -3150 22352 3149 22368
rect -3150 22288 3065 22352
rect 3129 22288 3149 22352
rect -3150 22272 3149 22288
rect -3150 22208 3065 22272
rect 3129 22208 3149 22272
rect -3150 22192 3149 22208
rect -3150 22128 3065 22192
rect 3129 22128 3149 22192
rect -3150 22100 3149 22128
rect 3169 28272 9468 28300
rect 3169 28208 9384 28272
rect 9448 28208 9468 28272
rect 3169 28192 9468 28208
rect 3169 28128 9384 28192
rect 9448 28128 9468 28192
rect 3169 28112 9468 28128
rect 3169 28048 9384 28112
rect 9448 28048 9468 28112
rect 3169 28032 9468 28048
rect 3169 27968 9384 28032
rect 9448 27968 9468 28032
rect 3169 27952 9468 27968
rect 3169 27888 9384 27952
rect 9448 27888 9468 27952
rect 3169 27872 9468 27888
rect 3169 27808 9384 27872
rect 9448 27808 9468 27872
rect 3169 27792 9468 27808
rect 3169 27728 9384 27792
rect 9448 27728 9468 27792
rect 3169 27712 9468 27728
rect 3169 27648 9384 27712
rect 9448 27648 9468 27712
rect 3169 27632 9468 27648
rect 3169 27568 9384 27632
rect 9448 27568 9468 27632
rect 3169 27552 9468 27568
rect 3169 27488 9384 27552
rect 9448 27488 9468 27552
rect 3169 27472 9468 27488
rect 3169 27408 9384 27472
rect 9448 27408 9468 27472
rect 3169 27392 9468 27408
rect 3169 27328 9384 27392
rect 9448 27328 9468 27392
rect 3169 27312 9468 27328
rect 3169 27248 9384 27312
rect 9448 27248 9468 27312
rect 3169 27232 9468 27248
rect 3169 27168 9384 27232
rect 9448 27168 9468 27232
rect 3169 27152 9468 27168
rect 3169 27088 9384 27152
rect 9448 27088 9468 27152
rect 3169 27072 9468 27088
rect 3169 27008 9384 27072
rect 9448 27008 9468 27072
rect 3169 26992 9468 27008
rect 3169 26928 9384 26992
rect 9448 26928 9468 26992
rect 3169 26912 9468 26928
rect 3169 26848 9384 26912
rect 9448 26848 9468 26912
rect 3169 26832 9468 26848
rect 3169 26768 9384 26832
rect 9448 26768 9468 26832
rect 3169 26752 9468 26768
rect 3169 26688 9384 26752
rect 9448 26688 9468 26752
rect 3169 26672 9468 26688
rect 3169 26608 9384 26672
rect 9448 26608 9468 26672
rect 3169 26592 9468 26608
rect 3169 26528 9384 26592
rect 9448 26528 9468 26592
rect 3169 26512 9468 26528
rect 3169 26448 9384 26512
rect 9448 26448 9468 26512
rect 3169 26432 9468 26448
rect 3169 26368 9384 26432
rect 9448 26368 9468 26432
rect 3169 26352 9468 26368
rect 3169 26288 9384 26352
rect 9448 26288 9468 26352
rect 3169 26272 9468 26288
rect 3169 26208 9384 26272
rect 9448 26208 9468 26272
rect 3169 26192 9468 26208
rect 3169 26128 9384 26192
rect 9448 26128 9468 26192
rect 3169 26112 9468 26128
rect 3169 26048 9384 26112
rect 9448 26048 9468 26112
rect 3169 26032 9468 26048
rect 3169 25968 9384 26032
rect 9448 25968 9468 26032
rect 3169 25952 9468 25968
rect 3169 25888 9384 25952
rect 9448 25888 9468 25952
rect 3169 25872 9468 25888
rect 3169 25808 9384 25872
rect 9448 25808 9468 25872
rect 3169 25792 9468 25808
rect 3169 25728 9384 25792
rect 9448 25728 9468 25792
rect 3169 25712 9468 25728
rect 3169 25648 9384 25712
rect 9448 25648 9468 25712
rect 3169 25632 9468 25648
rect 3169 25568 9384 25632
rect 9448 25568 9468 25632
rect 3169 25552 9468 25568
rect 3169 25488 9384 25552
rect 9448 25488 9468 25552
rect 3169 25472 9468 25488
rect 3169 25408 9384 25472
rect 9448 25408 9468 25472
rect 3169 25392 9468 25408
rect 3169 25328 9384 25392
rect 9448 25328 9468 25392
rect 3169 25312 9468 25328
rect 3169 25248 9384 25312
rect 9448 25248 9468 25312
rect 3169 25232 9468 25248
rect 3169 25168 9384 25232
rect 9448 25168 9468 25232
rect 3169 25152 9468 25168
rect 3169 25088 9384 25152
rect 9448 25088 9468 25152
rect 3169 25072 9468 25088
rect 3169 25008 9384 25072
rect 9448 25008 9468 25072
rect 3169 24992 9468 25008
rect 3169 24928 9384 24992
rect 9448 24928 9468 24992
rect 3169 24912 9468 24928
rect 3169 24848 9384 24912
rect 9448 24848 9468 24912
rect 3169 24832 9468 24848
rect 3169 24768 9384 24832
rect 9448 24768 9468 24832
rect 3169 24752 9468 24768
rect 3169 24688 9384 24752
rect 9448 24688 9468 24752
rect 3169 24672 9468 24688
rect 3169 24608 9384 24672
rect 9448 24608 9468 24672
rect 3169 24592 9468 24608
rect 3169 24528 9384 24592
rect 9448 24528 9468 24592
rect 3169 24512 9468 24528
rect 3169 24448 9384 24512
rect 9448 24448 9468 24512
rect 3169 24432 9468 24448
rect 3169 24368 9384 24432
rect 9448 24368 9468 24432
rect 3169 24352 9468 24368
rect 3169 24288 9384 24352
rect 9448 24288 9468 24352
rect 3169 24272 9468 24288
rect 3169 24208 9384 24272
rect 9448 24208 9468 24272
rect 3169 24192 9468 24208
rect 3169 24128 9384 24192
rect 9448 24128 9468 24192
rect 3169 24112 9468 24128
rect 3169 24048 9384 24112
rect 9448 24048 9468 24112
rect 3169 24032 9468 24048
rect 3169 23968 9384 24032
rect 9448 23968 9468 24032
rect 3169 23952 9468 23968
rect 3169 23888 9384 23952
rect 9448 23888 9468 23952
rect 3169 23872 9468 23888
rect 3169 23808 9384 23872
rect 9448 23808 9468 23872
rect 3169 23792 9468 23808
rect 3169 23728 9384 23792
rect 9448 23728 9468 23792
rect 3169 23712 9468 23728
rect 3169 23648 9384 23712
rect 9448 23648 9468 23712
rect 3169 23632 9468 23648
rect 3169 23568 9384 23632
rect 9448 23568 9468 23632
rect 3169 23552 9468 23568
rect 3169 23488 9384 23552
rect 9448 23488 9468 23552
rect 3169 23472 9468 23488
rect 3169 23408 9384 23472
rect 9448 23408 9468 23472
rect 3169 23392 9468 23408
rect 3169 23328 9384 23392
rect 9448 23328 9468 23392
rect 3169 23312 9468 23328
rect 3169 23248 9384 23312
rect 9448 23248 9468 23312
rect 3169 23232 9468 23248
rect 3169 23168 9384 23232
rect 9448 23168 9468 23232
rect 3169 23152 9468 23168
rect 3169 23088 9384 23152
rect 9448 23088 9468 23152
rect 3169 23072 9468 23088
rect 3169 23008 9384 23072
rect 9448 23008 9468 23072
rect 3169 22992 9468 23008
rect 3169 22928 9384 22992
rect 9448 22928 9468 22992
rect 3169 22912 9468 22928
rect 3169 22848 9384 22912
rect 9448 22848 9468 22912
rect 3169 22832 9468 22848
rect 3169 22768 9384 22832
rect 9448 22768 9468 22832
rect 3169 22752 9468 22768
rect 3169 22688 9384 22752
rect 9448 22688 9468 22752
rect 3169 22672 9468 22688
rect 3169 22608 9384 22672
rect 9448 22608 9468 22672
rect 3169 22592 9468 22608
rect 3169 22528 9384 22592
rect 9448 22528 9468 22592
rect 3169 22512 9468 22528
rect 3169 22448 9384 22512
rect 9448 22448 9468 22512
rect 3169 22432 9468 22448
rect 3169 22368 9384 22432
rect 9448 22368 9468 22432
rect 3169 22352 9468 22368
rect 3169 22288 9384 22352
rect 9448 22288 9468 22352
rect 3169 22272 9468 22288
rect 3169 22208 9384 22272
rect 9448 22208 9468 22272
rect 3169 22192 9468 22208
rect 3169 22128 9384 22192
rect 9448 22128 9468 22192
rect 3169 22100 9468 22128
rect 9488 28272 15787 28300
rect 9488 28208 15703 28272
rect 15767 28208 15787 28272
rect 9488 28192 15787 28208
rect 9488 28128 15703 28192
rect 15767 28128 15787 28192
rect 9488 28112 15787 28128
rect 9488 28048 15703 28112
rect 15767 28048 15787 28112
rect 9488 28032 15787 28048
rect 9488 27968 15703 28032
rect 15767 27968 15787 28032
rect 9488 27952 15787 27968
rect 9488 27888 15703 27952
rect 15767 27888 15787 27952
rect 9488 27872 15787 27888
rect 9488 27808 15703 27872
rect 15767 27808 15787 27872
rect 9488 27792 15787 27808
rect 9488 27728 15703 27792
rect 15767 27728 15787 27792
rect 9488 27712 15787 27728
rect 9488 27648 15703 27712
rect 15767 27648 15787 27712
rect 9488 27632 15787 27648
rect 9488 27568 15703 27632
rect 15767 27568 15787 27632
rect 9488 27552 15787 27568
rect 9488 27488 15703 27552
rect 15767 27488 15787 27552
rect 9488 27472 15787 27488
rect 9488 27408 15703 27472
rect 15767 27408 15787 27472
rect 9488 27392 15787 27408
rect 9488 27328 15703 27392
rect 15767 27328 15787 27392
rect 9488 27312 15787 27328
rect 9488 27248 15703 27312
rect 15767 27248 15787 27312
rect 9488 27232 15787 27248
rect 9488 27168 15703 27232
rect 15767 27168 15787 27232
rect 9488 27152 15787 27168
rect 9488 27088 15703 27152
rect 15767 27088 15787 27152
rect 9488 27072 15787 27088
rect 9488 27008 15703 27072
rect 15767 27008 15787 27072
rect 9488 26992 15787 27008
rect 9488 26928 15703 26992
rect 15767 26928 15787 26992
rect 9488 26912 15787 26928
rect 9488 26848 15703 26912
rect 15767 26848 15787 26912
rect 9488 26832 15787 26848
rect 9488 26768 15703 26832
rect 15767 26768 15787 26832
rect 9488 26752 15787 26768
rect 9488 26688 15703 26752
rect 15767 26688 15787 26752
rect 9488 26672 15787 26688
rect 9488 26608 15703 26672
rect 15767 26608 15787 26672
rect 9488 26592 15787 26608
rect 9488 26528 15703 26592
rect 15767 26528 15787 26592
rect 9488 26512 15787 26528
rect 9488 26448 15703 26512
rect 15767 26448 15787 26512
rect 9488 26432 15787 26448
rect 9488 26368 15703 26432
rect 15767 26368 15787 26432
rect 9488 26352 15787 26368
rect 9488 26288 15703 26352
rect 15767 26288 15787 26352
rect 9488 26272 15787 26288
rect 9488 26208 15703 26272
rect 15767 26208 15787 26272
rect 9488 26192 15787 26208
rect 9488 26128 15703 26192
rect 15767 26128 15787 26192
rect 9488 26112 15787 26128
rect 9488 26048 15703 26112
rect 15767 26048 15787 26112
rect 9488 26032 15787 26048
rect 9488 25968 15703 26032
rect 15767 25968 15787 26032
rect 9488 25952 15787 25968
rect 9488 25888 15703 25952
rect 15767 25888 15787 25952
rect 9488 25872 15787 25888
rect 9488 25808 15703 25872
rect 15767 25808 15787 25872
rect 9488 25792 15787 25808
rect 9488 25728 15703 25792
rect 15767 25728 15787 25792
rect 9488 25712 15787 25728
rect 9488 25648 15703 25712
rect 15767 25648 15787 25712
rect 9488 25632 15787 25648
rect 9488 25568 15703 25632
rect 15767 25568 15787 25632
rect 9488 25552 15787 25568
rect 9488 25488 15703 25552
rect 15767 25488 15787 25552
rect 9488 25472 15787 25488
rect 9488 25408 15703 25472
rect 15767 25408 15787 25472
rect 9488 25392 15787 25408
rect 9488 25328 15703 25392
rect 15767 25328 15787 25392
rect 9488 25312 15787 25328
rect 9488 25248 15703 25312
rect 15767 25248 15787 25312
rect 9488 25232 15787 25248
rect 9488 25168 15703 25232
rect 15767 25168 15787 25232
rect 9488 25152 15787 25168
rect 9488 25088 15703 25152
rect 15767 25088 15787 25152
rect 9488 25072 15787 25088
rect 9488 25008 15703 25072
rect 15767 25008 15787 25072
rect 9488 24992 15787 25008
rect 9488 24928 15703 24992
rect 15767 24928 15787 24992
rect 9488 24912 15787 24928
rect 9488 24848 15703 24912
rect 15767 24848 15787 24912
rect 9488 24832 15787 24848
rect 9488 24768 15703 24832
rect 15767 24768 15787 24832
rect 9488 24752 15787 24768
rect 9488 24688 15703 24752
rect 15767 24688 15787 24752
rect 9488 24672 15787 24688
rect 9488 24608 15703 24672
rect 15767 24608 15787 24672
rect 9488 24592 15787 24608
rect 9488 24528 15703 24592
rect 15767 24528 15787 24592
rect 9488 24512 15787 24528
rect 9488 24448 15703 24512
rect 15767 24448 15787 24512
rect 9488 24432 15787 24448
rect 9488 24368 15703 24432
rect 15767 24368 15787 24432
rect 9488 24352 15787 24368
rect 9488 24288 15703 24352
rect 15767 24288 15787 24352
rect 9488 24272 15787 24288
rect 9488 24208 15703 24272
rect 15767 24208 15787 24272
rect 9488 24192 15787 24208
rect 9488 24128 15703 24192
rect 15767 24128 15787 24192
rect 9488 24112 15787 24128
rect 9488 24048 15703 24112
rect 15767 24048 15787 24112
rect 9488 24032 15787 24048
rect 9488 23968 15703 24032
rect 15767 23968 15787 24032
rect 9488 23952 15787 23968
rect 9488 23888 15703 23952
rect 15767 23888 15787 23952
rect 9488 23872 15787 23888
rect 9488 23808 15703 23872
rect 15767 23808 15787 23872
rect 9488 23792 15787 23808
rect 9488 23728 15703 23792
rect 15767 23728 15787 23792
rect 9488 23712 15787 23728
rect 9488 23648 15703 23712
rect 15767 23648 15787 23712
rect 9488 23632 15787 23648
rect 9488 23568 15703 23632
rect 15767 23568 15787 23632
rect 9488 23552 15787 23568
rect 9488 23488 15703 23552
rect 15767 23488 15787 23552
rect 9488 23472 15787 23488
rect 9488 23408 15703 23472
rect 15767 23408 15787 23472
rect 9488 23392 15787 23408
rect 9488 23328 15703 23392
rect 15767 23328 15787 23392
rect 9488 23312 15787 23328
rect 9488 23248 15703 23312
rect 15767 23248 15787 23312
rect 9488 23232 15787 23248
rect 9488 23168 15703 23232
rect 15767 23168 15787 23232
rect 9488 23152 15787 23168
rect 9488 23088 15703 23152
rect 15767 23088 15787 23152
rect 9488 23072 15787 23088
rect 9488 23008 15703 23072
rect 15767 23008 15787 23072
rect 9488 22992 15787 23008
rect 9488 22928 15703 22992
rect 15767 22928 15787 22992
rect 9488 22912 15787 22928
rect 9488 22848 15703 22912
rect 15767 22848 15787 22912
rect 9488 22832 15787 22848
rect 9488 22768 15703 22832
rect 15767 22768 15787 22832
rect 9488 22752 15787 22768
rect 9488 22688 15703 22752
rect 15767 22688 15787 22752
rect 9488 22672 15787 22688
rect 9488 22608 15703 22672
rect 15767 22608 15787 22672
rect 9488 22592 15787 22608
rect 9488 22528 15703 22592
rect 15767 22528 15787 22592
rect 9488 22512 15787 22528
rect 9488 22448 15703 22512
rect 15767 22448 15787 22512
rect 9488 22432 15787 22448
rect 9488 22368 15703 22432
rect 15767 22368 15787 22432
rect 9488 22352 15787 22368
rect 9488 22288 15703 22352
rect 15767 22288 15787 22352
rect 9488 22272 15787 22288
rect 9488 22208 15703 22272
rect 15767 22208 15787 22272
rect 9488 22192 15787 22208
rect 9488 22128 15703 22192
rect 15767 22128 15787 22192
rect 9488 22100 15787 22128
rect 15807 28272 22106 28300
rect 15807 28208 22022 28272
rect 22086 28208 22106 28272
rect 15807 28192 22106 28208
rect 15807 28128 22022 28192
rect 22086 28128 22106 28192
rect 15807 28112 22106 28128
rect 15807 28048 22022 28112
rect 22086 28048 22106 28112
rect 15807 28032 22106 28048
rect 15807 27968 22022 28032
rect 22086 27968 22106 28032
rect 15807 27952 22106 27968
rect 15807 27888 22022 27952
rect 22086 27888 22106 27952
rect 15807 27872 22106 27888
rect 15807 27808 22022 27872
rect 22086 27808 22106 27872
rect 15807 27792 22106 27808
rect 15807 27728 22022 27792
rect 22086 27728 22106 27792
rect 15807 27712 22106 27728
rect 15807 27648 22022 27712
rect 22086 27648 22106 27712
rect 15807 27632 22106 27648
rect 15807 27568 22022 27632
rect 22086 27568 22106 27632
rect 15807 27552 22106 27568
rect 15807 27488 22022 27552
rect 22086 27488 22106 27552
rect 15807 27472 22106 27488
rect 15807 27408 22022 27472
rect 22086 27408 22106 27472
rect 15807 27392 22106 27408
rect 15807 27328 22022 27392
rect 22086 27328 22106 27392
rect 15807 27312 22106 27328
rect 15807 27248 22022 27312
rect 22086 27248 22106 27312
rect 15807 27232 22106 27248
rect 15807 27168 22022 27232
rect 22086 27168 22106 27232
rect 15807 27152 22106 27168
rect 15807 27088 22022 27152
rect 22086 27088 22106 27152
rect 15807 27072 22106 27088
rect 15807 27008 22022 27072
rect 22086 27008 22106 27072
rect 15807 26992 22106 27008
rect 15807 26928 22022 26992
rect 22086 26928 22106 26992
rect 15807 26912 22106 26928
rect 15807 26848 22022 26912
rect 22086 26848 22106 26912
rect 15807 26832 22106 26848
rect 15807 26768 22022 26832
rect 22086 26768 22106 26832
rect 15807 26752 22106 26768
rect 15807 26688 22022 26752
rect 22086 26688 22106 26752
rect 15807 26672 22106 26688
rect 15807 26608 22022 26672
rect 22086 26608 22106 26672
rect 15807 26592 22106 26608
rect 15807 26528 22022 26592
rect 22086 26528 22106 26592
rect 15807 26512 22106 26528
rect 15807 26448 22022 26512
rect 22086 26448 22106 26512
rect 15807 26432 22106 26448
rect 15807 26368 22022 26432
rect 22086 26368 22106 26432
rect 15807 26352 22106 26368
rect 15807 26288 22022 26352
rect 22086 26288 22106 26352
rect 15807 26272 22106 26288
rect 15807 26208 22022 26272
rect 22086 26208 22106 26272
rect 15807 26192 22106 26208
rect 15807 26128 22022 26192
rect 22086 26128 22106 26192
rect 15807 26112 22106 26128
rect 15807 26048 22022 26112
rect 22086 26048 22106 26112
rect 15807 26032 22106 26048
rect 15807 25968 22022 26032
rect 22086 25968 22106 26032
rect 15807 25952 22106 25968
rect 15807 25888 22022 25952
rect 22086 25888 22106 25952
rect 15807 25872 22106 25888
rect 15807 25808 22022 25872
rect 22086 25808 22106 25872
rect 15807 25792 22106 25808
rect 15807 25728 22022 25792
rect 22086 25728 22106 25792
rect 15807 25712 22106 25728
rect 15807 25648 22022 25712
rect 22086 25648 22106 25712
rect 15807 25632 22106 25648
rect 15807 25568 22022 25632
rect 22086 25568 22106 25632
rect 15807 25552 22106 25568
rect 15807 25488 22022 25552
rect 22086 25488 22106 25552
rect 15807 25472 22106 25488
rect 15807 25408 22022 25472
rect 22086 25408 22106 25472
rect 15807 25392 22106 25408
rect 15807 25328 22022 25392
rect 22086 25328 22106 25392
rect 15807 25312 22106 25328
rect 15807 25248 22022 25312
rect 22086 25248 22106 25312
rect 15807 25232 22106 25248
rect 15807 25168 22022 25232
rect 22086 25168 22106 25232
rect 15807 25152 22106 25168
rect 15807 25088 22022 25152
rect 22086 25088 22106 25152
rect 15807 25072 22106 25088
rect 15807 25008 22022 25072
rect 22086 25008 22106 25072
rect 15807 24992 22106 25008
rect 15807 24928 22022 24992
rect 22086 24928 22106 24992
rect 15807 24912 22106 24928
rect 15807 24848 22022 24912
rect 22086 24848 22106 24912
rect 15807 24832 22106 24848
rect 15807 24768 22022 24832
rect 22086 24768 22106 24832
rect 15807 24752 22106 24768
rect 15807 24688 22022 24752
rect 22086 24688 22106 24752
rect 15807 24672 22106 24688
rect 15807 24608 22022 24672
rect 22086 24608 22106 24672
rect 15807 24592 22106 24608
rect 15807 24528 22022 24592
rect 22086 24528 22106 24592
rect 15807 24512 22106 24528
rect 15807 24448 22022 24512
rect 22086 24448 22106 24512
rect 15807 24432 22106 24448
rect 15807 24368 22022 24432
rect 22086 24368 22106 24432
rect 15807 24352 22106 24368
rect 15807 24288 22022 24352
rect 22086 24288 22106 24352
rect 15807 24272 22106 24288
rect 15807 24208 22022 24272
rect 22086 24208 22106 24272
rect 15807 24192 22106 24208
rect 15807 24128 22022 24192
rect 22086 24128 22106 24192
rect 15807 24112 22106 24128
rect 15807 24048 22022 24112
rect 22086 24048 22106 24112
rect 15807 24032 22106 24048
rect 15807 23968 22022 24032
rect 22086 23968 22106 24032
rect 15807 23952 22106 23968
rect 15807 23888 22022 23952
rect 22086 23888 22106 23952
rect 15807 23872 22106 23888
rect 15807 23808 22022 23872
rect 22086 23808 22106 23872
rect 15807 23792 22106 23808
rect 15807 23728 22022 23792
rect 22086 23728 22106 23792
rect 15807 23712 22106 23728
rect 15807 23648 22022 23712
rect 22086 23648 22106 23712
rect 15807 23632 22106 23648
rect 15807 23568 22022 23632
rect 22086 23568 22106 23632
rect 15807 23552 22106 23568
rect 15807 23488 22022 23552
rect 22086 23488 22106 23552
rect 15807 23472 22106 23488
rect 15807 23408 22022 23472
rect 22086 23408 22106 23472
rect 15807 23392 22106 23408
rect 15807 23328 22022 23392
rect 22086 23328 22106 23392
rect 15807 23312 22106 23328
rect 15807 23248 22022 23312
rect 22086 23248 22106 23312
rect 15807 23232 22106 23248
rect 15807 23168 22022 23232
rect 22086 23168 22106 23232
rect 15807 23152 22106 23168
rect 15807 23088 22022 23152
rect 22086 23088 22106 23152
rect 15807 23072 22106 23088
rect 15807 23008 22022 23072
rect 22086 23008 22106 23072
rect 15807 22992 22106 23008
rect 15807 22928 22022 22992
rect 22086 22928 22106 22992
rect 15807 22912 22106 22928
rect 15807 22848 22022 22912
rect 22086 22848 22106 22912
rect 15807 22832 22106 22848
rect 15807 22768 22022 22832
rect 22086 22768 22106 22832
rect 15807 22752 22106 22768
rect 15807 22688 22022 22752
rect 22086 22688 22106 22752
rect 15807 22672 22106 22688
rect 15807 22608 22022 22672
rect 22086 22608 22106 22672
rect 15807 22592 22106 22608
rect 15807 22528 22022 22592
rect 22086 22528 22106 22592
rect 15807 22512 22106 22528
rect 15807 22448 22022 22512
rect 22086 22448 22106 22512
rect 15807 22432 22106 22448
rect 15807 22368 22022 22432
rect 22086 22368 22106 22432
rect 15807 22352 22106 22368
rect 15807 22288 22022 22352
rect 22086 22288 22106 22352
rect 15807 22272 22106 22288
rect 15807 22208 22022 22272
rect 22086 22208 22106 22272
rect 15807 22192 22106 22208
rect 15807 22128 22022 22192
rect 22086 22128 22106 22192
rect 15807 22100 22106 22128
rect 22126 28272 28425 28300
rect 22126 28208 28341 28272
rect 28405 28208 28425 28272
rect 22126 28192 28425 28208
rect 22126 28128 28341 28192
rect 28405 28128 28425 28192
rect 22126 28112 28425 28128
rect 22126 28048 28341 28112
rect 28405 28048 28425 28112
rect 22126 28032 28425 28048
rect 22126 27968 28341 28032
rect 28405 27968 28425 28032
rect 22126 27952 28425 27968
rect 22126 27888 28341 27952
rect 28405 27888 28425 27952
rect 22126 27872 28425 27888
rect 22126 27808 28341 27872
rect 28405 27808 28425 27872
rect 22126 27792 28425 27808
rect 22126 27728 28341 27792
rect 28405 27728 28425 27792
rect 22126 27712 28425 27728
rect 22126 27648 28341 27712
rect 28405 27648 28425 27712
rect 22126 27632 28425 27648
rect 22126 27568 28341 27632
rect 28405 27568 28425 27632
rect 22126 27552 28425 27568
rect 22126 27488 28341 27552
rect 28405 27488 28425 27552
rect 22126 27472 28425 27488
rect 22126 27408 28341 27472
rect 28405 27408 28425 27472
rect 22126 27392 28425 27408
rect 22126 27328 28341 27392
rect 28405 27328 28425 27392
rect 22126 27312 28425 27328
rect 22126 27248 28341 27312
rect 28405 27248 28425 27312
rect 22126 27232 28425 27248
rect 22126 27168 28341 27232
rect 28405 27168 28425 27232
rect 22126 27152 28425 27168
rect 22126 27088 28341 27152
rect 28405 27088 28425 27152
rect 22126 27072 28425 27088
rect 22126 27008 28341 27072
rect 28405 27008 28425 27072
rect 22126 26992 28425 27008
rect 22126 26928 28341 26992
rect 28405 26928 28425 26992
rect 22126 26912 28425 26928
rect 22126 26848 28341 26912
rect 28405 26848 28425 26912
rect 22126 26832 28425 26848
rect 22126 26768 28341 26832
rect 28405 26768 28425 26832
rect 22126 26752 28425 26768
rect 22126 26688 28341 26752
rect 28405 26688 28425 26752
rect 22126 26672 28425 26688
rect 22126 26608 28341 26672
rect 28405 26608 28425 26672
rect 22126 26592 28425 26608
rect 22126 26528 28341 26592
rect 28405 26528 28425 26592
rect 22126 26512 28425 26528
rect 22126 26448 28341 26512
rect 28405 26448 28425 26512
rect 22126 26432 28425 26448
rect 22126 26368 28341 26432
rect 28405 26368 28425 26432
rect 22126 26352 28425 26368
rect 22126 26288 28341 26352
rect 28405 26288 28425 26352
rect 22126 26272 28425 26288
rect 22126 26208 28341 26272
rect 28405 26208 28425 26272
rect 22126 26192 28425 26208
rect 22126 26128 28341 26192
rect 28405 26128 28425 26192
rect 22126 26112 28425 26128
rect 22126 26048 28341 26112
rect 28405 26048 28425 26112
rect 22126 26032 28425 26048
rect 22126 25968 28341 26032
rect 28405 25968 28425 26032
rect 22126 25952 28425 25968
rect 22126 25888 28341 25952
rect 28405 25888 28425 25952
rect 22126 25872 28425 25888
rect 22126 25808 28341 25872
rect 28405 25808 28425 25872
rect 22126 25792 28425 25808
rect 22126 25728 28341 25792
rect 28405 25728 28425 25792
rect 22126 25712 28425 25728
rect 22126 25648 28341 25712
rect 28405 25648 28425 25712
rect 22126 25632 28425 25648
rect 22126 25568 28341 25632
rect 28405 25568 28425 25632
rect 22126 25552 28425 25568
rect 22126 25488 28341 25552
rect 28405 25488 28425 25552
rect 22126 25472 28425 25488
rect 22126 25408 28341 25472
rect 28405 25408 28425 25472
rect 22126 25392 28425 25408
rect 22126 25328 28341 25392
rect 28405 25328 28425 25392
rect 22126 25312 28425 25328
rect 22126 25248 28341 25312
rect 28405 25248 28425 25312
rect 22126 25232 28425 25248
rect 22126 25168 28341 25232
rect 28405 25168 28425 25232
rect 22126 25152 28425 25168
rect 22126 25088 28341 25152
rect 28405 25088 28425 25152
rect 22126 25072 28425 25088
rect 22126 25008 28341 25072
rect 28405 25008 28425 25072
rect 22126 24992 28425 25008
rect 22126 24928 28341 24992
rect 28405 24928 28425 24992
rect 22126 24912 28425 24928
rect 22126 24848 28341 24912
rect 28405 24848 28425 24912
rect 22126 24832 28425 24848
rect 22126 24768 28341 24832
rect 28405 24768 28425 24832
rect 22126 24752 28425 24768
rect 22126 24688 28341 24752
rect 28405 24688 28425 24752
rect 22126 24672 28425 24688
rect 22126 24608 28341 24672
rect 28405 24608 28425 24672
rect 22126 24592 28425 24608
rect 22126 24528 28341 24592
rect 28405 24528 28425 24592
rect 22126 24512 28425 24528
rect 22126 24448 28341 24512
rect 28405 24448 28425 24512
rect 22126 24432 28425 24448
rect 22126 24368 28341 24432
rect 28405 24368 28425 24432
rect 22126 24352 28425 24368
rect 22126 24288 28341 24352
rect 28405 24288 28425 24352
rect 22126 24272 28425 24288
rect 22126 24208 28341 24272
rect 28405 24208 28425 24272
rect 22126 24192 28425 24208
rect 22126 24128 28341 24192
rect 28405 24128 28425 24192
rect 22126 24112 28425 24128
rect 22126 24048 28341 24112
rect 28405 24048 28425 24112
rect 22126 24032 28425 24048
rect 22126 23968 28341 24032
rect 28405 23968 28425 24032
rect 22126 23952 28425 23968
rect 22126 23888 28341 23952
rect 28405 23888 28425 23952
rect 22126 23872 28425 23888
rect 22126 23808 28341 23872
rect 28405 23808 28425 23872
rect 22126 23792 28425 23808
rect 22126 23728 28341 23792
rect 28405 23728 28425 23792
rect 22126 23712 28425 23728
rect 22126 23648 28341 23712
rect 28405 23648 28425 23712
rect 22126 23632 28425 23648
rect 22126 23568 28341 23632
rect 28405 23568 28425 23632
rect 22126 23552 28425 23568
rect 22126 23488 28341 23552
rect 28405 23488 28425 23552
rect 22126 23472 28425 23488
rect 22126 23408 28341 23472
rect 28405 23408 28425 23472
rect 22126 23392 28425 23408
rect 22126 23328 28341 23392
rect 28405 23328 28425 23392
rect 22126 23312 28425 23328
rect 22126 23248 28341 23312
rect 28405 23248 28425 23312
rect 22126 23232 28425 23248
rect 22126 23168 28341 23232
rect 28405 23168 28425 23232
rect 22126 23152 28425 23168
rect 22126 23088 28341 23152
rect 28405 23088 28425 23152
rect 22126 23072 28425 23088
rect 22126 23008 28341 23072
rect 28405 23008 28425 23072
rect 22126 22992 28425 23008
rect 22126 22928 28341 22992
rect 28405 22928 28425 22992
rect 22126 22912 28425 22928
rect 22126 22848 28341 22912
rect 28405 22848 28425 22912
rect 22126 22832 28425 22848
rect 22126 22768 28341 22832
rect 28405 22768 28425 22832
rect 22126 22752 28425 22768
rect 22126 22688 28341 22752
rect 28405 22688 28425 22752
rect 22126 22672 28425 22688
rect 22126 22608 28341 22672
rect 28405 22608 28425 22672
rect 22126 22592 28425 22608
rect 22126 22528 28341 22592
rect 28405 22528 28425 22592
rect 22126 22512 28425 22528
rect 22126 22448 28341 22512
rect 28405 22448 28425 22512
rect 22126 22432 28425 22448
rect 22126 22368 28341 22432
rect 28405 22368 28425 22432
rect 22126 22352 28425 22368
rect 22126 22288 28341 22352
rect 28405 22288 28425 22352
rect 22126 22272 28425 22288
rect 22126 22208 28341 22272
rect 28405 22208 28425 22272
rect 22126 22192 28425 22208
rect 22126 22128 28341 22192
rect 28405 22128 28425 22192
rect 22126 22100 28425 22128
rect 28445 28272 34744 28300
rect 28445 28208 34660 28272
rect 34724 28208 34744 28272
rect 28445 28192 34744 28208
rect 28445 28128 34660 28192
rect 34724 28128 34744 28192
rect 28445 28112 34744 28128
rect 28445 28048 34660 28112
rect 34724 28048 34744 28112
rect 28445 28032 34744 28048
rect 28445 27968 34660 28032
rect 34724 27968 34744 28032
rect 28445 27952 34744 27968
rect 28445 27888 34660 27952
rect 34724 27888 34744 27952
rect 28445 27872 34744 27888
rect 28445 27808 34660 27872
rect 34724 27808 34744 27872
rect 28445 27792 34744 27808
rect 28445 27728 34660 27792
rect 34724 27728 34744 27792
rect 28445 27712 34744 27728
rect 28445 27648 34660 27712
rect 34724 27648 34744 27712
rect 28445 27632 34744 27648
rect 28445 27568 34660 27632
rect 34724 27568 34744 27632
rect 28445 27552 34744 27568
rect 28445 27488 34660 27552
rect 34724 27488 34744 27552
rect 28445 27472 34744 27488
rect 28445 27408 34660 27472
rect 34724 27408 34744 27472
rect 28445 27392 34744 27408
rect 28445 27328 34660 27392
rect 34724 27328 34744 27392
rect 28445 27312 34744 27328
rect 28445 27248 34660 27312
rect 34724 27248 34744 27312
rect 28445 27232 34744 27248
rect 28445 27168 34660 27232
rect 34724 27168 34744 27232
rect 28445 27152 34744 27168
rect 28445 27088 34660 27152
rect 34724 27088 34744 27152
rect 28445 27072 34744 27088
rect 28445 27008 34660 27072
rect 34724 27008 34744 27072
rect 28445 26992 34744 27008
rect 28445 26928 34660 26992
rect 34724 26928 34744 26992
rect 28445 26912 34744 26928
rect 28445 26848 34660 26912
rect 34724 26848 34744 26912
rect 28445 26832 34744 26848
rect 28445 26768 34660 26832
rect 34724 26768 34744 26832
rect 28445 26752 34744 26768
rect 28445 26688 34660 26752
rect 34724 26688 34744 26752
rect 28445 26672 34744 26688
rect 28445 26608 34660 26672
rect 34724 26608 34744 26672
rect 28445 26592 34744 26608
rect 28445 26528 34660 26592
rect 34724 26528 34744 26592
rect 28445 26512 34744 26528
rect 28445 26448 34660 26512
rect 34724 26448 34744 26512
rect 28445 26432 34744 26448
rect 28445 26368 34660 26432
rect 34724 26368 34744 26432
rect 28445 26352 34744 26368
rect 28445 26288 34660 26352
rect 34724 26288 34744 26352
rect 28445 26272 34744 26288
rect 28445 26208 34660 26272
rect 34724 26208 34744 26272
rect 28445 26192 34744 26208
rect 28445 26128 34660 26192
rect 34724 26128 34744 26192
rect 28445 26112 34744 26128
rect 28445 26048 34660 26112
rect 34724 26048 34744 26112
rect 28445 26032 34744 26048
rect 28445 25968 34660 26032
rect 34724 25968 34744 26032
rect 28445 25952 34744 25968
rect 28445 25888 34660 25952
rect 34724 25888 34744 25952
rect 28445 25872 34744 25888
rect 28445 25808 34660 25872
rect 34724 25808 34744 25872
rect 28445 25792 34744 25808
rect 28445 25728 34660 25792
rect 34724 25728 34744 25792
rect 28445 25712 34744 25728
rect 28445 25648 34660 25712
rect 34724 25648 34744 25712
rect 28445 25632 34744 25648
rect 28445 25568 34660 25632
rect 34724 25568 34744 25632
rect 28445 25552 34744 25568
rect 28445 25488 34660 25552
rect 34724 25488 34744 25552
rect 28445 25472 34744 25488
rect 28445 25408 34660 25472
rect 34724 25408 34744 25472
rect 28445 25392 34744 25408
rect 28445 25328 34660 25392
rect 34724 25328 34744 25392
rect 28445 25312 34744 25328
rect 28445 25248 34660 25312
rect 34724 25248 34744 25312
rect 28445 25232 34744 25248
rect 28445 25168 34660 25232
rect 34724 25168 34744 25232
rect 28445 25152 34744 25168
rect 28445 25088 34660 25152
rect 34724 25088 34744 25152
rect 28445 25072 34744 25088
rect 28445 25008 34660 25072
rect 34724 25008 34744 25072
rect 28445 24992 34744 25008
rect 28445 24928 34660 24992
rect 34724 24928 34744 24992
rect 28445 24912 34744 24928
rect 28445 24848 34660 24912
rect 34724 24848 34744 24912
rect 28445 24832 34744 24848
rect 28445 24768 34660 24832
rect 34724 24768 34744 24832
rect 28445 24752 34744 24768
rect 28445 24688 34660 24752
rect 34724 24688 34744 24752
rect 28445 24672 34744 24688
rect 28445 24608 34660 24672
rect 34724 24608 34744 24672
rect 28445 24592 34744 24608
rect 28445 24528 34660 24592
rect 34724 24528 34744 24592
rect 28445 24512 34744 24528
rect 28445 24448 34660 24512
rect 34724 24448 34744 24512
rect 28445 24432 34744 24448
rect 28445 24368 34660 24432
rect 34724 24368 34744 24432
rect 28445 24352 34744 24368
rect 28445 24288 34660 24352
rect 34724 24288 34744 24352
rect 28445 24272 34744 24288
rect 28445 24208 34660 24272
rect 34724 24208 34744 24272
rect 28445 24192 34744 24208
rect 28445 24128 34660 24192
rect 34724 24128 34744 24192
rect 28445 24112 34744 24128
rect 28445 24048 34660 24112
rect 34724 24048 34744 24112
rect 28445 24032 34744 24048
rect 28445 23968 34660 24032
rect 34724 23968 34744 24032
rect 28445 23952 34744 23968
rect 28445 23888 34660 23952
rect 34724 23888 34744 23952
rect 28445 23872 34744 23888
rect 28445 23808 34660 23872
rect 34724 23808 34744 23872
rect 28445 23792 34744 23808
rect 28445 23728 34660 23792
rect 34724 23728 34744 23792
rect 28445 23712 34744 23728
rect 28445 23648 34660 23712
rect 34724 23648 34744 23712
rect 28445 23632 34744 23648
rect 28445 23568 34660 23632
rect 34724 23568 34744 23632
rect 28445 23552 34744 23568
rect 28445 23488 34660 23552
rect 34724 23488 34744 23552
rect 28445 23472 34744 23488
rect 28445 23408 34660 23472
rect 34724 23408 34744 23472
rect 28445 23392 34744 23408
rect 28445 23328 34660 23392
rect 34724 23328 34744 23392
rect 28445 23312 34744 23328
rect 28445 23248 34660 23312
rect 34724 23248 34744 23312
rect 28445 23232 34744 23248
rect 28445 23168 34660 23232
rect 34724 23168 34744 23232
rect 28445 23152 34744 23168
rect 28445 23088 34660 23152
rect 34724 23088 34744 23152
rect 28445 23072 34744 23088
rect 28445 23008 34660 23072
rect 34724 23008 34744 23072
rect 28445 22992 34744 23008
rect 28445 22928 34660 22992
rect 34724 22928 34744 22992
rect 28445 22912 34744 22928
rect 28445 22848 34660 22912
rect 34724 22848 34744 22912
rect 28445 22832 34744 22848
rect 28445 22768 34660 22832
rect 34724 22768 34744 22832
rect 28445 22752 34744 22768
rect 28445 22688 34660 22752
rect 34724 22688 34744 22752
rect 28445 22672 34744 22688
rect 28445 22608 34660 22672
rect 34724 22608 34744 22672
rect 28445 22592 34744 22608
rect 28445 22528 34660 22592
rect 34724 22528 34744 22592
rect 28445 22512 34744 22528
rect 28445 22448 34660 22512
rect 34724 22448 34744 22512
rect 28445 22432 34744 22448
rect 28445 22368 34660 22432
rect 34724 22368 34744 22432
rect 28445 22352 34744 22368
rect 28445 22288 34660 22352
rect 34724 22288 34744 22352
rect 28445 22272 34744 22288
rect 28445 22208 34660 22272
rect 34724 22208 34744 22272
rect 28445 22192 34744 22208
rect 28445 22128 34660 22192
rect 34724 22128 34744 22192
rect 28445 22100 34744 22128
rect 34764 28272 41063 28300
rect 34764 28208 40979 28272
rect 41043 28208 41063 28272
rect 34764 28192 41063 28208
rect 34764 28128 40979 28192
rect 41043 28128 41063 28192
rect 34764 28112 41063 28128
rect 34764 28048 40979 28112
rect 41043 28048 41063 28112
rect 34764 28032 41063 28048
rect 34764 27968 40979 28032
rect 41043 27968 41063 28032
rect 34764 27952 41063 27968
rect 34764 27888 40979 27952
rect 41043 27888 41063 27952
rect 34764 27872 41063 27888
rect 34764 27808 40979 27872
rect 41043 27808 41063 27872
rect 34764 27792 41063 27808
rect 34764 27728 40979 27792
rect 41043 27728 41063 27792
rect 34764 27712 41063 27728
rect 34764 27648 40979 27712
rect 41043 27648 41063 27712
rect 34764 27632 41063 27648
rect 34764 27568 40979 27632
rect 41043 27568 41063 27632
rect 34764 27552 41063 27568
rect 34764 27488 40979 27552
rect 41043 27488 41063 27552
rect 34764 27472 41063 27488
rect 34764 27408 40979 27472
rect 41043 27408 41063 27472
rect 34764 27392 41063 27408
rect 34764 27328 40979 27392
rect 41043 27328 41063 27392
rect 34764 27312 41063 27328
rect 34764 27248 40979 27312
rect 41043 27248 41063 27312
rect 34764 27232 41063 27248
rect 34764 27168 40979 27232
rect 41043 27168 41063 27232
rect 34764 27152 41063 27168
rect 34764 27088 40979 27152
rect 41043 27088 41063 27152
rect 34764 27072 41063 27088
rect 34764 27008 40979 27072
rect 41043 27008 41063 27072
rect 34764 26992 41063 27008
rect 34764 26928 40979 26992
rect 41043 26928 41063 26992
rect 34764 26912 41063 26928
rect 34764 26848 40979 26912
rect 41043 26848 41063 26912
rect 34764 26832 41063 26848
rect 34764 26768 40979 26832
rect 41043 26768 41063 26832
rect 34764 26752 41063 26768
rect 34764 26688 40979 26752
rect 41043 26688 41063 26752
rect 34764 26672 41063 26688
rect 34764 26608 40979 26672
rect 41043 26608 41063 26672
rect 34764 26592 41063 26608
rect 34764 26528 40979 26592
rect 41043 26528 41063 26592
rect 34764 26512 41063 26528
rect 34764 26448 40979 26512
rect 41043 26448 41063 26512
rect 34764 26432 41063 26448
rect 34764 26368 40979 26432
rect 41043 26368 41063 26432
rect 34764 26352 41063 26368
rect 34764 26288 40979 26352
rect 41043 26288 41063 26352
rect 34764 26272 41063 26288
rect 34764 26208 40979 26272
rect 41043 26208 41063 26272
rect 34764 26192 41063 26208
rect 34764 26128 40979 26192
rect 41043 26128 41063 26192
rect 34764 26112 41063 26128
rect 34764 26048 40979 26112
rect 41043 26048 41063 26112
rect 34764 26032 41063 26048
rect 34764 25968 40979 26032
rect 41043 25968 41063 26032
rect 34764 25952 41063 25968
rect 34764 25888 40979 25952
rect 41043 25888 41063 25952
rect 34764 25872 41063 25888
rect 34764 25808 40979 25872
rect 41043 25808 41063 25872
rect 34764 25792 41063 25808
rect 34764 25728 40979 25792
rect 41043 25728 41063 25792
rect 34764 25712 41063 25728
rect 34764 25648 40979 25712
rect 41043 25648 41063 25712
rect 34764 25632 41063 25648
rect 34764 25568 40979 25632
rect 41043 25568 41063 25632
rect 34764 25552 41063 25568
rect 34764 25488 40979 25552
rect 41043 25488 41063 25552
rect 34764 25472 41063 25488
rect 34764 25408 40979 25472
rect 41043 25408 41063 25472
rect 34764 25392 41063 25408
rect 34764 25328 40979 25392
rect 41043 25328 41063 25392
rect 34764 25312 41063 25328
rect 34764 25248 40979 25312
rect 41043 25248 41063 25312
rect 34764 25232 41063 25248
rect 34764 25168 40979 25232
rect 41043 25168 41063 25232
rect 34764 25152 41063 25168
rect 34764 25088 40979 25152
rect 41043 25088 41063 25152
rect 34764 25072 41063 25088
rect 34764 25008 40979 25072
rect 41043 25008 41063 25072
rect 34764 24992 41063 25008
rect 34764 24928 40979 24992
rect 41043 24928 41063 24992
rect 34764 24912 41063 24928
rect 34764 24848 40979 24912
rect 41043 24848 41063 24912
rect 34764 24832 41063 24848
rect 34764 24768 40979 24832
rect 41043 24768 41063 24832
rect 34764 24752 41063 24768
rect 34764 24688 40979 24752
rect 41043 24688 41063 24752
rect 34764 24672 41063 24688
rect 34764 24608 40979 24672
rect 41043 24608 41063 24672
rect 34764 24592 41063 24608
rect 34764 24528 40979 24592
rect 41043 24528 41063 24592
rect 34764 24512 41063 24528
rect 34764 24448 40979 24512
rect 41043 24448 41063 24512
rect 34764 24432 41063 24448
rect 34764 24368 40979 24432
rect 41043 24368 41063 24432
rect 34764 24352 41063 24368
rect 34764 24288 40979 24352
rect 41043 24288 41063 24352
rect 34764 24272 41063 24288
rect 34764 24208 40979 24272
rect 41043 24208 41063 24272
rect 34764 24192 41063 24208
rect 34764 24128 40979 24192
rect 41043 24128 41063 24192
rect 34764 24112 41063 24128
rect 34764 24048 40979 24112
rect 41043 24048 41063 24112
rect 34764 24032 41063 24048
rect 34764 23968 40979 24032
rect 41043 23968 41063 24032
rect 34764 23952 41063 23968
rect 34764 23888 40979 23952
rect 41043 23888 41063 23952
rect 34764 23872 41063 23888
rect 34764 23808 40979 23872
rect 41043 23808 41063 23872
rect 34764 23792 41063 23808
rect 34764 23728 40979 23792
rect 41043 23728 41063 23792
rect 34764 23712 41063 23728
rect 34764 23648 40979 23712
rect 41043 23648 41063 23712
rect 34764 23632 41063 23648
rect 34764 23568 40979 23632
rect 41043 23568 41063 23632
rect 34764 23552 41063 23568
rect 34764 23488 40979 23552
rect 41043 23488 41063 23552
rect 34764 23472 41063 23488
rect 34764 23408 40979 23472
rect 41043 23408 41063 23472
rect 34764 23392 41063 23408
rect 34764 23328 40979 23392
rect 41043 23328 41063 23392
rect 34764 23312 41063 23328
rect 34764 23248 40979 23312
rect 41043 23248 41063 23312
rect 34764 23232 41063 23248
rect 34764 23168 40979 23232
rect 41043 23168 41063 23232
rect 34764 23152 41063 23168
rect 34764 23088 40979 23152
rect 41043 23088 41063 23152
rect 34764 23072 41063 23088
rect 34764 23008 40979 23072
rect 41043 23008 41063 23072
rect 34764 22992 41063 23008
rect 34764 22928 40979 22992
rect 41043 22928 41063 22992
rect 34764 22912 41063 22928
rect 34764 22848 40979 22912
rect 41043 22848 41063 22912
rect 34764 22832 41063 22848
rect 34764 22768 40979 22832
rect 41043 22768 41063 22832
rect 34764 22752 41063 22768
rect 34764 22688 40979 22752
rect 41043 22688 41063 22752
rect 34764 22672 41063 22688
rect 34764 22608 40979 22672
rect 41043 22608 41063 22672
rect 34764 22592 41063 22608
rect 34764 22528 40979 22592
rect 41043 22528 41063 22592
rect 34764 22512 41063 22528
rect 34764 22448 40979 22512
rect 41043 22448 41063 22512
rect 34764 22432 41063 22448
rect 34764 22368 40979 22432
rect 41043 22368 41063 22432
rect 34764 22352 41063 22368
rect 34764 22288 40979 22352
rect 41043 22288 41063 22352
rect 34764 22272 41063 22288
rect 34764 22208 40979 22272
rect 41043 22208 41063 22272
rect 34764 22192 41063 22208
rect 34764 22128 40979 22192
rect 41043 22128 41063 22192
rect 34764 22100 41063 22128
rect 41083 28272 47382 28300
rect 41083 28208 47298 28272
rect 47362 28208 47382 28272
rect 41083 28192 47382 28208
rect 41083 28128 47298 28192
rect 47362 28128 47382 28192
rect 41083 28112 47382 28128
rect 41083 28048 47298 28112
rect 47362 28048 47382 28112
rect 41083 28032 47382 28048
rect 41083 27968 47298 28032
rect 47362 27968 47382 28032
rect 41083 27952 47382 27968
rect 41083 27888 47298 27952
rect 47362 27888 47382 27952
rect 41083 27872 47382 27888
rect 41083 27808 47298 27872
rect 47362 27808 47382 27872
rect 41083 27792 47382 27808
rect 41083 27728 47298 27792
rect 47362 27728 47382 27792
rect 41083 27712 47382 27728
rect 41083 27648 47298 27712
rect 47362 27648 47382 27712
rect 41083 27632 47382 27648
rect 41083 27568 47298 27632
rect 47362 27568 47382 27632
rect 41083 27552 47382 27568
rect 41083 27488 47298 27552
rect 47362 27488 47382 27552
rect 41083 27472 47382 27488
rect 41083 27408 47298 27472
rect 47362 27408 47382 27472
rect 41083 27392 47382 27408
rect 41083 27328 47298 27392
rect 47362 27328 47382 27392
rect 41083 27312 47382 27328
rect 41083 27248 47298 27312
rect 47362 27248 47382 27312
rect 41083 27232 47382 27248
rect 41083 27168 47298 27232
rect 47362 27168 47382 27232
rect 41083 27152 47382 27168
rect 41083 27088 47298 27152
rect 47362 27088 47382 27152
rect 41083 27072 47382 27088
rect 41083 27008 47298 27072
rect 47362 27008 47382 27072
rect 41083 26992 47382 27008
rect 41083 26928 47298 26992
rect 47362 26928 47382 26992
rect 41083 26912 47382 26928
rect 41083 26848 47298 26912
rect 47362 26848 47382 26912
rect 41083 26832 47382 26848
rect 41083 26768 47298 26832
rect 47362 26768 47382 26832
rect 41083 26752 47382 26768
rect 41083 26688 47298 26752
rect 47362 26688 47382 26752
rect 41083 26672 47382 26688
rect 41083 26608 47298 26672
rect 47362 26608 47382 26672
rect 41083 26592 47382 26608
rect 41083 26528 47298 26592
rect 47362 26528 47382 26592
rect 41083 26512 47382 26528
rect 41083 26448 47298 26512
rect 47362 26448 47382 26512
rect 41083 26432 47382 26448
rect 41083 26368 47298 26432
rect 47362 26368 47382 26432
rect 41083 26352 47382 26368
rect 41083 26288 47298 26352
rect 47362 26288 47382 26352
rect 41083 26272 47382 26288
rect 41083 26208 47298 26272
rect 47362 26208 47382 26272
rect 41083 26192 47382 26208
rect 41083 26128 47298 26192
rect 47362 26128 47382 26192
rect 41083 26112 47382 26128
rect 41083 26048 47298 26112
rect 47362 26048 47382 26112
rect 41083 26032 47382 26048
rect 41083 25968 47298 26032
rect 47362 25968 47382 26032
rect 41083 25952 47382 25968
rect 41083 25888 47298 25952
rect 47362 25888 47382 25952
rect 41083 25872 47382 25888
rect 41083 25808 47298 25872
rect 47362 25808 47382 25872
rect 41083 25792 47382 25808
rect 41083 25728 47298 25792
rect 47362 25728 47382 25792
rect 41083 25712 47382 25728
rect 41083 25648 47298 25712
rect 47362 25648 47382 25712
rect 41083 25632 47382 25648
rect 41083 25568 47298 25632
rect 47362 25568 47382 25632
rect 41083 25552 47382 25568
rect 41083 25488 47298 25552
rect 47362 25488 47382 25552
rect 41083 25472 47382 25488
rect 41083 25408 47298 25472
rect 47362 25408 47382 25472
rect 41083 25392 47382 25408
rect 41083 25328 47298 25392
rect 47362 25328 47382 25392
rect 41083 25312 47382 25328
rect 41083 25248 47298 25312
rect 47362 25248 47382 25312
rect 41083 25232 47382 25248
rect 41083 25168 47298 25232
rect 47362 25168 47382 25232
rect 41083 25152 47382 25168
rect 41083 25088 47298 25152
rect 47362 25088 47382 25152
rect 41083 25072 47382 25088
rect 41083 25008 47298 25072
rect 47362 25008 47382 25072
rect 41083 24992 47382 25008
rect 41083 24928 47298 24992
rect 47362 24928 47382 24992
rect 41083 24912 47382 24928
rect 41083 24848 47298 24912
rect 47362 24848 47382 24912
rect 41083 24832 47382 24848
rect 41083 24768 47298 24832
rect 47362 24768 47382 24832
rect 41083 24752 47382 24768
rect 41083 24688 47298 24752
rect 47362 24688 47382 24752
rect 41083 24672 47382 24688
rect 41083 24608 47298 24672
rect 47362 24608 47382 24672
rect 41083 24592 47382 24608
rect 41083 24528 47298 24592
rect 47362 24528 47382 24592
rect 41083 24512 47382 24528
rect 41083 24448 47298 24512
rect 47362 24448 47382 24512
rect 41083 24432 47382 24448
rect 41083 24368 47298 24432
rect 47362 24368 47382 24432
rect 41083 24352 47382 24368
rect 41083 24288 47298 24352
rect 47362 24288 47382 24352
rect 41083 24272 47382 24288
rect 41083 24208 47298 24272
rect 47362 24208 47382 24272
rect 41083 24192 47382 24208
rect 41083 24128 47298 24192
rect 47362 24128 47382 24192
rect 41083 24112 47382 24128
rect 41083 24048 47298 24112
rect 47362 24048 47382 24112
rect 41083 24032 47382 24048
rect 41083 23968 47298 24032
rect 47362 23968 47382 24032
rect 41083 23952 47382 23968
rect 41083 23888 47298 23952
rect 47362 23888 47382 23952
rect 41083 23872 47382 23888
rect 41083 23808 47298 23872
rect 47362 23808 47382 23872
rect 41083 23792 47382 23808
rect 41083 23728 47298 23792
rect 47362 23728 47382 23792
rect 41083 23712 47382 23728
rect 41083 23648 47298 23712
rect 47362 23648 47382 23712
rect 41083 23632 47382 23648
rect 41083 23568 47298 23632
rect 47362 23568 47382 23632
rect 41083 23552 47382 23568
rect 41083 23488 47298 23552
rect 47362 23488 47382 23552
rect 41083 23472 47382 23488
rect 41083 23408 47298 23472
rect 47362 23408 47382 23472
rect 41083 23392 47382 23408
rect 41083 23328 47298 23392
rect 47362 23328 47382 23392
rect 41083 23312 47382 23328
rect 41083 23248 47298 23312
rect 47362 23248 47382 23312
rect 41083 23232 47382 23248
rect 41083 23168 47298 23232
rect 47362 23168 47382 23232
rect 41083 23152 47382 23168
rect 41083 23088 47298 23152
rect 47362 23088 47382 23152
rect 41083 23072 47382 23088
rect 41083 23008 47298 23072
rect 47362 23008 47382 23072
rect 41083 22992 47382 23008
rect 41083 22928 47298 22992
rect 47362 22928 47382 22992
rect 41083 22912 47382 22928
rect 41083 22848 47298 22912
rect 47362 22848 47382 22912
rect 41083 22832 47382 22848
rect 41083 22768 47298 22832
rect 47362 22768 47382 22832
rect 41083 22752 47382 22768
rect 41083 22688 47298 22752
rect 47362 22688 47382 22752
rect 41083 22672 47382 22688
rect 41083 22608 47298 22672
rect 47362 22608 47382 22672
rect 41083 22592 47382 22608
rect 41083 22528 47298 22592
rect 47362 22528 47382 22592
rect 41083 22512 47382 22528
rect 41083 22448 47298 22512
rect 47362 22448 47382 22512
rect 41083 22432 47382 22448
rect 41083 22368 47298 22432
rect 47362 22368 47382 22432
rect 41083 22352 47382 22368
rect 41083 22288 47298 22352
rect 47362 22288 47382 22352
rect 41083 22272 47382 22288
rect 41083 22208 47298 22272
rect 47362 22208 47382 22272
rect 41083 22192 47382 22208
rect 41083 22128 47298 22192
rect 47362 22128 47382 22192
rect 41083 22100 47382 22128
rect -47383 21972 -41084 22000
rect -47383 21908 -41168 21972
rect -41104 21908 -41084 21972
rect -47383 21892 -41084 21908
rect -47383 21828 -41168 21892
rect -41104 21828 -41084 21892
rect -47383 21812 -41084 21828
rect -47383 21748 -41168 21812
rect -41104 21748 -41084 21812
rect -47383 21732 -41084 21748
rect -47383 21668 -41168 21732
rect -41104 21668 -41084 21732
rect -47383 21652 -41084 21668
rect -47383 21588 -41168 21652
rect -41104 21588 -41084 21652
rect -47383 21572 -41084 21588
rect -47383 21508 -41168 21572
rect -41104 21508 -41084 21572
rect -47383 21492 -41084 21508
rect -47383 21428 -41168 21492
rect -41104 21428 -41084 21492
rect -47383 21412 -41084 21428
rect -47383 21348 -41168 21412
rect -41104 21348 -41084 21412
rect -47383 21332 -41084 21348
rect -47383 21268 -41168 21332
rect -41104 21268 -41084 21332
rect -47383 21252 -41084 21268
rect -47383 21188 -41168 21252
rect -41104 21188 -41084 21252
rect -47383 21172 -41084 21188
rect -47383 21108 -41168 21172
rect -41104 21108 -41084 21172
rect -47383 21092 -41084 21108
rect -47383 21028 -41168 21092
rect -41104 21028 -41084 21092
rect -47383 21012 -41084 21028
rect -47383 20948 -41168 21012
rect -41104 20948 -41084 21012
rect -47383 20932 -41084 20948
rect -47383 20868 -41168 20932
rect -41104 20868 -41084 20932
rect -47383 20852 -41084 20868
rect -47383 20788 -41168 20852
rect -41104 20788 -41084 20852
rect -47383 20772 -41084 20788
rect -47383 20708 -41168 20772
rect -41104 20708 -41084 20772
rect -47383 20692 -41084 20708
rect -47383 20628 -41168 20692
rect -41104 20628 -41084 20692
rect -47383 20612 -41084 20628
rect -47383 20548 -41168 20612
rect -41104 20548 -41084 20612
rect -47383 20532 -41084 20548
rect -47383 20468 -41168 20532
rect -41104 20468 -41084 20532
rect -47383 20452 -41084 20468
rect -47383 20388 -41168 20452
rect -41104 20388 -41084 20452
rect -47383 20372 -41084 20388
rect -47383 20308 -41168 20372
rect -41104 20308 -41084 20372
rect -47383 20292 -41084 20308
rect -47383 20228 -41168 20292
rect -41104 20228 -41084 20292
rect -47383 20212 -41084 20228
rect -47383 20148 -41168 20212
rect -41104 20148 -41084 20212
rect -47383 20132 -41084 20148
rect -47383 20068 -41168 20132
rect -41104 20068 -41084 20132
rect -47383 20052 -41084 20068
rect -47383 19988 -41168 20052
rect -41104 19988 -41084 20052
rect -47383 19972 -41084 19988
rect -47383 19908 -41168 19972
rect -41104 19908 -41084 19972
rect -47383 19892 -41084 19908
rect -47383 19828 -41168 19892
rect -41104 19828 -41084 19892
rect -47383 19812 -41084 19828
rect -47383 19748 -41168 19812
rect -41104 19748 -41084 19812
rect -47383 19732 -41084 19748
rect -47383 19668 -41168 19732
rect -41104 19668 -41084 19732
rect -47383 19652 -41084 19668
rect -47383 19588 -41168 19652
rect -41104 19588 -41084 19652
rect -47383 19572 -41084 19588
rect -47383 19508 -41168 19572
rect -41104 19508 -41084 19572
rect -47383 19492 -41084 19508
rect -47383 19428 -41168 19492
rect -41104 19428 -41084 19492
rect -47383 19412 -41084 19428
rect -47383 19348 -41168 19412
rect -41104 19348 -41084 19412
rect -47383 19332 -41084 19348
rect -47383 19268 -41168 19332
rect -41104 19268 -41084 19332
rect -47383 19252 -41084 19268
rect -47383 19188 -41168 19252
rect -41104 19188 -41084 19252
rect -47383 19172 -41084 19188
rect -47383 19108 -41168 19172
rect -41104 19108 -41084 19172
rect -47383 19092 -41084 19108
rect -47383 19028 -41168 19092
rect -41104 19028 -41084 19092
rect -47383 19012 -41084 19028
rect -47383 18948 -41168 19012
rect -41104 18948 -41084 19012
rect -47383 18932 -41084 18948
rect -47383 18868 -41168 18932
rect -41104 18868 -41084 18932
rect -47383 18852 -41084 18868
rect -47383 18788 -41168 18852
rect -41104 18788 -41084 18852
rect -47383 18772 -41084 18788
rect -47383 18708 -41168 18772
rect -41104 18708 -41084 18772
rect -47383 18692 -41084 18708
rect -47383 18628 -41168 18692
rect -41104 18628 -41084 18692
rect -47383 18612 -41084 18628
rect -47383 18548 -41168 18612
rect -41104 18548 -41084 18612
rect -47383 18532 -41084 18548
rect -47383 18468 -41168 18532
rect -41104 18468 -41084 18532
rect -47383 18452 -41084 18468
rect -47383 18388 -41168 18452
rect -41104 18388 -41084 18452
rect -47383 18372 -41084 18388
rect -47383 18308 -41168 18372
rect -41104 18308 -41084 18372
rect -47383 18292 -41084 18308
rect -47383 18228 -41168 18292
rect -41104 18228 -41084 18292
rect -47383 18212 -41084 18228
rect -47383 18148 -41168 18212
rect -41104 18148 -41084 18212
rect -47383 18132 -41084 18148
rect -47383 18068 -41168 18132
rect -41104 18068 -41084 18132
rect -47383 18052 -41084 18068
rect -47383 17988 -41168 18052
rect -41104 17988 -41084 18052
rect -47383 17972 -41084 17988
rect -47383 17908 -41168 17972
rect -41104 17908 -41084 17972
rect -47383 17892 -41084 17908
rect -47383 17828 -41168 17892
rect -41104 17828 -41084 17892
rect -47383 17812 -41084 17828
rect -47383 17748 -41168 17812
rect -41104 17748 -41084 17812
rect -47383 17732 -41084 17748
rect -47383 17668 -41168 17732
rect -41104 17668 -41084 17732
rect -47383 17652 -41084 17668
rect -47383 17588 -41168 17652
rect -41104 17588 -41084 17652
rect -47383 17572 -41084 17588
rect -47383 17508 -41168 17572
rect -41104 17508 -41084 17572
rect -47383 17492 -41084 17508
rect -47383 17428 -41168 17492
rect -41104 17428 -41084 17492
rect -47383 17412 -41084 17428
rect -47383 17348 -41168 17412
rect -41104 17348 -41084 17412
rect -47383 17332 -41084 17348
rect -47383 17268 -41168 17332
rect -41104 17268 -41084 17332
rect -47383 17252 -41084 17268
rect -47383 17188 -41168 17252
rect -41104 17188 -41084 17252
rect -47383 17172 -41084 17188
rect -47383 17108 -41168 17172
rect -41104 17108 -41084 17172
rect -47383 17092 -41084 17108
rect -47383 17028 -41168 17092
rect -41104 17028 -41084 17092
rect -47383 17012 -41084 17028
rect -47383 16948 -41168 17012
rect -41104 16948 -41084 17012
rect -47383 16932 -41084 16948
rect -47383 16868 -41168 16932
rect -41104 16868 -41084 16932
rect -47383 16852 -41084 16868
rect -47383 16788 -41168 16852
rect -41104 16788 -41084 16852
rect -47383 16772 -41084 16788
rect -47383 16708 -41168 16772
rect -41104 16708 -41084 16772
rect -47383 16692 -41084 16708
rect -47383 16628 -41168 16692
rect -41104 16628 -41084 16692
rect -47383 16612 -41084 16628
rect -47383 16548 -41168 16612
rect -41104 16548 -41084 16612
rect -47383 16532 -41084 16548
rect -47383 16468 -41168 16532
rect -41104 16468 -41084 16532
rect -47383 16452 -41084 16468
rect -47383 16388 -41168 16452
rect -41104 16388 -41084 16452
rect -47383 16372 -41084 16388
rect -47383 16308 -41168 16372
rect -41104 16308 -41084 16372
rect -47383 16292 -41084 16308
rect -47383 16228 -41168 16292
rect -41104 16228 -41084 16292
rect -47383 16212 -41084 16228
rect -47383 16148 -41168 16212
rect -41104 16148 -41084 16212
rect -47383 16132 -41084 16148
rect -47383 16068 -41168 16132
rect -41104 16068 -41084 16132
rect -47383 16052 -41084 16068
rect -47383 15988 -41168 16052
rect -41104 15988 -41084 16052
rect -47383 15972 -41084 15988
rect -47383 15908 -41168 15972
rect -41104 15908 -41084 15972
rect -47383 15892 -41084 15908
rect -47383 15828 -41168 15892
rect -41104 15828 -41084 15892
rect -47383 15800 -41084 15828
rect -41064 21972 -34765 22000
rect -41064 21908 -34849 21972
rect -34785 21908 -34765 21972
rect -41064 21892 -34765 21908
rect -41064 21828 -34849 21892
rect -34785 21828 -34765 21892
rect -41064 21812 -34765 21828
rect -41064 21748 -34849 21812
rect -34785 21748 -34765 21812
rect -41064 21732 -34765 21748
rect -41064 21668 -34849 21732
rect -34785 21668 -34765 21732
rect -41064 21652 -34765 21668
rect -41064 21588 -34849 21652
rect -34785 21588 -34765 21652
rect -41064 21572 -34765 21588
rect -41064 21508 -34849 21572
rect -34785 21508 -34765 21572
rect -41064 21492 -34765 21508
rect -41064 21428 -34849 21492
rect -34785 21428 -34765 21492
rect -41064 21412 -34765 21428
rect -41064 21348 -34849 21412
rect -34785 21348 -34765 21412
rect -41064 21332 -34765 21348
rect -41064 21268 -34849 21332
rect -34785 21268 -34765 21332
rect -41064 21252 -34765 21268
rect -41064 21188 -34849 21252
rect -34785 21188 -34765 21252
rect -41064 21172 -34765 21188
rect -41064 21108 -34849 21172
rect -34785 21108 -34765 21172
rect -41064 21092 -34765 21108
rect -41064 21028 -34849 21092
rect -34785 21028 -34765 21092
rect -41064 21012 -34765 21028
rect -41064 20948 -34849 21012
rect -34785 20948 -34765 21012
rect -41064 20932 -34765 20948
rect -41064 20868 -34849 20932
rect -34785 20868 -34765 20932
rect -41064 20852 -34765 20868
rect -41064 20788 -34849 20852
rect -34785 20788 -34765 20852
rect -41064 20772 -34765 20788
rect -41064 20708 -34849 20772
rect -34785 20708 -34765 20772
rect -41064 20692 -34765 20708
rect -41064 20628 -34849 20692
rect -34785 20628 -34765 20692
rect -41064 20612 -34765 20628
rect -41064 20548 -34849 20612
rect -34785 20548 -34765 20612
rect -41064 20532 -34765 20548
rect -41064 20468 -34849 20532
rect -34785 20468 -34765 20532
rect -41064 20452 -34765 20468
rect -41064 20388 -34849 20452
rect -34785 20388 -34765 20452
rect -41064 20372 -34765 20388
rect -41064 20308 -34849 20372
rect -34785 20308 -34765 20372
rect -41064 20292 -34765 20308
rect -41064 20228 -34849 20292
rect -34785 20228 -34765 20292
rect -41064 20212 -34765 20228
rect -41064 20148 -34849 20212
rect -34785 20148 -34765 20212
rect -41064 20132 -34765 20148
rect -41064 20068 -34849 20132
rect -34785 20068 -34765 20132
rect -41064 20052 -34765 20068
rect -41064 19988 -34849 20052
rect -34785 19988 -34765 20052
rect -41064 19972 -34765 19988
rect -41064 19908 -34849 19972
rect -34785 19908 -34765 19972
rect -41064 19892 -34765 19908
rect -41064 19828 -34849 19892
rect -34785 19828 -34765 19892
rect -41064 19812 -34765 19828
rect -41064 19748 -34849 19812
rect -34785 19748 -34765 19812
rect -41064 19732 -34765 19748
rect -41064 19668 -34849 19732
rect -34785 19668 -34765 19732
rect -41064 19652 -34765 19668
rect -41064 19588 -34849 19652
rect -34785 19588 -34765 19652
rect -41064 19572 -34765 19588
rect -41064 19508 -34849 19572
rect -34785 19508 -34765 19572
rect -41064 19492 -34765 19508
rect -41064 19428 -34849 19492
rect -34785 19428 -34765 19492
rect -41064 19412 -34765 19428
rect -41064 19348 -34849 19412
rect -34785 19348 -34765 19412
rect -41064 19332 -34765 19348
rect -41064 19268 -34849 19332
rect -34785 19268 -34765 19332
rect -41064 19252 -34765 19268
rect -41064 19188 -34849 19252
rect -34785 19188 -34765 19252
rect -41064 19172 -34765 19188
rect -41064 19108 -34849 19172
rect -34785 19108 -34765 19172
rect -41064 19092 -34765 19108
rect -41064 19028 -34849 19092
rect -34785 19028 -34765 19092
rect -41064 19012 -34765 19028
rect -41064 18948 -34849 19012
rect -34785 18948 -34765 19012
rect -41064 18932 -34765 18948
rect -41064 18868 -34849 18932
rect -34785 18868 -34765 18932
rect -41064 18852 -34765 18868
rect -41064 18788 -34849 18852
rect -34785 18788 -34765 18852
rect -41064 18772 -34765 18788
rect -41064 18708 -34849 18772
rect -34785 18708 -34765 18772
rect -41064 18692 -34765 18708
rect -41064 18628 -34849 18692
rect -34785 18628 -34765 18692
rect -41064 18612 -34765 18628
rect -41064 18548 -34849 18612
rect -34785 18548 -34765 18612
rect -41064 18532 -34765 18548
rect -41064 18468 -34849 18532
rect -34785 18468 -34765 18532
rect -41064 18452 -34765 18468
rect -41064 18388 -34849 18452
rect -34785 18388 -34765 18452
rect -41064 18372 -34765 18388
rect -41064 18308 -34849 18372
rect -34785 18308 -34765 18372
rect -41064 18292 -34765 18308
rect -41064 18228 -34849 18292
rect -34785 18228 -34765 18292
rect -41064 18212 -34765 18228
rect -41064 18148 -34849 18212
rect -34785 18148 -34765 18212
rect -41064 18132 -34765 18148
rect -41064 18068 -34849 18132
rect -34785 18068 -34765 18132
rect -41064 18052 -34765 18068
rect -41064 17988 -34849 18052
rect -34785 17988 -34765 18052
rect -41064 17972 -34765 17988
rect -41064 17908 -34849 17972
rect -34785 17908 -34765 17972
rect -41064 17892 -34765 17908
rect -41064 17828 -34849 17892
rect -34785 17828 -34765 17892
rect -41064 17812 -34765 17828
rect -41064 17748 -34849 17812
rect -34785 17748 -34765 17812
rect -41064 17732 -34765 17748
rect -41064 17668 -34849 17732
rect -34785 17668 -34765 17732
rect -41064 17652 -34765 17668
rect -41064 17588 -34849 17652
rect -34785 17588 -34765 17652
rect -41064 17572 -34765 17588
rect -41064 17508 -34849 17572
rect -34785 17508 -34765 17572
rect -41064 17492 -34765 17508
rect -41064 17428 -34849 17492
rect -34785 17428 -34765 17492
rect -41064 17412 -34765 17428
rect -41064 17348 -34849 17412
rect -34785 17348 -34765 17412
rect -41064 17332 -34765 17348
rect -41064 17268 -34849 17332
rect -34785 17268 -34765 17332
rect -41064 17252 -34765 17268
rect -41064 17188 -34849 17252
rect -34785 17188 -34765 17252
rect -41064 17172 -34765 17188
rect -41064 17108 -34849 17172
rect -34785 17108 -34765 17172
rect -41064 17092 -34765 17108
rect -41064 17028 -34849 17092
rect -34785 17028 -34765 17092
rect -41064 17012 -34765 17028
rect -41064 16948 -34849 17012
rect -34785 16948 -34765 17012
rect -41064 16932 -34765 16948
rect -41064 16868 -34849 16932
rect -34785 16868 -34765 16932
rect -41064 16852 -34765 16868
rect -41064 16788 -34849 16852
rect -34785 16788 -34765 16852
rect -41064 16772 -34765 16788
rect -41064 16708 -34849 16772
rect -34785 16708 -34765 16772
rect -41064 16692 -34765 16708
rect -41064 16628 -34849 16692
rect -34785 16628 -34765 16692
rect -41064 16612 -34765 16628
rect -41064 16548 -34849 16612
rect -34785 16548 -34765 16612
rect -41064 16532 -34765 16548
rect -41064 16468 -34849 16532
rect -34785 16468 -34765 16532
rect -41064 16452 -34765 16468
rect -41064 16388 -34849 16452
rect -34785 16388 -34765 16452
rect -41064 16372 -34765 16388
rect -41064 16308 -34849 16372
rect -34785 16308 -34765 16372
rect -41064 16292 -34765 16308
rect -41064 16228 -34849 16292
rect -34785 16228 -34765 16292
rect -41064 16212 -34765 16228
rect -41064 16148 -34849 16212
rect -34785 16148 -34765 16212
rect -41064 16132 -34765 16148
rect -41064 16068 -34849 16132
rect -34785 16068 -34765 16132
rect -41064 16052 -34765 16068
rect -41064 15988 -34849 16052
rect -34785 15988 -34765 16052
rect -41064 15972 -34765 15988
rect -41064 15908 -34849 15972
rect -34785 15908 -34765 15972
rect -41064 15892 -34765 15908
rect -41064 15828 -34849 15892
rect -34785 15828 -34765 15892
rect -41064 15800 -34765 15828
rect -34745 21972 -28446 22000
rect -34745 21908 -28530 21972
rect -28466 21908 -28446 21972
rect -34745 21892 -28446 21908
rect -34745 21828 -28530 21892
rect -28466 21828 -28446 21892
rect -34745 21812 -28446 21828
rect -34745 21748 -28530 21812
rect -28466 21748 -28446 21812
rect -34745 21732 -28446 21748
rect -34745 21668 -28530 21732
rect -28466 21668 -28446 21732
rect -34745 21652 -28446 21668
rect -34745 21588 -28530 21652
rect -28466 21588 -28446 21652
rect -34745 21572 -28446 21588
rect -34745 21508 -28530 21572
rect -28466 21508 -28446 21572
rect -34745 21492 -28446 21508
rect -34745 21428 -28530 21492
rect -28466 21428 -28446 21492
rect -34745 21412 -28446 21428
rect -34745 21348 -28530 21412
rect -28466 21348 -28446 21412
rect -34745 21332 -28446 21348
rect -34745 21268 -28530 21332
rect -28466 21268 -28446 21332
rect -34745 21252 -28446 21268
rect -34745 21188 -28530 21252
rect -28466 21188 -28446 21252
rect -34745 21172 -28446 21188
rect -34745 21108 -28530 21172
rect -28466 21108 -28446 21172
rect -34745 21092 -28446 21108
rect -34745 21028 -28530 21092
rect -28466 21028 -28446 21092
rect -34745 21012 -28446 21028
rect -34745 20948 -28530 21012
rect -28466 20948 -28446 21012
rect -34745 20932 -28446 20948
rect -34745 20868 -28530 20932
rect -28466 20868 -28446 20932
rect -34745 20852 -28446 20868
rect -34745 20788 -28530 20852
rect -28466 20788 -28446 20852
rect -34745 20772 -28446 20788
rect -34745 20708 -28530 20772
rect -28466 20708 -28446 20772
rect -34745 20692 -28446 20708
rect -34745 20628 -28530 20692
rect -28466 20628 -28446 20692
rect -34745 20612 -28446 20628
rect -34745 20548 -28530 20612
rect -28466 20548 -28446 20612
rect -34745 20532 -28446 20548
rect -34745 20468 -28530 20532
rect -28466 20468 -28446 20532
rect -34745 20452 -28446 20468
rect -34745 20388 -28530 20452
rect -28466 20388 -28446 20452
rect -34745 20372 -28446 20388
rect -34745 20308 -28530 20372
rect -28466 20308 -28446 20372
rect -34745 20292 -28446 20308
rect -34745 20228 -28530 20292
rect -28466 20228 -28446 20292
rect -34745 20212 -28446 20228
rect -34745 20148 -28530 20212
rect -28466 20148 -28446 20212
rect -34745 20132 -28446 20148
rect -34745 20068 -28530 20132
rect -28466 20068 -28446 20132
rect -34745 20052 -28446 20068
rect -34745 19988 -28530 20052
rect -28466 19988 -28446 20052
rect -34745 19972 -28446 19988
rect -34745 19908 -28530 19972
rect -28466 19908 -28446 19972
rect -34745 19892 -28446 19908
rect -34745 19828 -28530 19892
rect -28466 19828 -28446 19892
rect -34745 19812 -28446 19828
rect -34745 19748 -28530 19812
rect -28466 19748 -28446 19812
rect -34745 19732 -28446 19748
rect -34745 19668 -28530 19732
rect -28466 19668 -28446 19732
rect -34745 19652 -28446 19668
rect -34745 19588 -28530 19652
rect -28466 19588 -28446 19652
rect -34745 19572 -28446 19588
rect -34745 19508 -28530 19572
rect -28466 19508 -28446 19572
rect -34745 19492 -28446 19508
rect -34745 19428 -28530 19492
rect -28466 19428 -28446 19492
rect -34745 19412 -28446 19428
rect -34745 19348 -28530 19412
rect -28466 19348 -28446 19412
rect -34745 19332 -28446 19348
rect -34745 19268 -28530 19332
rect -28466 19268 -28446 19332
rect -34745 19252 -28446 19268
rect -34745 19188 -28530 19252
rect -28466 19188 -28446 19252
rect -34745 19172 -28446 19188
rect -34745 19108 -28530 19172
rect -28466 19108 -28446 19172
rect -34745 19092 -28446 19108
rect -34745 19028 -28530 19092
rect -28466 19028 -28446 19092
rect -34745 19012 -28446 19028
rect -34745 18948 -28530 19012
rect -28466 18948 -28446 19012
rect -34745 18932 -28446 18948
rect -34745 18868 -28530 18932
rect -28466 18868 -28446 18932
rect -34745 18852 -28446 18868
rect -34745 18788 -28530 18852
rect -28466 18788 -28446 18852
rect -34745 18772 -28446 18788
rect -34745 18708 -28530 18772
rect -28466 18708 -28446 18772
rect -34745 18692 -28446 18708
rect -34745 18628 -28530 18692
rect -28466 18628 -28446 18692
rect -34745 18612 -28446 18628
rect -34745 18548 -28530 18612
rect -28466 18548 -28446 18612
rect -34745 18532 -28446 18548
rect -34745 18468 -28530 18532
rect -28466 18468 -28446 18532
rect -34745 18452 -28446 18468
rect -34745 18388 -28530 18452
rect -28466 18388 -28446 18452
rect -34745 18372 -28446 18388
rect -34745 18308 -28530 18372
rect -28466 18308 -28446 18372
rect -34745 18292 -28446 18308
rect -34745 18228 -28530 18292
rect -28466 18228 -28446 18292
rect -34745 18212 -28446 18228
rect -34745 18148 -28530 18212
rect -28466 18148 -28446 18212
rect -34745 18132 -28446 18148
rect -34745 18068 -28530 18132
rect -28466 18068 -28446 18132
rect -34745 18052 -28446 18068
rect -34745 17988 -28530 18052
rect -28466 17988 -28446 18052
rect -34745 17972 -28446 17988
rect -34745 17908 -28530 17972
rect -28466 17908 -28446 17972
rect -34745 17892 -28446 17908
rect -34745 17828 -28530 17892
rect -28466 17828 -28446 17892
rect -34745 17812 -28446 17828
rect -34745 17748 -28530 17812
rect -28466 17748 -28446 17812
rect -34745 17732 -28446 17748
rect -34745 17668 -28530 17732
rect -28466 17668 -28446 17732
rect -34745 17652 -28446 17668
rect -34745 17588 -28530 17652
rect -28466 17588 -28446 17652
rect -34745 17572 -28446 17588
rect -34745 17508 -28530 17572
rect -28466 17508 -28446 17572
rect -34745 17492 -28446 17508
rect -34745 17428 -28530 17492
rect -28466 17428 -28446 17492
rect -34745 17412 -28446 17428
rect -34745 17348 -28530 17412
rect -28466 17348 -28446 17412
rect -34745 17332 -28446 17348
rect -34745 17268 -28530 17332
rect -28466 17268 -28446 17332
rect -34745 17252 -28446 17268
rect -34745 17188 -28530 17252
rect -28466 17188 -28446 17252
rect -34745 17172 -28446 17188
rect -34745 17108 -28530 17172
rect -28466 17108 -28446 17172
rect -34745 17092 -28446 17108
rect -34745 17028 -28530 17092
rect -28466 17028 -28446 17092
rect -34745 17012 -28446 17028
rect -34745 16948 -28530 17012
rect -28466 16948 -28446 17012
rect -34745 16932 -28446 16948
rect -34745 16868 -28530 16932
rect -28466 16868 -28446 16932
rect -34745 16852 -28446 16868
rect -34745 16788 -28530 16852
rect -28466 16788 -28446 16852
rect -34745 16772 -28446 16788
rect -34745 16708 -28530 16772
rect -28466 16708 -28446 16772
rect -34745 16692 -28446 16708
rect -34745 16628 -28530 16692
rect -28466 16628 -28446 16692
rect -34745 16612 -28446 16628
rect -34745 16548 -28530 16612
rect -28466 16548 -28446 16612
rect -34745 16532 -28446 16548
rect -34745 16468 -28530 16532
rect -28466 16468 -28446 16532
rect -34745 16452 -28446 16468
rect -34745 16388 -28530 16452
rect -28466 16388 -28446 16452
rect -34745 16372 -28446 16388
rect -34745 16308 -28530 16372
rect -28466 16308 -28446 16372
rect -34745 16292 -28446 16308
rect -34745 16228 -28530 16292
rect -28466 16228 -28446 16292
rect -34745 16212 -28446 16228
rect -34745 16148 -28530 16212
rect -28466 16148 -28446 16212
rect -34745 16132 -28446 16148
rect -34745 16068 -28530 16132
rect -28466 16068 -28446 16132
rect -34745 16052 -28446 16068
rect -34745 15988 -28530 16052
rect -28466 15988 -28446 16052
rect -34745 15972 -28446 15988
rect -34745 15908 -28530 15972
rect -28466 15908 -28446 15972
rect -34745 15892 -28446 15908
rect -34745 15828 -28530 15892
rect -28466 15828 -28446 15892
rect -34745 15800 -28446 15828
rect -28426 21972 -22127 22000
rect -28426 21908 -22211 21972
rect -22147 21908 -22127 21972
rect -28426 21892 -22127 21908
rect -28426 21828 -22211 21892
rect -22147 21828 -22127 21892
rect -28426 21812 -22127 21828
rect -28426 21748 -22211 21812
rect -22147 21748 -22127 21812
rect -28426 21732 -22127 21748
rect -28426 21668 -22211 21732
rect -22147 21668 -22127 21732
rect -28426 21652 -22127 21668
rect -28426 21588 -22211 21652
rect -22147 21588 -22127 21652
rect -28426 21572 -22127 21588
rect -28426 21508 -22211 21572
rect -22147 21508 -22127 21572
rect -28426 21492 -22127 21508
rect -28426 21428 -22211 21492
rect -22147 21428 -22127 21492
rect -28426 21412 -22127 21428
rect -28426 21348 -22211 21412
rect -22147 21348 -22127 21412
rect -28426 21332 -22127 21348
rect -28426 21268 -22211 21332
rect -22147 21268 -22127 21332
rect -28426 21252 -22127 21268
rect -28426 21188 -22211 21252
rect -22147 21188 -22127 21252
rect -28426 21172 -22127 21188
rect -28426 21108 -22211 21172
rect -22147 21108 -22127 21172
rect -28426 21092 -22127 21108
rect -28426 21028 -22211 21092
rect -22147 21028 -22127 21092
rect -28426 21012 -22127 21028
rect -28426 20948 -22211 21012
rect -22147 20948 -22127 21012
rect -28426 20932 -22127 20948
rect -28426 20868 -22211 20932
rect -22147 20868 -22127 20932
rect -28426 20852 -22127 20868
rect -28426 20788 -22211 20852
rect -22147 20788 -22127 20852
rect -28426 20772 -22127 20788
rect -28426 20708 -22211 20772
rect -22147 20708 -22127 20772
rect -28426 20692 -22127 20708
rect -28426 20628 -22211 20692
rect -22147 20628 -22127 20692
rect -28426 20612 -22127 20628
rect -28426 20548 -22211 20612
rect -22147 20548 -22127 20612
rect -28426 20532 -22127 20548
rect -28426 20468 -22211 20532
rect -22147 20468 -22127 20532
rect -28426 20452 -22127 20468
rect -28426 20388 -22211 20452
rect -22147 20388 -22127 20452
rect -28426 20372 -22127 20388
rect -28426 20308 -22211 20372
rect -22147 20308 -22127 20372
rect -28426 20292 -22127 20308
rect -28426 20228 -22211 20292
rect -22147 20228 -22127 20292
rect -28426 20212 -22127 20228
rect -28426 20148 -22211 20212
rect -22147 20148 -22127 20212
rect -28426 20132 -22127 20148
rect -28426 20068 -22211 20132
rect -22147 20068 -22127 20132
rect -28426 20052 -22127 20068
rect -28426 19988 -22211 20052
rect -22147 19988 -22127 20052
rect -28426 19972 -22127 19988
rect -28426 19908 -22211 19972
rect -22147 19908 -22127 19972
rect -28426 19892 -22127 19908
rect -28426 19828 -22211 19892
rect -22147 19828 -22127 19892
rect -28426 19812 -22127 19828
rect -28426 19748 -22211 19812
rect -22147 19748 -22127 19812
rect -28426 19732 -22127 19748
rect -28426 19668 -22211 19732
rect -22147 19668 -22127 19732
rect -28426 19652 -22127 19668
rect -28426 19588 -22211 19652
rect -22147 19588 -22127 19652
rect -28426 19572 -22127 19588
rect -28426 19508 -22211 19572
rect -22147 19508 -22127 19572
rect -28426 19492 -22127 19508
rect -28426 19428 -22211 19492
rect -22147 19428 -22127 19492
rect -28426 19412 -22127 19428
rect -28426 19348 -22211 19412
rect -22147 19348 -22127 19412
rect -28426 19332 -22127 19348
rect -28426 19268 -22211 19332
rect -22147 19268 -22127 19332
rect -28426 19252 -22127 19268
rect -28426 19188 -22211 19252
rect -22147 19188 -22127 19252
rect -28426 19172 -22127 19188
rect -28426 19108 -22211 19172
rect -22147 19108 -22127 19172
rect -28426 19092 -22127 19108
rect -28426 19028 -22211 19092
rect -22147 19028 -22127 19092
rect -28426 19012 -22127 19028
rect -28426 18948 -22211 19012
rect -22147 18948 -22127 19012
rect -28426 18932 -22127 18948
rect -28426 18868 -22211 18932
rect -22147 18868 -22127 18932
rect -28426 18852 -22127 18868
rect -28426 18788 -22211 18852
rect -22147 18788 -22127 18852
rect -28426 18772 -22127 18788
rect -28426 18708 -22211 18772
rect -22147 18708 -22127 18772
rect -28426 18692 -22127 18708
rect -28426 18628 -22211 18692
rect -22147 18628 -22127 18692
rect -28426 18612 -22127 18628
rect -28426 18548 -22211 18612
rect -22147 18548 -22127 18612
rect -28426 18532 -22127 18548
rect -28426 18468 -22211 18532
rect -22147 18468 -22127 18532
rect -28426 18452 -22127 18468
rect -28426 18388 -22211 18452
rect -22147 18388 -22127 18452
rect -28426 18372 -22127 18388
rect -28426 18308 -22211 18372
rect -22147 18308 -22127 18372
rect -28426 18292 -22127 18308
rect -28426 18228 -22211 18292
rect -22147 18228 -22127 18292
rect -28426 18212 -22127 18228
rect -28426 18148 -22211 18212
rect -22147 18148 -22127 18212
rect -28426 18132 -22127 18148
rect -28426 18068 -22211 18132
rect -22147 18068 -22127 18132
rect -28426 18052 -22127 18068
rect -28426 17988 -22211 18052
rect -22147 17988 -22127 18052
rect -28426 17972 -22127 17988
rect -28426 17908 -22211 17972
rect -22147 17908 -22127 17972
rect -28426 17892 -22127 17908
rect -28426 17828 -22211 17892
rect -22147 17828 -22127 17892
rect -28426 17812 -22127 17828
rect -28426 17748 -22211 17812
rect -22147 17748 -22127 17812
rect -28426 17732 -22127 17748
rect -28426 17668 -22211 17732
rect -22147 17668 -22127 17732
rect -28426 17652 -22127 17668
rect -28426 17588 -22211 17652
rect -22147 17588 -22127 17652
rect -28426 17572 -22127 17588
rect -28426 17508 -22211 17572
rect -22147 17508 -22127 17572
rect -28426 17492 -22127 17508
rect -28426 17428 -22211 17492
rect -22147 17428 -22127 17492
rect -28426 17412 -22127 17428
rect -28426 17348 -22211 17412
rect -22147 17348 -22127 17412
rect -28426 17332 -22127 17348
rect -28426 17268 -22211 17332
rect -22147 17268 -22127 17332
rect -28426 17252 -22127 17268
rect -28426 17188 -22211 17252
rect -22147 17188 -22127 17252
rect -28426 17172 -22127 17188
rect -28426 17108 -22211 17172
rect -22147 17108 -22127 17172
rect -28426 17092 -22127 17108
rect -28426 17028 -22211 17092
rect -22147 17028 -22127 17092
rect -28426 17012 -22127 17028
rect -28426 16948 -22211 17012
rect -22147 16948 -22127 17012
rect -28426 16932 -22127 16948
rect -28426 16868 -22211 16932
rect -22147 16868 -22127 16932
rect -28426 16852 -22127 16868
rect -28426 16788 -22211 16852
rect -22147 16788 -22127 16852
rect -28426 16772 -22127 16788
rect -28426 16708 -22211 16772
rect -22147 16708 -22127 16772
rect -28426 16692 -22127 16708
rect -28426 16628 -22211 16692
rect -22147 16628 -22127 16692
rect -28426 16612 -22127 16628
rect -28426 16548 -22211 16612
rect -22147 16548 -22127 16612
rect -28426 16532 -22127 16548
rect -28426 16468 -22211 16532
rect -22147 16468 -22127 16532
rect -28426 16452 -22127 16468
rect -28426 16388 -22211 16452
rect -22147 16388 -22127 16452
rect -28426 16372 -22127 16388
rect -28426 16308 -22211 16372
rect -22147 16308 -22127 16372
rect -28426 16292 -22127 16308
rect -28426 16228 -22211 16292
rect -22147 16228 -22127 16292
rect -28426 16212 -22127 16228
rect -28426 16148 -22211 16212
rect -22147 16148 -22127 16212
rect -28426 16132 -22127 16148
rect -28426 16068 -22211 16132
rect -22147 16068 -22127 16132
rect -28426 16052 -22127 16068
rect -28426 15988 -22211 16052
rect -22147 15988 -22127 16052
rect -28426 15972 -22127 15988
rect -28426 15908 -22211 15972
rect -22147 15908 -22127 15972
rect -28426 15892 -22127 15908
rect -28426 15828 -22211 15892
rect -22147 15828 -22127 15892
rect -28426 15800 -22127 15828
rect -22107 21972 -15808 22000
rect -22107 21908 -15892 21972
rect -15828 21908 -15808 21972
rect -22107 21892 -15808 21908
rect -22107 21828 -15892 21892
rect -15828 21828 -15808 21892
rect -22107 21812 -15808 21828
rect -22107 21748 -15892 21812
rect -15828 21748 -15808 21812
rect -22107 21732 -15808 21748
rect -22107 21668 -15892 21732
rect -15828 21668 -15808 21732
rect -22107 21652 -15808 21668
rect -22107 21588 -15892 21652
rect -15828 21588 -15808 21652
rect -22107 21572 -15808 21588
rect -22107 21508 -15892 21572
rect -15828 21508 -15808 21572
rect -22107 21492 -15808 21508
rect -22107 21428 -15892 21492
rect -15828 21428 -15808 21492
rect -22107 21412 -15808 21428
rect -22107 21348 -15892 21412
rect -15828 21348 -15808 21412
rect -22107 21332 -15808 21348
rect -22107 21268 -15892 21332
rect -15828 21268 -15808 21332
rect -22107 21252 -15808 21268
rect -22107 21188 -15892 21252
rect -15828 21188 -15808 21252
rect -22107 21172 -15808 21188
rect -22107 21108 -15892 21172
rect -15828 21108 -15808 21172
rect -22107 21092 -15808 21108
rect -22107 21028 -15892 21092
rect -15828 21028 -15808 21092
rect -22107 21012 -15808 21028
rect -22107 20948 -15892 21012
rect -15828 20948 -15808 21012
rect -22107 20932 -15808 20948
rect -22107 20868 -15892 20932
rect -15828 20868 -15808 20932
rect -22107 20852 -15808 20868
rect -22107 20788 -15892 20852
rect -15828 20788 -15808 20852
rect -22107 20772 -15808 20788
rect -22107 20708 -15892 20772
rect -15828 20708 -15808 20772
rect -22107 20692 -15808 20708
rect -22107 20628 -15892 20692
rect -15828 20628 -15808 20692
rect -22107 20612 -15808 20628
rect -22107 20548 -15892 20612
rect -15828 20548 -15808 20612
rect -22107 20532 -15808 20548
rect -22107 20468 -15892 20532
rect -15828 20468 -15808 20532
rect -22107 20452 -15808 20468
rect -22107 20388 -15892 20452
rect -15828 20388 -15808 20452
rect -22107 20372 -15808 20388
rect -22107 20308 -15892 20372
rect -15828 20308 -15808 20372
rect -22107 20292 -15808 20308
rect -22107 20228 -15892 20292
rect -15828 20228 -15808 20292
rect -22107 20212 -15808 20228
rect -22107 20148 -15892 20212
rect -15828 20148 -15808 20212
rect -22107 20132 -15808 20148
rect -22107 20068 -15892 20132
rect -15828 20068 -15808 20132
rect -22107 20052 -15808 20068
rect -22107 19988 -15892 20052
rect -15828 19988 -15808 20052
rect -22107 19972 -15808 19988
rect -22107 19908 -15892 19972
rect -15828 19908 -15808 19972
rect -22107 19892 -15808 19908
rect -22107 19828 -15892 19892
rect -15828 19828 -15808 19892
rect -22107 19812 -15808 19828
rect -22107 19748 -15892 19812
rect -15828 19748 -15808 19812
rect -22107 19732 -15808 19748
rect -22107 19668 -15892 19732
rect -15828 19668 -15808 19732
rect -22107 19652 -15808 19668
rect -22107 19588 -15892 19652
rect -15828 19588 -15808 19652
rect -22107 19572 -15808 19588
rect -22107 19508 -15892 19572
rect -15828 19508 -15808 19572
rect -22107 19492 -15808 19508
rect -22107 19428 -15892 19492
rect -15828 19428 -15808 19492
rect -22107 19412 -15808 19428
rect -22107 19348 -15892 19412
rect -15828 19348 -15808 19412
rect -22107 19332 -15808 19348
rect -22107 19268 -15892 19332
rect -15828 19268 -15808 19332
rect -22107 19252 -15808 19268
rect -22107 19188 -15892 19252
rect -15828 19188 -15808 19252
rect -22107 19172 -15808 19188
rect -22107 19108 -15892 19172
rect -15828 19108 -15808 19172
rect -22107 19092 -15808 19108
rect -22107 19028 -15892 19092
rect -15828 19028 -15808 19092
rect -22107 19012 -15808 19028
rect -22107 18948 -15892 19012
rect -15828 18948 -15808 19012
rect -22107 18932 -15808 18948
rect -22107 18868 -15892 18932
rect -15828 18868 -15808 18932
rect -22107 18852 -15808 18868
rect -22107 18788 -15892 18852
rect -15828 18788 -15808 18852
rect -22107 18772 -15808 18788
rect -22107 18708 -15892 18772
rect -15828 18708 -15808 18772
rect -22107 18692 -15808 18708
rect -22107 18628 -15892 18692
rect -15828 18628 -15808 18692
rect -22107 18612 -15808 18628
rect -22107 18548 -15892 18612
rect -15828 18548 -15808 18612
rect -22107 18532 -15808 18548
rect -22107 18468 -15892 18532
rect -15828 18468 -15808 18532
rect -22107 18452 -15808 18468
rect -22107 18388 -15892 18452
rect -15828 18388 -15808 18452
rect -22107 18372 -15808 18388
rect -22107 18308 -15892 18372
rect -15828 18308 -15808 18372
rect -22107 18292 -15808 18308
rect -22107 18228 -15892 18292
rect -15828 18228 -15808 18292
rect -22107 18212 -15808 18228
rect -22107 18148 -15892 18212
rect -15828 18148 -15808 18212
rect -22107 18132 -15808 18148
rect -22107 18068 -15892 18132
rect -15828 18068 -15808 18132
rect -22107 18052 -15808 18068
rect -22107 17988 -15892 18052
rect -15828 17988 -15808 18052
rect -22107 17972 -15808 17988
rect -22107 17908 -15892 17972
rect -15828 17908 -15808 17972
rect -22107 17892 -15808 17908
rect -22107 17828 -15892 17892
rect -15828 17828 -15808 17892
rect -22107 17812 -15808 17828
rect -22107 17748 -15892 17812
rect -15828 17748 -15808 17812
rect -22107 17732 -15808 17748
rect -22107 17668 -15892 17732
rect -15828 17668 -15808 17732
rect -22107 17652 -15808 17668
rect -22107 17588 -15892 17652
rect -15828 17588 -15808 17652
rect -22107 17572 -15808 17588
rect -22107 17508 -15892 17572
rect -15828 17508 -15808 17572
rect -22107 17492 -15808 17508
rect -22107 17428 -15892 17492
rect -15828 17428 -15808 17492
rect -22107 17412 -15808 17428
rect -22107 17348 -15892 17412
rect -15828 17348 -15808 17412
rect -22107 17332 -15808 17348
rect -22107 17268 -15892 17332
rect -15828 17268 -15808 17332
rect -22107 17252 -15808 17268
rect -22107 17188 -15892 17252
rect -15828 17188 -15808 17252
rect -22107 17172 -15808 17188
rect -22107 17108 -15892 17172
rect -15828 17108 -15808 17172
rect -22107 17092 -15808 17108
rect -22107 17028 -15892 17092
rect -15828 17028 -15808 17092
rect -22107 17012 -15808 17028
rect -22107 16948 -15892 17012
rect -15828 16948 -15808 17012
rect -22107 16932 -15808 16948
rect -22107 16868 -15892 16932
rect -15828 16868 -15808 16932
rect -22107 16852 -15808 16868
rect -22107 16788 -15892 16852
rect -15828 16788 -15808 16852
rect -22107 16772 -15808 16788
rect -22107 16708 -15892 16772
rect -15828 16708 -15808 16772
rect -22107 16692 -15808 16708
rect -22107 16628 -15892 16692
rect -15828 16628 -15808 16692
rect -22107 16612 -15808 16628
rect -22107 16548 -15892 16612
rect -15828 16548 -15808 16612
rect -22107 16532 -15808 16548
rect -22107 16468 -15892 16532
rect -15828 16468 -15808 16532
rect -22107 16452 -15808 16468
rect -22107 16388 -15892 16452
rect -15828 16388 -15808 16452
rect -22107 16372 -15808 16388
rect -22107 16308 -15892 16372
rect -15828 16308 -15808 16372
rect -22107 16292 -15808 16308
rect -22107 16228 -15892 16292
rect -15828 16228 -15808 16292
rect -22107 16212 -15808 16228
rect -22107 16148 -15892 16212
rect -15828 16148 -15808 16212
rect -22107 16132 -15808 16148
rect -22107 16068 -15892 16132
rect -15828 16068 -15808 16132
rect -22107 16052 -15808 16068
rect -22107 15988 -15892 16052
rect -15828 15988 -15808 16052
rect -22107 15972 -15808 15988
rect -22107 15908 -15892 15972
rect -15828 15908 -15808 15972
rect -22107 15892 -15808 15908
rect -22107 15828 -15892 15892
rect -15828 15828 -15808 15892
rect -22107 15800 -15808 15828
rect -15788 21972 -9489 22000
rect -15788 21908 -9573 21972
rect -9509 21908 -9489 21972
rect -15788 21892 -9489 21908
rect -15788 21828 -9573 21892
rect -9509 21828 -9489 21892
rect -15788 21812 -9489 21828
rect -15788 21748 -9573 21812
rect -9509 21748 -9489 21812
rect -15788 21732 -9489 21748
rect -15788 21668 -9573 21732
rect -9509 21668 -9489 21732
rect -15788 21652 -9489 21668
rect -15788 21588 -9573 21652
rect -9509 21588 -9489 21652
rect -15788 21572 -9489 21588
rect -15788 21508 -9573 21572
rect -9509 21508 -9489 21572
rect -15788 21492 -9489 21508
rect -15788 21428 -9573 21492
rect -9509 21428 -9489 21492
rect -15788 21412 -9489 21428
rect -15788 21348 -9573 21412
rect -9509 21348 -9489 21412
rect -15788 21332 -9489 21348
rect -15788 21268 -9573 21332
rect -9509 21268 -9489 21332
rect -15788 21252 -9489 21268
rect -15788 21188 -9573 21252
rect -9509 21188 -9489 21252
rect -15788 21172 -9489 21188
rect -15788 21108 -9573 21172
rect -9509 21108 -9489 21172
rect -15788 21092 -9489 21108
rect -15788 21028 -9573 21092
rect -9509 21028 -9489 21092
rect -15788 21012 -9489 21028
rect -15788 20948 -9573 21012
rect -9509 20948 -9489 21012
rect -15788 20932 -9489 20948
rect -15788 20868 -9573 20932
rect -9509 20868 -9489 20932
rect -15788 20852 -9489 20868
rect -15788 20788 -9573 20852
rect -9509 20788 -9489 20852
rect -15788 20772 -9489 20788
rect -15788 20708 -9573 20772
rect -9509 20708 -9489 20772
rect -15788 20692 -9489 20708
rect -15788 20628 -9573 20692
rect -9509 20628 -9489 20692
rect -15788 20612 -9489 20628
rect -15788 20548 -9573 20612
rect -9509 20548 -9489 20612
rect -15788 20532 -9489 20548
rect -15788 20468 -9573 20532
rect -9509 20468 -9489 20532
rect -15788 20452 -9489 20468
rect -15788 20388 -9573 20452
rect -9509 20388 -9489 20452
rect -15788 20372 -9489 20388
rect -15788 20308 -9573 20372
rect -9509 20308 -9489 20372
rect -15788 20292 -9489 20308
rect -15788 20228 -9573 20292
rect -9509 20228 -9489 20292
rect -15788 20212 -9489 20228
rect -15788 20148 -9573 20212
rect -9509 20148 -9489 20212
rect -15788 20132 -9489 20148
rect -15788 20068 -9573 20132
rect -9509 20068 -9489 20132
rect -15788 20052 -9489 20068
rect -15788 19988 -9573 20052
rect -9509 19988 -9489 20052
rect -15788 19972 -9489 19988
rect -15788 19908 -9573 19972
rect -9509 19908 -9489 19972
rect -15788 19892 -9489 19908
rect -15788 19828 -9573 19892
rect -9509 19828 -9489 19892
rect -15788 19812 -9489 19828
rect -15788 19748 -9573 19812
rect -9509 19748 -9489 19812
rect -15788 19732 -9489 19748
rect -15788 19668 -9573 19732
rect -9509 19668 -9489 19732
rect -15788 19652 -9489 19668
rect -15788 19588 -9573 19652
rect -9509 19588 -9489 19652
rect -15788 19572 -9489 19588
rect -15788 19508 -9573 19572
rect -9509 19508 -9489 19572
rect -15788 19492 -9489 19508
rect -15788 19428 -9573 19492
rect -9509 19428 -9489 19492
rect -15788 19412 -9489 19428
rect -15788 19348 -9573 19412
rect -9509 19348 -9489 19412
rect -15788 19332 -9489 19348
rect -15788 19268 -9573 19332
rect -9509 19268 -9489 19332
rect -15788 19252 -9489 19268
rect -15788 19188 -9573 19252
rect -9509 19188 -9489 19252
rect -15788 19172 -9489 19188
rect -15788 19108 -9573 19172
rect -9509 19108 -9489 19172
rect -15788 19092 -9489 19108
rect -15788 19028 -9573 19092
rect -9509 19028 -9489 19092
rect -15788 19012 -9489 19028
rect -15788 18948 -9573 19012
rect -9509 18948 -9489 19012
rect -15788 18932 -9489 18948
rect -15788 18868 -9573 18932
rect -9509 18868 -9489 18932
rect -15788 18852 -9489 18868
rect -15788 18788 -9573 18852
rect -9509 18788 -9489 18852
rect -15788 18772 -9489 18788
rect -15788 18708 -9573 18772
rect -9509 18708 -9489 18772
rect -15788 18692 -9489 18708
rect -15788 18628 -9573 18692
rect -9509 18628 -9489 18692
rect -15788 18612 -9489 18628
rect -15788 18548 -9573 18612
rect -9509 18548 -9489 18612
rect -15788 18532 -9489 18548
rect -15788 18468 -9573 18532
rect -9509 18468 -9489 18532
rect -15788 18452 -9489 18468
rect -15788 18388 -9573 18452
rect -9509 18388 -9489 18452
rect -15788 18372 -9489 18388
rect -15788 18308 -9573 18372
rect -9509 18308 -9489 18372
rect -15788 18292 -9489 18308
rect -15788 18228 -9573 18292
rect -9509 18228 -9489 18292
rect -15788 18212 -9489 18228
rect -15788 18148 -9573 18212
rect -9509 18148 -9489 18212
rect -15788 18132 -9489 18148
rect -15788 18068 -9573 18132
rect -9509 18068 -9489 18132
rect -15788 18052 -9489 18068
rect -15788 17988 -9573 18052
rect -9509 17988 -9489 18052
rect -15788 17972 -9489 17988
rect -15788 17908 -9573 17972
rect -9509 17908 -9489 17972
rect -15788 17892 -9489 17908
rect -15788 17828 -9573 17892
rect -9509 17828 -9489 17892
rect -15788 17812 -9489 17828
rect -15788 17748 -9573 17812
rect -9509 17748 -9489 17812
rect -15788 17732 -9489 17748
rect -15788 17668 -9573 17732
rect -9509 17668 -9489 17732
rect -15788 17652 -9489 17668
rect -15788 17588 -9573 17652
rect -9509 17588 -9489 17652
rect -15788 17572 -9489 17588
rect -15788 17508 -9573 17572
rect -9509 17508 -9489 17572
rect -15788 17492 -9489 17508
rect -15788 17428 -9573 17492
rect -9509 17428 -9489 17492
rect -15788 17412 -9489 17428
rect -15788 17348 -9573 17412
rect -9509 17348 -9489 17412
rect -15788 17332 -9489 17348
rect -15788 17268 -9573 17332
rect -9509 17268 -9489 17332
rect -15788 17252 -9489 17268
rect -15788 17188 -9573 17252
rect -9509 17188 -9489 17252
rect -15788 17172 -9489 17188
rect -15788 17108 -9573 17172
rect -9509 17108 -9489 17172
rect -15788 17092 -9489 17108
rect -15788 17028 -9573 17092
rect -9509 17028 -9489 17092
rect -15788 17012 -9489 17028
rect -15788 16948 -9573 17012
rect -9509 16948 -9489 17012
rect -15788 16932 -9489 16948
rect -15788 16868 -9573 16932
rect -9509 16868 -9489 16932
rect -15788 16852 -9489 16868
rect -15788 16788 -9573 16852
rect -9509 16788 -9489 16852
rect -15788 16772 -9489 16788
rect -15788 16708 -9573 16772
rect -9509 16708 -9489 16772
rect -15788 16692 -9489 16708
rect -15788 16628 -9573 16692
rect -9509 16628 -9489 16692
rect -15788 16612 -9489 16628
rect -15788 16548 -9573 16612
rect -9509 16548 -9489 16612
rect -15788 16532 -9489 16548
rect -15788 16468 -9573 16532
rect -9509 16468 -9489 16532
rect -15788 16452 -9489 16468
rect -15788 16388 -9573 16452
rect -9509 16388 -9489 16452
rect -15788 16372 -9489 16388
rect -15788 16308 -9573 16372
rect -9509 16308 -9489 16372
rect -15788 16292 -9489 16308
rect -15788 16228 -9573 16292
rect -9509 16228 -9489 16292
rect -15788 16212 -9489 16228
rect -15788 16148 -9573 16212
rect -9509 16148 -9489 16212
rect -15788 16132 -9489 16148
rect -15788 16068 -9573 16132
rect -9509 16068 -9489 16132
rect -15788 16052 -9489 16068
rect -15788 15988 -9573 16052
rect -9509 15988 -9489 16052
rect -15788 15972 -9489 15988
rect -15788 15908 -9573 15972
rect -9509 15908 -9489 15972
rect -15788 15892 -9489 15908
rect -15788 15828 -9573 15892
rect -9509 15828 -9489 15892
rect -15788 15800 -9489 15828
rect -9469 21972 -3170 22000
rect -9469 21908 -3254 21972
rect -3190 21908 -3170 21972
rect -9469 21892 -3170 21908
rect -9469 21828 -3254 21892
rect -3190 21828 -3170 21892
rect -9469 21812 -3170 21828
rect -9469 21748 -3254 21812
rect -3190 21748 -3170 21812
rect -9469 21732 -3170 21748
rect -9469 21668 -3254 21732
rect -3190 21668 -3170 21732
rect -9469 21652 -3170 21668
rect -9469 21588 -3254 21652
rect -3190 21588 -3170 21652
rect -9469 21572 -3170 21588
rect -9469 21508 -3254 21572
rect -3190 21508 -3170 21572
rect -9469 21492 -3170 21508
rect -9469 21428 -3254 21492
rect -3190 21428 -3170 21492
rect -9469 21412 -3170 21428
rect -9469 21348 -3254 21412
rect -3190 21348 -3170 21412
rect -9469 21332 -3170 21348
rect -9469 21268 -3254 21332
rect -3190 21268 -3170 21332
rect -9469 21252 -3170 21268
rect -9469 21188 -3254 21252
rect -3190 21188 -3170 21252
rect -9469 21172 -3170 21188
rect -9469 21108 -3254 21172
rect -3190 21108 -3170 21172
rect -9469 21092 -3170 21108
rect -9469 21028 -3254 21092
rect -3190 21028 -3170 21092
rect -9469 21012 -3170 21028
rect -9469 20948 -3254 21012
rect -3190 20948 -3170 21012
rect -9469 20932 -3170 20948
rect -9469 20868 -3254 20932
rect -3190 20868 -3170 20932
rect -9469 20852 -3170 20868
rect -9469 20788 -3254 20852
rect -3190 20788 -3170 20852
rect -9469 20772 -3170 20788
rect -9469 20708 -3254 20772
rect -3190 20708 -3170 20772
rect -9469 20692 -3170 20708
rect -9469 20628 -3254 20692
rect -3190 20628 -3170 20692
rect -9469 20612 -3170 20628
rect -9469 20548 -3254 20612
rect -3190 20548 -3170 20612
rect -9469 20532 -3170 20548
rect -9469 20468 -3254 20532
rect -3190 20468 -3170 20532
rect -9469 20452 -3170 20468
rect -9469 20388 -3254 20452
rect -3190 20388 -3170 20452
rect -9469 20372 -3170 20388
rect -9469 20308 -3254 20372
rect -3190 20308 -3170 20372
rect -9469 20292 -3170 20308
rect -9469 20228 -3254 20292
rect -3190 20228 -3170 20292
rect -9469 20212 -3170 20228
rect -9469 20148 -3254 20212
rect -3190 20148 -3170 20212
rect -9469 20132 -3170 20148
rect -9469 20068 -3254 20132
rect -3190 20068 -3170 20132
rect -9469 20052 -3170 20068
rect -9469 19988 -3254 20052
rect -3190 19988 -3170 20052
rect -9469 19972 -3170 19988
rect -9469 19908 -3254 19972
rect -3190 19908 -3170 19972
rect -9469 19892 -3170 19908
rect -9469 19828 -3254 19892
rect -3190 19828 -3170 19892
rect -9469 19812 -3170 19828
rect -9469 19748 -3254 19812
rect -3190 19748 -3170 19812
rect -9469 19732 -3170 19748
rect -9469 19668 -3254 19732
rect -3190 19668 -3170 19732
rect -9469 19652 -3170 19668
rect -9469 19588 -3254 19652
rect -3190 19588 -3170 19652
rect -9469 19572 -3170 19588
rect -9469 19508 -3254 19572
rect -3190 19508 -3170 19572
rect -9469 19492 -3170 19508
rect -9469 19428 -3254 19492
rect -3190 19428 -3170 19492
rect -9469 19412 -3170 19428
rect -9469 19348 -3254 19412
rect -3190 19348 -3170 19412
rect -9469 19332 -3170 19348
rect -9469 19268 -3254 19332
rect -3190 19268 -3170 19332
rect -9469 19252 -3170 19268
rect -9469 19188 -3254 19252
rect -3190 19188 -3170 19252
rect -9469 19172 -3170 19188
rect -9469 19108 -3254 19172
rect -3190 19108 -3170 19172
rect -9469 19092 -3170 19108
rect -9469 19028 -3254 19092
rect -3190 19028 -3170 19092
rect -9469 19012 -3170 19028
rect -9469 18948 -3254 19012
rect -3190 18948 -3170 19012
rect -9469 18932 -3170 18948
rect -9469 18868 -3254 18932
rect -3190 18868 -3170 18932
rect -9469 18852 -3170 18868
rect -9469 18788 -3254 18852
rect -3190 18788 -3170 18852
rect -9469 18772 -3170 18788
rect -9469 18708 -3254 18772
rect -3190 18708 -3170 18772
rect -9469 18692 -3170 18708
rect -9469 18628 -3254 18692
rect -3190 18628 -3170 18692
rect -9469 18612 -3170 18628
rect -9469 18548 -3254 18612
rect -3190 18548 -3170 18612
rect -9469 18532 -3170 18548
rect -9469 18468 -3254 18532
rect -3190 18468 -3170 18532
rect -9469 18452 -3170 18468
rect -9469 18388 -3254 18452
rect -3190 18388 -3170 18452
rect -9469 18372 -3170 18388
rect -9469 18308 -3254 18372
rect -3190 18308 -3170 18372
rect -9469 18292 -3170 18308
rect -9469 18228 -3254 18292
rect -3190 18228 -3170 18292
rect -9469 18212 -3170 18228
rect -9469 18148 -3254 18212
rect -3190 18148 -3170 18212
rect -9469 18132 -3170 18148
rect -9469 18068 -3254 18132
rect -3190 18068 -3170 18132
rect -9469 18052 -3170 18068
rect -9469 17988 -3254 18052
rect -3190 17988 -3170 18052
rect -9469 17972 -3170 17988
rect -9469 17908 -3254 17972
rect -3190 17908 -3170 17972
rect -9469 17892 -3170 17908
rect -9469 17828 -3254 17892
rect -3190 17828 -3170 17892
rect -9469 17812 -3170 17828
rect -9469 17748 -3254 17812
rect -3190 17748 -3170 17812
rect -9469 17732 -3170 17748
rect -9469 17668 -3254 17732
rect -3190 17668 -3170 17732
rect -9469 17652 -3170 17668
rect -9469 17588 -3254 17652
rect -3190 17588 -3170 17652
rect -9469 17572 -3170 17588
rect -9469 17508 -3254 17572
rect -3190 17508 -3170 17572
rect -9469 17492 -3170 17508
rect -9469 17428 -3254 17492
rect -3190 17428 -3170 17492
rect -9469 17412 -3170 17428
rect -9469 17348 -3254 17412
rect -3190 17348 -3170 17412
rect -9469 17332 -3170 17348
rect -9469 17268 -3254 17332
rect -3190 17268 -3170 17332
rect -9469 17252 -3170 17268
rect -9469 17188 -3254 17252
rect -3190 17188 -3170 17252
rect -9469 17172 -3170 17188
rect -9469 17108 -3254 17172
rect -3190 17108 -3170 17172
rect -9469 17092 -3170 17108
rect -9469 17028 -3254 17092
rect -3190 17028 -3170 17092
rect -9469 17012 -3170 17028
rect -9469 16948 -3254 17012
rect -3190 16948 -3170 17012
rect -9469 16932 -3170 16948
rect -9469 16868 -3254 16932
rect -3190 16868 -3170 16932
rect -9469 16852 -3170 16868
rect -9469 16788 -3254 16852
rect -3190 16788 -3170 16852
rect -9469 16772 -3170 16788
rect -9469 16708 -3254 16772
rect -3190 16708 -3170 16772
rect -9469 16692 -3170 16708
rect -9469 16628 -3254 16692
rect -3190 16628 -3170 16692
rect -9469 16612 -3170 16628
rect -9469 16548 -3254 16612
rect -3190 16548 -3170 16612
rect -9469 16532 -3170 16548
rect -9469 16468 -3254 16532
rect -3190 16468 -3170 16532
rect -9469 16452 -3170 16468
rect -9469 16388 -3254 16452
rect -3190 16388 -3170 16452
rect -9469 16372 -3170 16388
rect -9469 16308 -3254 16372
rect -3190 16308 -3170 16372
rect -9469 16292 -3170 16308
rect -9469 16228 -3254 16292
rect -3190 16228 -3170 16292
rect -9469 16212 -3170 16228
rect -9469 16148 -3254 16212
rect -3190 16148 -3170 16212
rect -9469 16132 -3170 16148
rect -9469 16068 -3254 16132
rect -3190 16068 -3170 16132
rect -9469 16052 -3170 16068
rect -9469 15988 -3254 16052
rect -3190 15988 -3170 16052
rect -9469 15972 -3170 15988
rect -9469 15908 -3254 15972
rect -3190 15908 -3170 15972
rect -9469 15892 -3170 15908
rect -9469 15828 -3254 15892
rect -3190 15828 -3170 15892
rect -9469 15800 -3170 15828
rect -3150 21972 3149 22000
rect -3150 21908 3065 21972
rect 3129 21908 3149 21972
rect -3150 21892 3149 21908
rect -3150 21828 3065 21892
rect 3129 21828 3149 21892
rect -3150 21812 3149 21828
rect -3150 21748 3065 21812
rect 3129 21748 3149 21812
rect -3150 21732 3149 21748
rect -3150 21668 3065 21732
rect 3129 21668 3149 21732
rect -3150 21652 3149 21668
rect -3150 21588 3065 21652
rect 3129 21588 3149 21652
rect -3150 21572 3149 21588
rect -3150 21508 3065 21572
rect 3129 21508 3149 21572
rect -3150 21492 3149 21508
rect -3150 21428 3065 21492
rect 3129 21428 3149 21492
rect -3150 21412 3149 21428
rect -3150 21348 3065 21412
rect 3129 21348 3149 21412
rect -3150 21332 3149 21348
rect -3150 21268 3065 21332
rect 3129 21268 3149 21332
rect -3150 21252 3149 21268
rect -3150 21188 3065 21252
rect 3129 21188 3149 21252
rect -3150 21172 3149 21188
rect -3150 21108 3065 21172
rect 3129 21108 3149 21172
rect -3150 21092 3149 21108
rect -3150 21028 3065 21092
rect 3129 21028 3149 21092
rect -3150 21012 3149 21028
rect -3150 20948 3065 21012
rect 3129 20948 3149 21012
rect -3150 20932 3149 20948
rect -3150 20868 3065 20932
rect 3129 20868 3149 20932
rect -3150 20852 3149 20868
rect -3150 20788 3065 20852
rect 3129 20788 3149 20852
rect -3150 20772 3149 20788
rect -3150 20708 3065 20772
rect 3129 20708 3149 20772
rect -3150 20692 3149 20708
rect -3150 20628 3065 20692
rect 3129 20628 3149 20692
rect -3150 20612 3149 20628
rect -3150 20548 3065 20612
rect 3129 20548 3149 20612
rect -3150 20532 3149 20548
rect -3150 20468 3065 20532
rect 3129 20468 3149 20532
rect -3150 20452 3149 20468
rect -3150 20388 3065 20452
rect 3129 20388 3149 20452
rect -3150 20372 3149 20388
rect -3150 20308 3065 20372
rect 3129 20308 3149 20372
rect -3150 20292 3149 20308
rect -3150 20228 3065 20292
rect 3129 20228 3149 20292
rect -3150 20212 3149 20228
rect -3150 20148 3065 20212
rect 3129 20148 3149 20212
rect -3150 20132 3149 20148
rect -3150 20068 3065 20132
rect 3129 20068 3149 20132
rect -3150 20052 3149 20068
rect -3150 19988 3065 20052
rect 3129 19988 3149 20052
rect -3150 19972 3149 19988
rect -3150 19908 3065 19972
rect 3129 19908 3149 19972
rect -3150 19892 3149 19908
rect -3150 19828 3065 19892
rect 3129 19828 3149 19892
rect -3150 19812 3149 19828
rect -3150 19748 3065 19812
rect 3129 19748 3149 19812
rect -3150 19732 3149 19748
rect -3150 19668 3065 19732
rect 3129 19668 3149 19732
rect -3150 19652 3149 19668
rect -3150 19588 3065 19652
rect 3129 19588 3149 19652
rect -3150 19572 3149 19588
rect -3150 19508 3065 19572
rect 3129 19508 3149 19572
rect -3150 19492 3149 19508
rect -3150 19428 3065 19492
rect 3129 19428 3149 19492
rect -3150 19412 3149 19428
rect -3150 19348 3065 19412
rect 3129 19348 3149 19412
rect -3150 19332 3149 19348
rect -3150 19268 3065 19332
rect 3129 19268 3149 19332
rect -3150 19252 3149 19268
rect -3150 19188 3065 19252
rect 3129 19188 3149 19252
rect -3150 19172 3149 19188
rect -3150 19108 3065 19172
rect 3129 19108 3149 19172
rect -3150 19092 3149 19108
rect -3150 19028 3065 19092
rect 3129 19028 3149 19092
rect -3150 19012 3149 19028
rect -3150 18948 3065 19012
rect 3129 18948 3149 19012
rect -3150 18932 3149 18948
rect -3150 18868 3065 18932
rect 3129 18868 3149 18932
rect -3150 18852 3149 18868
rect -3150 18788 3065 18852
rect 3129 18788 3149 18852
rect -3150 18772 3149 18788
rect -3150 18708 3065 18772
rect 3129 18708 3149 18772
rect -3150 18692 3149 18708
rect -3150 18628 3065 18692
rect 3129 18628 3149 18692
rect -3150 18612 3149 18628
rect -3150 18548 3065 18612
rect 3129 18548 3149 18612
rect -3150 18532 3149 18548
rect -3150 18468 3065 18532
rect 3129 18468 3149 18532
rect -3150 18452 3149 18468
rect -3150 18388 3065 18452
rect 3129 18388 3149 18452
rect -3150 18372 3149 18388
rect -3150 18308 3065 18372
rect 3129 18308 3149 18372
rect -3150 18292 3149 18308
rect -3150 18228 3065 18292
rect 3129 18228 3149 18292
rect -3150 18212 3149 18228
rect -3150 18148 3065 18212
rect 3129 18148 3149 18212
rect -3150 18132 3149 18148
rect -3150 18068 3065 18132
rect 3129 18068 3149 18132
rect -3150 18052 3149 18068
rect -3150 17988 3065 18052
rect 3129 17988 3149 18052
rect -3150 17972 3149 17988
rect -3150 17908 3065 17972
rect 3129 17908 3149 17972
rect -3150 17892 3149 17908
rect -3150 17828 3065 17892
rect 3129 17828 3149 17892
rect -3150 17812 3149 17828
rect -3150 17748 3065 17812
rect 3129 17748 3149 17812
rect -3150 17732 3149 17748
rect -3150 17668 3065 17732
rect 3129 17668 3149 17732
rect -3150 17652 3149 17668
rect -3150 17588 3065 17652
rect 3129 17588 3149 17652
rect -3150 17572 3149 17588
rect -3150 17508 3065 17572
rect 3129 17508 3149 17572
rect -3150 17492 3149 17508
rect -3150 17428 3065 17492
rect 3129 17428 3149 17492
rect -3150 17412 3149 17428
rect -3150 17348 3065 17412
rect 3129 17348 3149 17412
rect -3150 17332 3149 17348
rect -3150 17268 3065 17332
rect 3129 17268 3149 17332
rect -3150 17252 3149 17268
rect -3150 17188 3065 17252
rect 3129 17188 3149 17252
rect -3150 17172 3149 17188
rect -3150 17108 3065 17172
rect 3129 17108 3149 17172
rect -3150 17092 3149 17108
rect -3150 17028 3065 17092
rect 3129 17028 3149 17092
rect -3150 17012 3149 17028
rect -3150 16948 3065 17012
rect 3129 16948 3149 17012
rect -3150 16932 3149 16948
rect -3150 16868 3065 16932
rect 3129 16868 3149 16932
rect -3150 16852 3149 16868
rect -3150 16788 3065 16852
rect 3129 16788 3149 16852
rect -3150 16772 3149 16788
rect -3150 16708 3065 16772
rect 3129 16708 3149 16772
rect -3150 16692 3149 16708
rect -3150 16628 3065 16692
rect 3129 16628 3149 16692
rect -3150 16612 3149 16628
rect -3150 16548 3065 16612
rect 3129 16548 3149 16612
rect -3150 16532 3149 16548
rect -3150 16468 3065 16532
rect 3129 16468 3149 16532
rect -3150 16452 3149 16468
rect -3150 16388 3065 16452
rect 3129 16388 3149 16452
rect -3150 16372 3149 16388
rect -3150 16308 3065 16372
rect 3129 16308 3149 16372
rect -3150 16292 3149 16308
rect -3150 16228 3065 16292
rect 3129 16228 3149 16292
rect -3150 16212 3149 16228
rect -3150 16148 3065 16212
rect 3129 16148 3149 16212
rect -3150 16132 3149 16148
rect -3150 16068 3065 16132
rect 3129 16068 3149 16132
rect -3150 16052 3149 16068
rect -3150 15988 3065 16052
rect 3129 15988 3149 16052
rect -3150 15972 3149 15988
rect -3150 15908 3065 15972
rect 3129 15908 3149 15972
rect -3150 15892 3149 15908
rect -3150 15828 3065 15892
rect 3129 15828 3149 15892
rect -3150 15800 3149 15828
rect 3169 21972 9468 22000
rect 3169 21908 9384 21972
rect 9448 21908 9468 21972
rect 3169 21892 9468 21908
rect 3169 21828 9384 21892
rect 9448 21828 9468 21892
rect 3169 21812 9468 21828
rect 3169 21748 9384 21812
rect 9448 21748 9468 21812
rect 3169 21732 9468 21748
rect 3169 21668 9384 21732
rect 9448 21668 9468 21732
rect 3169 21652 9468 21668
rect 3169 21588 9384 21652
rect 9448 21588 9468 21652
rect 3169 21572 9468 21588
rect 3169 21508 9384 21572
rect 9448 21508 9468 21572
rect 3169 21492 9468 21508
rect 3169 21428 9384 21492
rect 9448 21428 9468 21492
rect 3169 21412 9468 21428
rect 3169 21348 9384 21412
rect 9448 21348 9468 21412
rect 3169 21332 9468 21348
rect 3169 21268 9384 21332
rect 9448 21268 9468 21332
rect 3169 21252 9468 21268
rect 3169 21188 9384 21252
rect 9448 21188 9468 21252
rect 3169 21172 9468 21188
rect 3169 21108 9384 21172
rect 9448 21108 9468 21172
rect 3169 21092 9468 21108
rect 3169 21028 9384 21092
rect 9448 21028 9468 21092
rect 3169 21012 9468 21028
rect 3169 20948 9384 21012
rect 9448 20948 9468 21012
rect 3169 20932 9468 20948
rect 3169 20868 9384 20932
rect 9448 20868 9468 20932
rect 3169 20852 9468 20868
rect 3169 20788 9384 20852
rect 9448 20788 9468 20852
rect 3169 20772 9468 20788
rect 3169 20708 9384 20772
rect 9448 20708 9468 20772
rect 3169 20692 9468 20708
rect 3169 20628 9384 20692
rect 9448 20628 9468 20692
rect 3169 20612 9468 20628
rect 3169 20548 9384 20612
rect 9448 20548 9468 20612
rect 3169 20532 9468 20548
rect 3169 20468 9384 20532
rect 9448 20468 9468 20532
rect 3169 20452 9468 20468
rect 3169 20388 9384 20452
rect 9448 20388 9468 20452
rect 3169 20372 9468 20388
rect 3169 20308 9384 20372
rect 9448 20308 9468 20372
rect 3169 20292 9468 20308
rect 3169 20228 9384 20292
rect 9448 20228 9468 20292
rect 3169 20212 9468 20228
rect 3169 20148 9384 20212
rect 9448 20148 9468 20212
rect 3169 20132 9468 20148
rect 3169 20068 9384 20132
rect 9448 20068 9468 20132
rect 3169 20052 9468 20068
rect 3169 19988 9384 20052
rect 9448 19988 9468 20052
rect 3169 19972 9468 19988
rect 3169 19908 9384 19972
rect 9448 19908 9468 19972
rect 3169 19892 9468 19908
rect 3169 19828 9384 19892
rect 9448 19828 9468 19892
rect 3169 19812 9468 19828
rect 3169 19748 9384 19812
rect 9448 19748 9468 19812
rect 3169 19732 9468 19748
rect 3169 19668 9384 19732
rect 9448 19668 9468 19732
rect 3169 19652 9468 19668
rect 3169 19588 9384 19652
rect 9448 19588 9468 19652
rect 3169 19572 9468 19588
rect 3169 19508 9384 19572
rect 9448 19508 9468 19572
rect 3169 19492 9468 19508
rect 3169 19428 9384 19492
rect 9448 19428 9468 19492
rect 3169 19412 9468 19428
rect 3169 19348 9384 19412
rect 9448 19348 9468 19412
rect 3169 19332 9468 19348
rect 3169 19268 9384 19332
rect 9448 19268 9468 19332
rect 3169 19252 9468 19268
rect 3169 19188 9384 19252
rect 9448 19188 9468 19252
rect 3169 19172 9468 19188
rect 3169 19108 9384 19172
rect 9448 19108 9468 19172
rect 3169 19092 9468 19108
rect 3169 19028 9384 19092
rect 9448 19028 9468 19092
rect 3169 19012 9468 19028
rect 3169 18948 9384 19012
rect 9448 18948 9468 19012
rect 3169 18932 9468 18948
rect 3169 18868 9384 18932
rect 9448 18868 9468 18932
rect 3169 18852 9468 18868
rect 3169 18788 9384 18852
rect 9448 18788 9468 18852
rect 3169 18772 9468 18788
rect 3169 18708 9384 18772
rect 9448 18708 9468 18772
rect 3169 18692 9468 18708
rect 3169 18628 9384 18692
rect 9448 18628 9468 18692
rect 3169 18612 9468 18628
rect 3169 18548 9384 18612
rect 9448 18548 9468 18612
rect 3169 18532 9468 18548
rect 3169 18468 9384 18532
rect 9448 18468 9468 18532
rect 3169 18452 9468 18468
rect 3169 18388 9384 18452
rect 9448 18388 9468 18452
rect 3169 18372 9468 18388
rect 3169 18308 9384 18372
rect 9448 18308 9468 18372
rect 3169 18292 9468 18308
rect 3169 18228 9384 18292
rect 9448 18228 9468 18292
rect 3169 18212 9468 18228
rect 3169 18148 9384 18212
rect 9448 18148 9468 18212
rect 3169 18132 9468 18148
rect 3169 18068 9384 18132
rect 9448 18068 9468 18132
rect 3169 18052 9468 18068
rect 3169 17988 9384 18052
rect 9448 17988 9468 18052
rect 3169 17972 9468 17988
rect 3169 17908 9384 17972
rect 9448 17908 9468 17972
rect 3169 17892 9468 17908
rect 3169 17828 9384 17892
rect 9448 17828 9468 17892
rect 3169 17812 9468 17828
rect 3169 17748 9384 17812
rect 9448 17748 9468 17812
rect 3169 17732 9468 17748
rect 3169 17668 9384 17732
rect 9448 17668 9468 17732
rect 3169 17652 9468 17668
rect 3169 17588 9384 17652
rect 9448 17588 9468 17652
rect 3169 17572 9468 17588
rect 3169 17508 9384 17572
rect 9448 17508 9468 17572
rect 3169 17492 9468 17508
rect 3169 17428 9384 17492
rect 9448 17428 9468 17492
rect 3169 17412 9468 17428
rect 3169 17348 9384 17412
rect 9448 17348 9468 17412
rect 3169 17332 9468 17348
rect 3169 17268 9384 17332
rect 9448 17268 9468 17332
rect 3169 17252 9468 17268
rect 3169 17188 9384 17252
rect 9448 17188 9468 17252
rect 3169 17172 9468 17188
rect 3169 17108 9384 17172
rect 9448 17108 9468 17172
rect 3169 17092 9468 17108
rect 3169 17028 9384 17092
rect 9448 17028 9468 17092
rect 3169 17012 9468 17028
rect 3169 16948 9384 17012
rect 9448 16948 9468 17012
rect 3169 16932 9468 16948
rect 3169 16868 9384 16932
rect 9448 16868 9468 16932
rect 3169 16852 9468 16868
rect 3169 16788 9384 16852
rect 9448 16788 9468 16852
rect 3169 16772 9468 16788
rect 3169 16708 9384 16772
rect 9448 16708 9468 16772
rect 3169 16692 9468 16708
rect 3169 16628 9384 16692
rect 9448 16628 9468 16692
rect 3169 16612 9468 16628
rect 3169 16548 9384 16612
rect 9448 16548 9468 16612
rect 3169 16532 9468 16548
rect 3169 16468 9384 16532
rect 9448 16468 9468 16532
rect 3169 16452 9468 16468
rect 3169 16388 9384 16452
rect 9448 16388 9468 16452
rect 3169 16372 9468 16388
rect 3169 16308 9384 16372
rect 9448 16308 9468 16372
rect 3169 16292 9468 16308
rect 3169 16228 9384 16292
rect 9448 16228 9468 16292
rect 3169 16212 9468 16228
rect 3169 16148 9384 16212
rect 9448 16148 9468 16212
rect 3169 16132 9468 16148
rect 3169 16068 9384 16132
rect 9448 16068 9468 16132
rect 3169 16052 9468 16068
rect 3169 15988 9384 16052
rect 9448 15988 9468 16052
rect 3169 15972 9468 15988
rect 3169 15908 9384 15972
rect 9448 15908 9468 15972
rect 3169 15892 9468 15908
rect 3169 15828 9384 15892
rect 9448 15828 9468 15892
rect 3169 15800 9468 15828
rect 9488 21972 15787 22000
rect 9488 21908 15703 21972
rect 15767 21908 15787 21972
rect 9488 21892 15787 21908
rect 9488 21828 15703 21892
rect 15767 21828 15787 21892
rect 9488 21812 15787 21828
rect 9488 21748 15703 21812
rect 15767 21748 15787 21812
rect 9488 21732 15787 21748
rect 9488 21668 15703 21732
rect 15767 21668 15787 21732
rect 9488 21652 15787 21668
rect 9488 21588 15703 21652
rect 15767 21588 15787 21652
rect 9488 21572 15787 21588
rect 9488 21508 15703 21572
rect 15767 21508 15787 21572
rect 9488 21492 15787 21508
rect 9488 21428 15703 21492
rect 15767 21428 15787 21492
rect 9488 21412 15787 21428
rect 9488 21348 15703 21412
rect 15767 21348 15787 21412
rect 9488 21332 15787 21348
rect 9488 21268 15703 21332
rect 15767 21268 15787 21332
rect 9488 21252 15787 21268
rect 9488 21188 15703 21252
rect 15767 21188 15787 21252
rect 9488 21172 15787 21188
rect 9488 21108 15703 21172
rect 15767 21108 15787 21172
rect 9488 21092 15787 21108
rect 9488 21028 15703 21092
rect 15767 21028 15787 21092
rect 9488 21012 15787 21028
rect 9488 20948 15703 21012
rect 15767 20948 15787 21012
rect 9488 20932 15787 20948
rect 9488 20868 15703 20932
rect 15767 20868 15787 20932
rect 9488 20852 15787 20868
rect 9488 20788 15703 20852
rect 15767 20788 15787 20852
rect 9488 20772 15787 20788
rect 9488 20708 15703 20772
rect 15767 20708 15787 20772
rect 9488 20692 15787 20708
rect 9488 20628 15703 20692
rect 15767 20628 15787 20692
rect 9488 20612 15787 20628
rect 9488 20548 15703 20612
rect 15767 20548 15787 20612
rect 9488 20532 15787 20548
rect 9488 20468 15703 20532
rect 15767 20468 15787 20532
rect 9488 20452 15787 20468
rect 9488 20388 15703 20452
rect 15767 20388 15787 20452
rect 9488 20372 15787 20388
rect 9488 20308 15703 20372
rect 15767 20308 15787 20372
rect 9488 20292 15787 20308
rect 9488 20228 15703 20292
rect 15767 20228 15787 20292
rect 9488 20212 15787 20228
rect 9488 20148 15703 20212
rect 15767 20148 15787 20212
rect 9488 20132 15787 20148
rect 9488 20068 15703 20132
rect 15767 20068 15787 20132
rect 9488 20052 15787 20068
rect 9488 19988 15703 20052
rect 15767 19988 15787 20052
rect 9488 19972 15787 19988
rect 9488 19908 15703 19972
rect 15767 19908 15787 19972
rect 9488 19892 15787 19908
rect 9488 19828 15703 19892
rect 15767 19828 15787 19892
rect 9488 19812 15787 19828
rect 9488 19748 15703 19812
rect 15767 19748 15787 19812
rect 9488 19732 15787 19748
rect 9488 19668 15703 19732
rect 15767 19668 15787 19732
rect 9488 19652 15787 19668
rect 9488 19588 15703 19652
rect 15767 19588 15787 19652
rect 9488 19572 15787 19588
rect 9488 19508 15703 19572
rect 15767 19508 15787 19572
rect 9488 19492 15787 19508
rect 9488 19428 15703 19492
rect 15767 19428 15787 19492
rect 9488 19412 15787 19428
rect 9488 19348 15703 19412
rect 15767 19348 15787 19412
rect 9488 19332 15787 19348
rect 9488 19268 15703 19332
rect 15767 19268 15787 19332
rect 9488 19252 15787 19268
rect 9488 19188 15703 19252
rect 15767 19188 15787 19252
rect 9488 19172 15787 19188
rect 9488 19108 15703 19172
rect 15767 19108 15787 19172
rect 9488 19092 15787 19108
rect 9488 19028 15703 19092
rect 15767 19028 15787 19092
rect 9488 19012 15787 19028
rect 9488 18948 15703 19012
rect 15767 18948 15787 19012
rect 9488 18932 15787 18948
rect 9488 18868 15703 18932
rect 15767 18868 15787 18932
rect 9488 18852 15787 18868
rect 9488 18788 15703 18852
rect 15767 18788 15787 18852
rect 9488 18772 15787 18788
rect 9488 18708 15703 18772
rect 15767 18708 15787 18772
rect 9488 18692 15787 18708
rect 9488 18628 15703 18692
rect 15767 18628 15787 18692
rect 9488 18612 15787 18628
rect 9488 18548 15703 18612
rect 15767 18548 15787 18612
rect 9488 18532 15787 18548
rect 9488 18468 15703 18532
rect 15767 18468 15787 18532
rect 9488 18452 15787 18468
rect 9488 18388 15703 18452
rect 15767 18388 15787 18452
rect 9488 18372 15787 18388
rect 9488 18308 15703 18372
rect 15767 18308 15787 18372
rect 9488 18292 15787 18308
rect 9488 18228 15703 18292
rect 15767 18228 15787 18292
rect 9488 18212 15787 18228
rect 9488 18148 15703 18212
rect 15767 18148 15787 18212
rect 9488 18132 15787 18148
rect 9488 18068 15703 18132
rect 15767 18068 15787 18132
rect 9488 18052 15787 18068
rect 9488 17988 15703 18052
rect 15767 17988 15787 18052
rect 9488 17972 15787 17988
rect 9488 17908 15703 17972
rect 15767 17908 15787 17972
rect 9488 17892 15787 17908
rect 9488 17828 15703 17892
rect 15767 17828 15787 17892
rect 9488 17812 15787 17828
rect 9488 17748 15703 17812
rect 15767 17748 15787 17812
rect 9488 17732 15787 17748
rect 9488 17668 15703 17732
rect 15767 17668 15787 17732
rect 9488 17652 15787 17668
rect 9488 17588 15703 17652
rect 15767 17588 15787 17652
rect 9488 17572 15787 17588
rect 9488 17508 15703 17572
rect 15767 17508 15787 17572
rect 9488 17492 15787 17508
rect 9488 17428 15703 17492
rect 15767 17428 15787 17492
rect 9488 17412 15787 17428
rect 9488 17348 15703 17412
rect 15767 17348 15787 17412
rect 9488 17332 15787 17348
rect 9488 17268 15703 17332
rect 15767 17268 15787 17332
rect 9488 17252 15787 17268
rect 9488 17188 15703 17252
rect 15767 17188 15787 17252
rect 9488 17172 15787 17188
rect 9488 17108 15703 17172
rect 15767 17108 15787 17172
rect 9488 17092 15787 17108
rect 9488 17028 15703 17092
rect 15767 17028 15787 17092
rect 9488 17012 15787 17028
rect 9488 16948 15703 17012
rect 15767 16948 15787 17012
rect 9488 16932 15787 16948
rect 9488 16868 15703 16932
rect 15767 16868 15787 16932
rect 9488 16852 15787 16868
rect 9488 16788 15703 16852
rect 15767 16788 15787 16852
rect 9488 16772 15787 16788
rect 9488 16708 15703 16772
rect 15767 16708 15787 16772
rect 9488 16692 15787 16708
rect 9488 16628 15703 16692
rect 15767 16628 15787 16692
rect 9488 16612 15787 16628
rect 9488 16548 15703 16612
rect 15767 16548 15787 16612
rect 9488 16532 15787 16548
rect 9488 16468 15703 16532
rect 15767 16468 15787 16532
rect 9488 16452 15787 16468
rect 9488 16388 15703 16452
rect 15767 16388 15787 16452
rect 9488 16372 15787 16388
rect 9488 16308 15703 16372
rect 15767 16308 15787 16372
rect 9488 16292 15787 16308
rect 9488 16228 15703 16292
rect 15767 16228 15787 16292
rect 9488 16212 15787 16228
rect 9488 16148 15703 16212
rect 15767 16148 15787 16212
rect 9488 16132 15787 16148
rect 9488 16068 15703 16132
rect 15767 16068 15787 16132
rect 9488 16052 15787 16068
rect 9488 15988 15703 16052
rect 15767 15988 15787 16052
rect 9488 15972 15787 15988
rect 9488 15908 15703 15972
rect 15767 15908 15787 15972
rect 9488 15892 15787 15908
rect 9488 15828 15703 15892
rect 15767 15828 15787 15892
rect 9488 15800 15787 15828
rect 15807 21972 22106 22000
rect 15807 21908 22022 21972
rect 22086 21908 22106 21972
rect 15807 21892 22106 21908
rect 15807 21828 22022 21892
rect 22086 21828 22106 21892
rect 15807 21812 22106 21828
rect 15807 21748 22022 21812
rect 22086 21748 22106 21812
rect 15807 21732 22106 21748
rect 15807 21668 22022 21732
rect 22086 21668 22106 21732
rect 15807 21652 22106 21668
rect 15807 21588 22022 21652
rect 22086 21588 22106 21652
rect 15807 21572 22106 21588
rect 15807 21508 22022 21572
rect 22086 21508 22106 21572
rect 15807 21492 22106 21508
rect 15807 21428 22022 21492
rect 22086 21428 22106 21492
rect 15807 21412 22106 21428
rect 15807 21348 22022 21412
rect 22086 21348 22106 21412
rect 15807 21332 22106 21348
rect 15807 21268 22022 21332
rect 22086 21268 22106 21332
rect 15807 21252 22106 21268
rect 15807 21188 22022 21252
rect 22086 21188 22106 21252
rect 15807 21172 22106 21188
rect 15807 21108 22022 21172
rect 22086 21108 22106 21172
rect 15807 21092 22106 21108
rect 15807 21028 22022 21092
rect 22086 21028 22106 21092
rect 15807 21012 22106 21028
rect 15807 20948 22022 21012
rect 22086 20948 22106 21012
rect 15807 20932 22106 20948
rect 15807 20868 22022 20932
rect 22086 20868 22106 20932
rect 15807 20852 22106 20868
rect 15807 20788 22022 20852
rect 22086 20788 22106 20852
rect 15807 20772 22106 20788
rect 15807 20708 22022 20772
rect 22086 20708 22106 20772
rect 15807 20692 22106 20708
rect 15807 20628 22022 20692
rect 22086 20628 22106 20692
rect 15807 20612 22106 20628
rect 15807 20548 22022 20612
rect 22086 20548 22106 20612
rect 15807 20532 22106 20548
rect 15807 20468 22022 20532
rect 22086 20468 22106 20532
rect 15807 20452 22106 20468
rect 15807 20388 22022 20452
rect 22086 20388 22106 20452
rect 15807 20372 22106 20388
rect 15807 20308 22022 20372
rect 22086 20308 22106 20372
rect 15807 20292 22106 20308
rect 15807 20228 22022 20292
rect 22086 20228 22106 20292
rect 15807 20212 22106 20228
rect 15807 20148 22022 20212
rect 22086 20148 22106 20212
rect 15807 20132 22106 20148
rect 15807 20068 22022 20132
rect 22086 20068 22106 20132
rect 15807 20052 22106 20068
rect 15807 19988 22022 20052
rect 22086 19988 22106 20052
rect 15807 19972 22106 19988
rect 15807 19908 22022 19972
rect 22086 19908 22106 19972
rect 15807 19892 22106 19908
rect 15807 19828 22022 19892
rect 22086 19828 22106 19892
rect 15807 19812 22106 19828
rect 15807 19748 22022 19812
rect 22086 19748 22106 19812
rect 15807 19732 22106 19748
rect 15807 19668 22022 19732
rect 22086 19668 22106 19732
rect 15807 19652 22106 19668
rect 15807 19588 22022 19652
rect 22086 19588 22106 19652
rect 15807 19572 22106 19588
rect 15807 19508 22022 19572
rect 22086 19508 22106 19572
rect 15807 19492 22106 19508
rect 15807 19428 22022 19492
rect 22086 19428 22106 19492
rect 15807 19412 22106 19428
rect 15807 19348 22022 19412
rect 22086 19348 22106 19412
rect 15807 19332 22106 19348
rect 15807 19268 22022 19332
rect 22086 19268 22106 19332
rect 15807 19252 22106 19268
rect 15807 19188 22022 19252
rect 22086 19188 22106 19252
rect 15807 19172 22106 19188
rect 15807 19108 22022 19172
rect 22086 19108 22106 19172
rect 15807 19092 22106 19108
rect 15807 19028 22022 19092
rect 22086 19028 22106 19092
rect 15807 19012 22106 19028
rect 15807 18948 22022 19012
rect 22086 18948 22106 19012
rect 15807 18932 22106 18948
rect 15807 18868 22022 18932
rect 22086 18868 22106 18932
rect 15807 18852 22106 18868
rect 15807 18788 22022 18852
rect 22086 18788 22106 18852
rect 15807 18772 22106 18788
rect 15807 18708 22022 18772
rect 22086 18708 22106 18772
rect 15807 18692 22106 18708
rect 15807 18628 22022 18692
rect 22086 18628 22106 18692
rect 15807 18612 22106 18628
rect 15807 18548 22022 18612
rect 22086 18548 22106 18612
rect 15807 18532 22106 18548
rect 15807 18468 22022 18532
rect 22086 18468 22106 18532
rect 15807 18452 22106 18468
rect 15807 18388 22022 18452
rect 22086 18388 22106 18452
rect 15807 18372 22106 18388
rect 15807 18308 22022 18372
rect 22086 18308 22106 18372
rect 15807 18292 22106 18308
rect 15807 18228 22022 18292
rect 22086 18228 22106 18292
rect 15807 18212 22106 18228
rect 15807 18148 22022 18212
rect 22086 18148 22106 18212
rect 15807 18132 22106 18148
rect 15807 18068 22022 18132
rect 22086 18068 22106 18132
rect 15807 18052 22106 18068
rect 15807 17988 22022 18052
rect 22086 17988 22106 18052
rect 15807 17972 22106 17988
rect 15807 17908 22022 17972
rect 22086 17908 22106 17972
rect 15807 17892 22106 17908
rect 15807 17828 22022 17892
rect 22086 17828 22106 17892
rect 15807 17812 22106 17828
rect 15807 17748 22022 17812
rect 22086 17748 22106 17812
rect 15807 17732 22106 17748
rect 15807 17668 22022 17732
rect 22086 17668 22106 17732
rect 15807 17652 22106 17668
rect 15807 17588 22022 17652
rect 22086 17588 22106 17652
rect 15807 17572 22106 17588
rect 15807 17508 22022 17572
rect 22086 17508 22106 17572
rect 15807 17492 22106 17508
rect 15807 17428 22022 17492
rect 22086 17428 22106 17492
rect 15807 17412 22106 17428
rect 15807 17348 22022 17412
rect 22086 17348 22106 17412
rect 15807 17332 22106 17348
rect 15807 17268 22022 17332
rect 22086 17268 22106 17332
rect 15807 17252 22106 17268
rect 15807 17188 22022 17252
rect 22086 17188 22106 17252
rect 15807 17172 22106 17188
rect 15807 17108 22022 17172
rect 22086 17108 22106 17172
rect 15807 17092 22106 17108
rect 15807 17028 22022 17092
rect 22086 17028 22106 17092
rect 15807 17012 22106 17028
rect 15807 16948 22022 17012
rect 22086 16948 22106 17012
rect 15807 16932 22106 16948
rect 15807 16868 22022 16932
rect 22086 16868 22106 16932
rect 15807 16852 22106 16868
rect 15807 16788 22022 16852
rect 22086 16788 22106 16852
rect 15807 16772 22106 16788
rect 15807 16708 22022 16772
rect 22086 16708 22106 16772
rect 15807 16692 22106 16708
rect 15807 16628 22022 16692
rect 22086 16628 22106 16692
rect 15807 16612 22106 16628
rect 15807 16548 22022 16612
rect 22086 16548 22106 16612
rect 15807 16532 22106 16548
rect 15807 16468 22022 16532
rect 22086 16468 22106 16532
rect 15807 16452 22106 16468
rect 15807 16388 22022 16452
rect 22086 16388 22106 16452
rect 15807 16372 22106 16388
rect 15807 16308 22022 16372
rect 22086 16308 22106 16372
rect 15807 16292 22106 16308
rect 15807 16228 22022 16292
rect 22086 16228 22106 16292
rect 15807 16212 22106 16228
rect 15807 16148 22022 16212
rect 22086 16148 22106 16212
rect 15807 16132 22106 16148
rect 15807 16068 22022 16132
rect 22086 16068 22106 16132
rect 15807 16052 22106 16068
rect 15807 15988 22022 16052
rect 22086 15988 22106 16052
rect 15807 15972 22106 15988
rect 15807 15908 22022 15972
rect 22086 15908 22106 15972
rect 15807 15892 22106 15908
rect 15807 15828 22022 15892
rect 22086 15828 22106 15892
rect 15807 15800 22106 15828
rect 22126 21972 28425 22000
rect 22126 21908 28341 21972
rect 28405 21908 28425 21972
rect 22126 21892 28425 21908
rect 22126 21828 28341 21892
rect 28405 21828 28425 21892
rect 22126 21812 28425 21828
rect 22126 21748 28341 21812
rect 28405 21748 28425 21812
rect 22126 21732 28425 21748
rect 22126 21668 28341 21732
rect 28405 21668 28425 21732
rect 22126 21652 28425 21668
rect 22126 21588 28341 21652
rect 28405 21588 28425 21652
rect 22126 21572 28425 21588
rect 22126 21508 28341 21572
rect 28405 21508 28425 21572
rect 22126 21492 28425 21508
rect 22126 21428 28341 21492
rect 28405 21428 28425 21492
rect 22126 21412 28425 21428
rect 22126 21348 28341 21412
rect 28405 21348 28425 21412
rect 22126 21332 28425 21348
rect 22126 21268 28341 21332
rect 28405 21268 28425 21332
rect 22126 21252 28425 21268
rect 22126 21188 28341 21252
rect 28405 21188 28425 21252
rect 22126 21172 28425 21188
rect 22126 21108 28341 21172
rect 28405 21108 28425 21172
rect 22126 21092 28425 21108
rect 22126 21028 28341 21092
rect 28405 21028 28425 21092
rect 22126 21012 28425 21028
rect 22126 20948 28341 21012
rect 28405 20948 28425 21012
rect 22126 20932 28425 20948
rect 22126 20868 28341 20932
rect 28405 20868 28425 20932
rect 22126 20852 28425 20868
rect 22126 20788 28341 20852
rect 28405 20788 28425 20852
rect 22126 20772 28425 20788
rect 22126 20708 28341 20772
rect 28405 20708 28425 20772
rect 22126 20692 28425 20708
rect 22126 20628 28341 20692
rect 28405 20628 28425 20692
rect 22126 20612 28425 20628
rect 22126 20548 28341 20612
rect 28405 20548 28425 20612
rect 22126 20532 28425 20548
rect 22126 20468 28341 20532
rect 28405 20468 28425 20532
rect 22126 20452 28425 20468
rect 22126 20388 28341 20452
rect 28405 20388 28425 20452
rect 22126 20372 28425 20388
rect 22126 20308 28341 20372
rect 28405 20308 28425 20372
rect 22126 20292 28425 20308
rect 22126 20228 28341 20292
rect 28405 20228 28425 20292
rect 22126 20212 28425 20228
rect 22126 20148 28341 20212
rect 28405 20148 28425 20212
rect 22126 20132 28425 20148
rect 22126 20068 28341 20132
rect 28405 20068 28425 20132
rect 22126 20052 28425 20068
rect 22126 19988 28341 20052
rect 28405 19988 28425 20052
rect 22126 19972 28425 19988
rect 22126 19908 28341 19972
rect 28405 19908 28425 19972
rect 22126 19892 28425 19908
rect 22126 19828 28341 19892
rect 28405 19828 28425 19892
rect 22126 19812 28425 19828
rect 22126 19748 28341 19812
rect 28405 19748 28425 19812
rect 22126 19732 28425 19748
rect 22126 19668 28341 19732
rect 28405 19668 28425 19732
rect 22126 19652 28425 19668
rect 22126 19588 28341 19652
rect 28405 19588 28425 19652
rect 22126 19572 28425 19588
rect 22126 19508 28341 19572
rect 28405 19508 28425 19572
rect 22126 19492 28425 19508
rect 22126 19428 28341 19492
rect 28405 19428 28425 19492
rect 22126 19412 28425 19428
rect 22126 19348 28341 19412
rect 28405 19348 28425 19412
rect 22126 19332 28425 19348
rect 22126 19268 28341 19332
rect 28405 19268 28425 19332
rect 22126 19252 28425 19268
rect 22126 19188 28341 19252
rect 28405 19188 28425 19252
rect 22126 19172 28425 19188
rect 22126 19108 28341 19172
rect 28405 19108 28425 19172
rect 22126 19092 28425 19108
rect 22126 19028 28341 19092
rect 28405 19028 28425 19092
rect 22126 19012 28425 19028
rect 22126 18948 28341 19012
rect 28405 18948 28425 19012
rect 22126 18932 28425 18948
rect 22126 18868 28341 18932
rect 28405 18868 28425 18932
rect 22126 18852 28425 18868
rect 22126 18788 28341 18852
rect 28405 18788 28425 18852
rect 22126 18772 28425 18788
rect 22126 18708 28341 18772
rect 28405 18708 28425 18772
rect 22126 18692 28425 18708
rect 22126 18628 28341 18692
rect 28405 18628 28425 18692
rect 22126 18612 28425 18628
rect 22126 18548 28341 18612
rect 28405 18548 28425 18612
rect 22126 18532 28425 18548
rect 22126 18468 28341 18532
rect 28405 18468 28425 18532
rect 22126 18452 28425 18468
rect 22126 18388 28341 18452
rect 28405 18388 28425 18452
rect 22126 18372 28425 18388
rect 22126 18308 28341 18372
rect 28405 18308 28425 18372
rect 22126 18292 28425 18308
rect 22126 18228 28341 18292
rect 28405 18228 28425 18292
rect 22126 18212 28425 18228
rect 22126 18148 28341 18212
rect 28405 18148 28425 18212
rect 22126 18132 28425 18148
rect 22126 18068 28341 18132
rect 28405 18068 28425 18132
rect 22126 18052 28425 18068
rect 22126 17988 28341 18052
rect 28405 17988 28425 18052
rect 22126 17972 28425 17988
rect 22126 17908 28341 17972
rect 28405 17908 28425 17972
rect 22126 17892 28425 17908
rect 22126 17828 28341 17892
rect 28405 17828 28425 17892
rect 22126 17812 28425 17828
rect 22126 17748 28341 17812
rect 28405 17748 28425 17812
rect 22126 17732 28425 17748
rect 22126 17668 28341 17732
rect 28405 17668 28425 17732
rect 22126 17652 28425 17668
rect 22126 17588 28341 17652
rect 28405 17588 28425 17652
rect 22126 17572 28425 17588
rect 22126 17508 28341 17572
rect 28405 17508 28425 17572
rect 22126 17492 28425 17508
rect 22126 17428 28341 17492
rect 28405 17428 28425 17492
rect 22126 17412 28425 17428
rect 22126 17348 28341 17412
rect 28405 17348 28425 17412
rect 22126 17332 28425 17348
rect 22126 17268 28341 17332
rect 28405 17268 28425 17332
rect 22126 17252 28425 17268
rect 22126 17188 28341 17252
rect 28405 17188 28425 17252
rect 22126 17172 28425 17188
rect 22126 17108 28341 17172
rect 28405 17108 28425 17172
rect 22126 17092 28425 17108
rect 22126 17028 28341 17092
rect 28405 17028 28425 17092
rect 22126 17012 28425 17028
rect 22126 16948 28341 17012
rect 28405 16948 28425 17012
rect 22126 16932 28425 16948
rect 22126 16868 28341 16932
rect 28405 16868 28425 16932
rect 22126 16852 28425 16868
rect 22126 16788 28341 16852
rect 28405 16788 28425 16852
rect 22126 16772 28425 16788
rect 22126 16708 28341 16772
rect 28405 16708 28425 16772
rect 22126 16692 28425 16708
rect 22126 16628 28341 16692
rect 28405 16628 28425 16692
rect 22126 16612 28425 16628
rect 22126 16548 28341 16612
rect 28405 16548 28425 16612
rect 22126 16532 28425 16548
rect 22126 16468 28341 16532
rect 28405 16468 28425 16532
rect 22126 16452 28425 16468
rect 22126 16388 28341 16452
rect 28405 16388 28425 16452
rect 22126 16372 28425 16388
rect 22126 16308 28341 16372
rect 28405 16308 28425 16372
rect 22126 16292 28425 16308
rect 22126 16228 28341 16292
rect 28405 16228 28425 16292
rect 22126 16212 28425 16228
rect 22126 16148 28341 16212
rect 28405 16148 28425 16212
rect 22126 16132 28425 16148
rect 22126 16068 28341 16132
rect 28405 16068 28425 16132
rect 22126 16052 28425 16068
rect 22126 15988 28341 16052
rect 28405 15988 28425 16052
rect 22126 15972 28425 15988
rect 22126 15908 28341 15972
rect 28405 15908 28425 15972
rect 22126 15892 28425 15908
rect 22126 15828 28341 15892
rect 28405 15828 28425 15892
rect 22126 15800 28425 15828
rect 28445 21972 34744 22000
rect 28445 21908 34660 21972
rect 34724 21908 34744 21972
rect 28445 21892 34744 21908
rect 28445 21828 34660 21892
rect 34724 21828 34744 21892
rect 28445 21812 34744 21828
rect 28445 21748 34660 21812
rect 34724 21748 34744 21812
rect 28445 21732 34744 21748
rect 28445 21668 34660 21732
rect 34724 21668 34744 21732
rect 28445 21652 34744 21668
rect 28445 21588 34660 21652
rect 34724 21588 34744 21652
rect 28445 21572 34744 21588
rect 28445 21508 34660 21572
rect 34724 21508 34744 21572
rect 28445 21492 34744 21508
rect 28445 21428 34660 21492
rect 34724 21428 34744 21492
rect 28445 21412 34744 21428
rect 28445 21348 34660 21412
rect 34724 21348 34744 21412
rect 28445 21332 34744 21348
rect 28445 21268 34660 21332
rect 34724 21268 34744 21332
rect 28445 21252 34744 21268
rect 28445 21188 34660 21252
rect 34724 21188 34744 21252
rect 28445 21172 34744 21188
rect 28445 21108 34660 21172
rect 34724 21108 34744 21172
rect 28445 21092 34744 21108
rect 28445 21028 34660 21092
rect 34724 21028 34744 21092
rect 28445 21012 34744 21028
rect 28445 20948 34660 21012
rect 34724 20948 34744 21012
rect 28445 20932 34744 20948
rect 28445 20868 34660 20932
rect 34724 20868 34744 20932
rect 28445 20852 34744 20868
rect 28445 20788 34660 20852
rect 34724 20788 34744 20852
rect 28445 20772 34744 20788
rect 28445 20708 34660 20772
rect 34724 20708 34744 20772
rect 28445 20692 34744 20708
rect 28445 20628 34660 20692
rect 34724 20628 34744 20692
rect 28445 20612 34744 20628
rect 28445 20548 34660 20612
rect 34724 20548 34744 20612
rect 28445 20532 34744 20548
rect 28445 20468 34660 20532
rect 34724 20468 34744 20532
rect 28445 20452 34744 20468
rect 28445 20388 34660 20452
rect 34724 20388 34744 20452
rect 28445 20372 34744 20388
rect 28445 20308 34660 20372
rect 34724 20308 34744 20372
rect 28445 20292 34744 20308
rect 28445 20228 34660 20292
rect 34724 20228 34744 20292
rect 28445 20212 34744 20228
rect 28445 20148 34660 20212
rect 34724 20148 34744 20212
rect 28445 20132 34744 20148
rect 28445 20068 34660 20132
rect 34724 20068 34744 20132
rect 28445 20052 34744 20068
rect 28445 19988 34660 20052
rect 34724 19988 34744 20052
rect 28445 19972 34744 19988
rect 28445 19908 34660 19972
rect 34724 19908 34744 19972
rect 28445 19892 34744 19908
rect 28445 19828 34660 19892
rect 34724 19828 34744 19892
rect 28445 19812 34744 19828
rect 28445 19748 34660 19812
rect 34724 19748 34744 19812
rect 28445 19732 34744 19748
rect 28445 19668 34660 19732
rect 34724 19668 34744 19732
rect 28445 19652 34744 19668
rect 28445 19588 34660 19652
rect 34724 19588 34744 19652
rect 28445 19572 34744 19588
rect 28445 19508 34660 19572
rect 34724 19508 34744 19572
rect 28445 19492 34744 19508
rect 28445 19428 34660 19492
rect 34724 19428 34744 19492
rect 28445 19412 34744 19428
rect 28445 19348 34660 19412
rect 34724 19348 34744 19412
rect 28445 19332 34744 19348
rect 28445 19268 34660 19332
rect 34724 19268 34744 19332
rect 28445 19252 34744 19268
rect 28445 19188 34660 19252
rect 34724 19188 34744 19252
rect 28445 19172 34744 19188
rect 28445 19108 34660 19172
rect 34724 19108 34744 19172
rect 28445 19092 34744 19108
rect 28445 19028 34660 19092
rect 34724 19028 34744 19092
rect 28445 19012 34744 19028
rect 28445 18948 34660 19012
rect 34724 18948 34744 19012
rect 28445 18932 34744 18948
rect 28445 18868 34660 18932
rect 34724 18868 34744 18932
rect 28445 18852 34744 18868
rect 28445 18788 34660 18852
rect 34724 18788 34744 18852
rect 28445 18772 34744 18788
rect 28445 18708 34660 18772
rect 34724 18708 34744 18772
rect 28445 18692 34744 18708
rect 28445 18628 34660 18692
rect 34724 18628 34744 18692
rect 28445 18612 34744 18628
rect 28445 18548 34660 18612
rect 34724 18548 34744 18612
rect 28445 18532 34744 18548
rect 28445 18468 34660 18532
rect 34724 18468 34744 18532
rect 28445 18452 34744 18468
rect 28445 18388 34660 18452
rect 34724 18388 34744 18452
rect 28445 18372 34744 18388
rect 28445 18308 34660 18372
rect 34724 18308 34744 18372
rect 28445 18292 34744 18308
rect 28445 18228 34660 18292
rect 34724 18228 34744 18292
rect 28445 18212 34744 18228
rect 28445 18148 34660 18212
rect 34724 18148 34744 18212
rect 28445 18132 34744 18148
rect 28445 18068 34660 18132
rect 34724 18068 34744 18132
rect 28445 18052 34744 18068
rect 28445 17988 34660 18052
rect 34724 17988 34744 18052
rect 28445 17972 34744 17988
rect 28445 17908 34660 17972
rect 34724 17908 34744 17972
rect 28445 17892 34744 17908
rect 28445 17828 34660 17892
rect 34724 17828 34744 17892
rect 28445 17812 34744 17828
rect 28445 17748 34660 17812
rect 34724 17748 34744 17812
rect 28445 17732 34744 17748
rect 28445 17668 34660 17732
rect 34724 17668 34744 17732
rect 28445 17652 34744 17668
rect 28445 17588 34660 17652
rect 34724 17588 34744 17652
rect 28445 17572 34744 17588
rect 28445 17508 34660 17572
rect 34724 17508 34744 17572
rect 28445 17492 34744 17508
rect 28445 17428 34660 17492
rect 34724 17428 34744 17492
rect 28445 17412 34744 17428
rect 28445 17348 34660 17412
rect 34724 17348 34744 17412
rect 28445 17332 34744 17348
rect 28445 17268 34660 17332
rect 34724 17268 34744 17332
rect 28445 17252 34744 17268
rect 28445 17188 34660 17252
rect 34724 17188 34744 17252
rect 28445 17172 34744 17188
rect 28445 17108 34660 17172
rect 34724 17108 34744 17172
rect 28445 17092 34744 17108
rect 28445 17028 34660 17092
rect 34724 17028 34744 17092
rect 28445 17012 34744 17028
rect 28445 16948 34660 17012
rect 34724 16948 34744 17012
rect 28445 16932 34744 16948
rect 28445 16868 34660 16932
rect 34724 16868 34744 16932
rect 28445 16852 34744 16868
rect 28445 16788 34660 16852
rect 34724 16788 34744 16852
rect 28445 16772 34744 16788
rect 28445 16708 34660 16772
rect 34724 16708 34744 16772
rect 28445 16692 34744 16708
rect 28445 16628 34660 16692
rect 34724 16628 34744 16692
rect 28445 16612 34744 16628
rect 28445 16548 34660 16612
rect 34724 16548 34744 16612
rect 28445 16532 34744 16548
rect 28445 16468 34660 16532
rect 34724 16468 34744 16532
rect 28445 16452 34744 16468
rect 28445 16388 34660 16452
rect 34724 16388 34744 16452
rect 28445 16372 34744 16388
rect 28445 16308 34660 16372
rect 34724 16308 34744 16372
rect 28445 16292 34744 16308
rect 28445 16228 34660 16292
rect 34724 16228 34744 16292
rect 28445 16212 34744 16228
rect 28445 16148 34660 16212
rect 34724 16148 34744 16212
rect 28445 16132 34744 16148
rect 28445 16068 34660 16132
rect 34724 16068 34744 16132
rect 28445 16052 34744 16068
rect 28445 15988 34660 16052
rect 34724 15988 34744 16052
rect 28445 15972 34744 15988
rect 28445 15908 34660 15972
rect 34724 15908 34744 15972
rect 28445 15892 34744 15908
rect 28445 15828 34660 15892
rect 34724 15828 34744 15892
rect 28445 15800 34744 15828
rect 34764 21972 41063 22000
rect 34764 21908 40979 21972
rect 41043 21908 41063 21972
rect 34764 21892 41063 21908
rect 34764 21828 40979 21892
rect 41043 21828 41063 21892
rect 34764 21812 41063 21828
rect 34764 21748 40979 21812
rect 41043 21748 41063 21812
rect 34764 21732 41063 21748
rect 34764 21668 40979 21732
rect 41043 21668 41063 21732
rect 34764 21652 41063 21668
rect 34764 21588 40979 21652
rect 41043 21588 41063 21652
rect 34764 21572 41063 21588
rect 34764 21508 40979 21572
rect 41043 21508 41063 21572
rect 34764 21492 41063 21508
rect 34764 21428 40979 21492
rect 41043 21428 41063 21492
rect 34764 21412 41063 21428
rect 34764 21348 40979 21412
rect 41043 21348 41063 21412
rect 34764 21332 41063 21348
rect 34764 21268 40979 21332
rect 41043 21268 41063 21332
rect 34764 21252 41063 21268
rect 34764 21188 40979 21252
rect 41043 21188 41063 21252
rect 34764 21172 41063 21188
rect 34764 21108 40979 21172
rect 41043 21108 41063 21172
rect 34764 21092 41063 21108
rect 34764 21028 40979 21092
rect 41043 21028 41063 21092
rect 34764 21012 41063 21028
rect 34764 20948 40979 21012
rect 41043 20948 41063 21012
rect 34764 20932 41063 20948
rect 34764 20868 40979 20932
rect 41043 20868 41063 20932
rect 34764 20852 41063 20868
rect 34764 20788 40979 20852
rect 41043 20788 41063 20852
rect 34764 20772 41063 20788
rect 34764 20708 40979 20772
rect 41043 20708 41063 20772
rect 34764 20692 41063 20708
rect 34764 20628 40979 20692
rect 41043 20628 41063 20692
rect 34764 20612 41063 20628
rect 34764 20548 40979 20612
rect 41043 20548 41063 20612
rect 34764 20532 41063 20548
rect 34764 20468 40979 20532
rect 41043 20468 41063 20532
rect 34764 20452 41063 20468
rect 34764 20388 40979 20452
rect 41043 20388 41063 20452
rect 34764 20372 41063 20388
rect 34764 20308 40979 20372
rect 41043 20308 41063 20372
rect 34764 20292 41063 20308
rect 34764 20228 40979 20292
rect 41043 20228 41063 20292
rect 34764 20212 41063 20228
rect 34764 20148 40979 20212
rect 41043 20148 41063 20212
rect 34764 20132 41063 20148
rect 34764 20068 40979 20132
rect 41043 20068 41063 20132
rect 34764 20052 41063 20068
rect 34764 19988 40979 20052
rect 41043 19988 41063 20052
rect 34764 19972 41063 19988
rect 34764 19908 40979 19972
rect 41043 19908 41063 19972
rect 34764 19892 41063 19908
rect 34764 19828 40979 19892
rect 41043 19828 41063 19892
rect 34764 19812 41063 19828
rect 34764 19748 40979 19812
rect 41043 19748 41063 19812
rect 34764 19732 41063 19748
rect 34764 19668 40979 19732
rect 41043 19668 41063 19732
rect 34764 19652 41063 19668
rect 34764 19588 40979 19652
rect 41043 19588 41063 19652
rect 34764 19572 41063 19588
rect 34764 19508 40979 19572
rect 41043 19508 41063 19572
rect 34764 19492 41063 19508
rect 34764 19428 40979 19492
rect 41043 19428 41063 19492
rect 34764 19412 41063 19428
rect 34764 19348 40979 19412
rect 41043 19348 41063 19412
rect 34764 19332 41063 19348
rect 34764 19268 40979 19332
rect 41043 19268 41063 19332
rect 34764 19252 41063 19268
rect 34764 19188 40979 19252
rect 41043 19188 41063 19252
rect 34764 19172 41063 19188
rect 34764 19108 40979 19172
rect 41043 19108 41063 19172
rect 34764 19092 41063 19108
rect 34764 19028 40979 19092
rect 41043 19028 41063 19092
rect 34764 19012 41063 19028
rect 34764 18948 40979 19012
rect 41043 18948 41063 19012
rect 34764 18932 41063 18948
rect 34764 18868 40979 18932
rect 41043 18868 41063 18932
rect 34764 18852 41063 18868
rect 34764 18788 40979 18852
rect 41043 18788 41063 18852
rect 34764 18772 41063 18788
rect 34764 18708 40979 18772
rect 41043 18708 41063 18772
rect 34764 18692 41063 18708
rect 34764 18628 40979 18692
rect 41043 18628 41063 18692
rect 34764 18612 41063 18628
rect 34764 18548 40979 18612
rect 41043 18548 41063 18612
rect 34764 18532 41063 18548
rect 34764 18468 40979 18532
rect 41043 18468 41063 18532
rect 34764 18452 41063 18468
rect 34764 18388 40979 18452
rect 41043 18388 41063 18452
rect 34764 18372 41063 18388
rect 34764 18308 40979 18372
rect 41043 18308 41063 18372
rect 34764 18292 41063 18308
rect 34764 18228 40979 18292
rect 41043 18228 41063 18292
rect 34764 18212 41063 18228
rect 34764 18148 40979 18212
rect 41043 18148 41063 18212
rect 34764 18132 41063 18148
rect 34764 18068 40979 18132
rect 41043 18068 41063 18132
rect 34764 18052 41063 18068
rect 34764 17988 40979 18052
rect 41043 17988 41063 18052
rect 34764 17972 41063 17988
rect 34764 17908 40979 17972
rect 41043 17908 41063 17972
rect 34764 17892 41063 17908
rect 34764 17828 40979 17892
rect 41043 17828 41063 17892
rect 34764 17812 41063 17828
rect 34764 17748 40979 17812
rect 41043 17748 41063 17812
rect 34764 17732 41063 17748
rect 34764 17668 40979 17732
rect 41043 17668 41063 17732
rect 34764 17652 41063 17668
rect 34764 17588 40979 17652
rect 41043 17588 41063 17652
rect 34764 17572 41063 17588
rect 34764 17508 40979 17572
rect 41043 17508 41063 17572
rect 34764 17492 41063 17508
rect 34764 17428 40979 17492
rect 41043 17428 41063 17492
rect 34764 17412 41063 17428
rect 34764 17348 40979 17412
rect 41043 17348 41063 17412
rect 34764 17332 41063 17348
rect 34764 17268 40979 17332
rect 41043 17268 41063 17332
rect 34764 17252 41063 17268
rect 34764 17188 40979 17252
rect 41043 17188 41063 17252
rect 34764 17172 41063 17188
rect 34764 17108 40979 17172
rect 41043 17108 41063 17172
rect 34764 17092 41063 17108
rect 34764 17028 40979 17092
rect 41043 17028 41063 17092
rect 34764 17012 41063 17028
rect 34764 16948 40979 17012
rect 41043 16948 41063 17012
rect 34764 16932 41063 16948
rect 34764 16868 40979 16932
rect 41043 16868 41063 16932
rect 34764 16852 41063 16868
rect 34764 16788 40979 16852
rect 41043 16788 41063 16852
rect 34764 16772 41063 16788
rect 34764 16708 40979 16772
rect 41043 16708 41063 16772
rect 34764 16692 41063 16708
rect 34764 16628 40979 16692
rect 41043 16628 41063 16692
rect 34764 16612 41063 16628
rect 34764 16548 40979 16612
rect 41043 16548 41063 16612
rect 34764 16532 41063 16548
rect 34764 16468 40979 16532
rect 41043 16468 41063 16532
rect 34764 16452 41063 16468
rect 34764 16388 40979 16452
rect 41043 16388 41063 16452
rect 34764 16372 41063 16388
rect 34764 16308 40979 16372
rect 41043 16308 41063 16372
rect 34764 16292 41063 16308
rect 34764 16228 40979 16292
rect 41043 16228 41063 16292
rect 34764 16212 41063 16228
rect 34764 16148 40979 16212
rect 41043 16148 41063 16212
rect 34764 16132 41063 16148
rect 34764 16068 40979 16132
rect 41043 16068 41063 16132
rect 34764 16052 41063 16068
rect 34764 15988 40979 16052
rect 41043 15988 41063 16052
rect 34764 15972 41063 15988
rect 34764 15908 40979 15972
rect 41043 15908 41063 15972
rect 34764 15892 41063 15908
rect 34764 15828 40979 15892
rect 41043 15828 41063 15892
rect 34764 15800 41063 15828
rect 41083 21972 47382 22000
rect 41083 21908 47298 21972
rect 47362 21908 47382 21972
rect 41083 21892 47382 21908
rect 41083 21828 47298 21892
rect 47362 21828 47382 21892
rect 41083 21812 47382 21828
rect 41083 21748 47298 21812
rect 47362 21748 47382 21812
rect 41083 21732 47382 21748
rect 41083 21668 47298 21732
rect 47362 21668 47382 21732
rect 41083 21652 47382 21668
rect 41083 21588 47298 21652
rect 47362 21588 47382 21652
rect 41083 21572 47382 21588
rect 41083 21508 47298 21572
rect 47362 21508 47382 21572
rect 41083 21492 47382 21508
rect 41083 21428 47298 21492
rect 47362 21428 47382 21492
rect 41083 21412 47382 21428
rect 41083 21348 47298 21412
rect 47362 21348 47382 21412
rect 41083 21332 47382 21348
rect 41083 21268 47298 21332
rect 47362 21268 47382 21332
rect 41083 21252 47382 21268
rect 41083 21188 47298 21252
rect 47362 21188 47382 21252
rect 41083 21172 47382 21188
rect 41083 21108 47298 21172
rect 47362 21108 47382 21172
rect 41083 21092 47382 21108
rect 41083 21028 47298 21092
rect 47362 21028 47382 21092
rect 41083 21012 47382 21028
rect 41083 20948 47298 21012
rect 47362 20948 47382 21012
rect 41083 20932 47382 20948
rect 41083 20868 47298 20932
rect 47362 20868 47382 20932
rect 41083 20852 47382 20868
rect 41083 20788 47298 20852
rect 47362 20788 47382 20852
rect 41083 20772 47382 20788
rect 41083 20708 47298 20772
rect 47362 20708 47382 20772
rect 41083 20692 47382 20708
rect 41083 20628 47298 20692
rect 47362 20628 47382 20692
rect 41083 20612 47382 20628
rect 41083 20548 47298 20612
rect 47362 20548 47382 20612
rect 41083 20532 47382 20548
rect 41083 20468 47298 20532
rect 47362 20468 47382 20532
rect 41083 20452 47382 20468
rect 41083 20388 47298 20452
rect 47362 20388 47382 20452
rect 41083 20372 47382 20388
rect 41083 20308 47298 20372
rect 47362 20308 47382 20372
rect 41083 20292 47382 20308
rect 41083 20228 47298 20292
rect 47362 20228 47382 20292
rect 41083 20212 47382 20228
rect 41083 20148 47298 20212
rect 47362 20148 47382 20212
rect 41083 20132 47382 20148
rect 41083 20068 47298 20132
rect 47362 20068 47382 20132
rect 41083 20052 47382 20068
rect 41083 19988 47298 20052
rect 47362 19988 47382 20052
rect 41083 19972 47382 19988
rect 41083 19908 47298 19972
rect 47362 19908 47382 19972
rect 41083 19892 47382 19908
rect 41083 19828 47298 19892
rect 47362 19828 47382 19892
rect 41083 19812 47382 19828
rect 41083 19748 47298 19812
rect 47362 19748 47382 19812
rect 41083 19732 47382 19748
rect 41083 19668 47298 19732
rect 47362 19668 47382 19732
rect 41083 19652 47382 19668
rect 41083 19588 47298 19652
rect 47362 19588 47382 19652
rect 41083 19572 47382 19588
rect 41083 19508 47298 19572
rect 47362 19508 47382 19572
rect 41083 19492 47382 19508
rect 41083 19428 47298 19492
rect 47362 19428 47382 19492
rect 41083 19412 47382 19428
rect 41083 19348 47298 19412
rect 47362 19348 47382 19412
rect 41083 19332 47382 19348
rect 41083 19268 47298 19332
rect 47362 19268 47382 19332
rect 41083 19252 47382 19268
rect 41083 19188 47298 19252
rect 47362 19188 47382 19252
rect 41083 19172 47382 19188
rect 41083 19108 47298 19172
rect 47362 19108 47382 19172
rect 41083 19092 47382 19108
rect 41083 19028 47298 19092
rect 47362 19028 47382 19092
rect 41083 19012 47382 19028
rect 41083 18948 47298 19012
rect 47362 18948 47382 19012
rect 41083 18932 47382 18948
rect 41083 18868 47298 18932
rect 47362 18868 47382 18932
rect 41083 18852 47382 18868
rect 41083 18788 47298 18852
rect 47362 18788 47382 18852
rect 41083 18772 47382 18788
rect 41083 18708 47298 18772
rect 47362 18708 47382 18772
rect 41083 18692 47382 18708
rect 41083 18628 47298 18692
rect 47362 18628 47382 18692
rect 41083 18612 47382 18628
rect 41083 18548 47298 18612
rect 47362 18548 47382 18612
rect 41083 18532 47382 18548
rect 41083 18468 47298 18532
rect 47362 18468 47382 18532
rect 41083 18452 47382 18468
rect 41083 18388 47298 18452
rect 47362 18388 47382 18452
rect 41083 18372 47382 18388
rect 41083 18308 47298 18372
rect 47362 18308 47382 18372
rect 41083 18292 47382 18308
rect 41083 18228 47298 18292
rect 47362 18228 47382 18292
rect 41083 18212 47382 18228
rect 41083 18148 47298 18212
rect 47362 18148 47382 18212
rect 41083 18132 47382 18148
rect 41083 18068 47298 18132
rect 47362 18068 47382 18132
rect 41083 18052 47382 18068
rect 41083 17988 47298 18052
rect 47362 17988 47382 18052
rect 41083 17972 47382 17988
rect 41083 17908 47298 17972
rect 47362 17908 47382 17972
rect 41083 17892 47382 17908
rect 41083 17828 47298 17892
rect 47362 17828 47382 17892
rect 41083 17812 47382 17828
rect 41083 17748 47298 17812
rect 47362 17748 47382 17812
rect 41083 17732 47382 17748
rect 41083 17668 47298 17732
rect 47362 17668 47382 17732
rect 41083 17652 47382 17668
rect 41083 17588 47298 17652
rect 47362 17588 47382 17652
rect 41083 17572 47382 17588
rect 41083 17508 47298 17572
rect 47362 17508 47382 17572
rect 41083 17492 47382 17508
rect 41083 17428 47298 17492
rect 47362 17428 47382 17492
rect 41083 17412 47382 17428
rect 41083 17348 47298 17412
rect 47362 17348 47382 17412
rect 41083 17332 47382 17348
rect 41083 17268 47298 17332
rect 47362 17268 47382 17332
rect 41083 17252 47382 17268
rect 41083 17188 47298 17252
rect 47362 17188 47382 17252
rect 41083 17172 47382 17188
rect 41083 17108 47298 17172
rect 47362 17108 47382 17172
rect 41083 17092 47382 17108
rect 41083 17028 47298 17092
rect 47362 17028 47382 17092
rect 41083 17012 47382 17028
rect 41083 16948 47298 17012
rect 47362 16948 47382 17012
rect 41083 16932 47382 16948
rect 41083 16868 47298 16932
rect 47362 16868 47382 16932
rect 41083 16852 47382 16868
rect 41083 16788 47298 16852
rect 47362 16788 47382 16852
rect 41083 16772 47382 16788
rect 41083 16708 47298 16772
rect 47362 16708 47382 16772
rect 41083 16692 47382 16708
rect 41083 16628 47298 16692
rect 47362 16628 47382 16692
rect 41083 16612 47382 16628
rect 41083 16548 47298 16612
rect 47362 16548 47382 16612
rect 41083 16532 47382 16548
rect 41083 16468 47298 16532
rect 47362 16468 47382 16532
rect 41083 16452 47382 16468
rect 41083 16388 47298 16452
rect 47362 16388 47382 16452
rect 41083 16372 47382 16388
rect 41083 16308 47298 16372
rect 47362 16308 47382 16372
rect 41083 16292 47382 16308
rect 41083 16228 47298 16292
rect 47362 16228 47382 16292
rect 41083 16212 47382 16228
rect 41083 16148 47298 16212
rect 47362 16148 47382 16212
rect 41083 16132 47382 16148
rect 41083 16068 47298 16132
rect 47362 16068 47382 16132
rect 41083 16052 47382 16068
rect 41083 15988 47298 16052
rect 47362 15988 47382 16052
rect 41083 15972 47382 15988
rect 41083 15908 47298 15972
rect 47362 15908 47382 15972
rect 41083 15892 47382 15908
rect 41083 15828 47298 15892
rect 47362 15828 47382 15892
rect 41083 15800 47382 15828
rect -47383 15672 -41084 15700
rect -47383 15608 -41168 15672
rect -41104 15608 -41084 15672
rect -47383 15592 -41084 15608
rect -47383 15528 -41168 15592
rect -41104 15528 -41084 15592
rect -47383 15512 -41084 15528
rect -47383 15448 -41168 15512
rect -41104 15448 -41084 15512
rect -47383 15432 -41084 15448
rect -47383 15368 -41168 15432
rect -41104 15368 -41084 15432
rect -47383 15352 -41084 15368
rect -47383 15288 -41168 15352
rect -41104 15288 -41084 15352
rect -47383 15272 -41084 15288
rect -47383 15208 -41168 15272
rect -41104 15208 -41084 15272
rect -47383 15192 -41084 15208
rect -47383 15128 -41168 15192
rect -41104 15128 -41084 15192
rect -47383 15112 -41084 15128
rect -47383 15048 -41168 15112
rect -41104 15048 -41084 15112
rect -47383 15032 -41084 15048
rect -47383 14968 -41168 15032
rect -41104 14968 -41084 15032
rect -47383 14952 -41084 14968
rect -47383 14888 -41168 14952
rect -41104 14888 -41084 14952
rect -47383 14872 -41084 14888
rect -47383 14808 -41168 14872
rect -41104 14808 -41084 14872
rect -47383 14792 -41084 14808
rect -47383 14728 -41168 14792
rect -41104 14728 -41084 14792
rect -47383 14712 -41084 14728
rect -47383 14648 -41168 14712
rect -41104 14648 -41084 14712
rect -47383 14632 -41084 14648
rect -47383 14568 -41168 14632
rect -41104 14568 -41084 14632
rect -47383 14552 -41084 14568
rect -47383 14488 -41168 14552
rect -41104 14488 -41084 14552
rect -47383 14472 -41084 14488
rect -47383 14408 -41168 14472
rect -41104 14408 -41084 14472
rect -47383 14392 -41084 14408
rect -47383 14328 -41168 14392
rect -41104 14328 -41084 14392
rect -47383 14312 -41084 14328
rect -47383 14248 -41168 14312
rect -41104 14248 -41084 14312
rect -47383 14232 -41084 14248
rect -47383 14168 -41168 14232
rect -41104 14168 -41084 14232
rect -47383 14152 -41084 14168
rect -47383 14088 -41168 14152
rect -41104 14088 -41084 14152
rect -47383 14072 -41084 14088
rect -47383 14008 -41168 14072
rect -41104 14008 -41084 14072
rect -47383 13992 -41084 14008
rect -47383 13928 -41168 13992
rect -41104 13928 -41084 13992
rect -47383 13912 -41084 13928
rect -47383 13848 -41168 13912
rect -41104 13848 -41084 13912
rect -47383 13832 -41084 13848
rect -47383 13768 -41168 13832
rect -41104 13768 -41084 13832
rect -47383 13752 -41084 13768
rect -47383 13688 -41168 13752
rect -41104 13688 -41084 13752
rect -47383 13672 -41084 13688
rect -47383 13608 -41168 13672
rect -41104 13608 -41084 13672
rect -47383 13592 -41084 13608
rect -47383 13528 -41168 13592
rect -41104 13528 -41084 13592
rect -47383 13512 -41084 13528
rect -47383 13448 -41168 13512
rect -41104 13448 -41084 13512
rect -47383 13432 -41084 13448
rect -47383 13368 -41168 13432
rect -41104 13368 -41084 13432
rect -47383 13352 -41084 13368
rect -47383 13288 -41168 13352
rect -41104 13288 -41084 13352
rect -47383 13272 -41084 13288
rect -47383 13208 -41168 13272
rect -41104 13208 -41084 13272
rect -47383 13192 -41084 13208
rect -47383 13128 -41168 13192
rect -41104 13128 -41084 13192
rect -47383 13112 -41084 13128
rect -47383 13048 -41168 13112
rect -41104 13048 -41084 13112
rect -47383 13032 -41084 13048
rect -47383 12968 -41168 13032
rect -41104 12968 -41084 13032
rect -47383 12952 -41084 12968
rect -47383 12888 -41168 12952
rect -41104 12888 -41084 12952
rect -47383 12872 -41084 12888
rect -47383 12808 -41168 12872
rect -41104 12808 -41084 12872
rect -47383 12792 -41084 12808
rect -47383 12728 -41168 12792
rect -41104 12728 -41084 12792
rect -47383 12712 -41084 12728
rect -47383 12648 -41168 12712
rect -41104 12648 -41084 12712
rect -47383 12632 -41084 12648
rect -47383 12568 -41168 12632
rect -41104 12568 -41084 12632
rect -47383 12552 -41084 12568
rect -47383 12488 -41168 12552
rect -41104 12488 -41084 12552
rect -47383 12472 -41084 12488
rect -47383 12408 -41168 12472
rect -41104 12408 -41084 12472
rect -47383 12392 -41084 12408
rect -47383 12328 -41168 12392
rect -41104 12328 -41084 12392
rect -47383 12312 -41084 12328
rect -47383 12248 -41168 12312
rect -41104 12248 -41084 12312
rect -47383 12232 -41084 12248
rect -47383 12168 -41168 12232
rect -41104 12168 -41084 12232
rect -47383 12152 -41084 12168
rect -47383 12088 -41168 12152
rect -41104 12088 -41084 12152
rect -47383 12072 -41084 12088
rect -47383 12008 -41168 12072
rect -41104 12008 -41084 12072
rect -47383 11992 -41084 12008
rect -47383 11928 -41168 11992
rect -41104 11928 -41084 11992
rect -47383 11912 -41084 11928
rect -47383 11848 -41168 11912
rect -41104 11848 -41084 11912
rect -47383 11832 -41084 11848
rect -47383 11768 -41168 11832
rect -41104 11768 -41084 11832
rect -47383 11752 -41084 11768
rect -47383 11688 -41168 11752
rect -41104 11688 -41084 11752
rect -47383 11672 -41084 11688
rect -47383 11608 -41168 11672
rect -41104 11608 -41084 11672
rect -47383 11592 -41084 11608
rect -47383 11528 -41168 11592
rect -41104 11528 -41084 11592
rect -47383 11512 -41084 11528
rect -47383 11448 -41168 11512
rect -41104 11448 -41084 11512
rect -47383 11432 -41084 11448
rect -47383 11368 -41168 11432
rect -41104 11368 -41084 11432
rect -47383 11352 -41084 11368
rect -47383 11288 -41168 11352
rect -41104 11288 -41084 11352
rect -47383 11272 -41084 11288
rect -47383 11208 -41168 11272
rect -41104 11208 -41084 11272
rect -47383 11192 -41084 11208
rect -47383 11128 -41168 11192
rect -41104 11128 -41084 11192
rect -47383 11112 -41084 11128
rect -47383 11048 -41168 11112
rect -41104 11048 -41084 11112
rect -47383 11032 -41084 11048
rect -47383 10968 -41168 11032
rect -41104 10968 -41084 11032
rect -47383 10952 -41084 10968
rect -47383 10888 -41168 10952
rect -41104 10888 -41084 10952
rect -47383 10872 -41084 10888
rect -47383 10808 -41168 10872
rect -41104 10808 -41084 10872
rect -47383 10792 -41084 10808
rect -47383 10728 -41168 10792
rect -41104 10728 -41084 10792
rect -47383 10712 -41084 10728
rect -47383 10648 -41168 10712
rect -41104 10648 -41084 10712
rect -47383 10632 -41084 10648
rect -47383 10568 -41168 10632
rect -41104 10568 -41084 10632
rect -47383 10552 -41084 10568
rect -47383 10488 -41168 10552
rect -41104 10488 -41084 10552
rect -47383 10472 -41084 10488
rect -47383 10408 -41168 10472
rect -41104 10408 -41084 10472
rect -47383 10392 -41084 10408
rect -47383 10328 -41168 10392
rect -41104 10328 -41084 10392
rect -47383 10312 -41084 10328
rect -47383 10248 -41168 10312
rect -41104 10248 -41084 10312
rect -47383 10232 -41084 10248
rect -47383 10168 -41168 10232
rect -41104 10168 -41084 10232
rect -47383 10152 -41084 10168
rect -47383 10088 -41168 10152
rect -41104 10088 -41084 10152
rect -47383 10072 -41084 10088
rect -47383 10008 -41168 10072
rect -41104 10008 -41084 10072
rect -47383 9992 -41084 10008
rect -47383 9928 -41168 9992
rect -41104 9928 -41084 9992
rect -47383 9912 -41084 9928
rect -47383 9848 -41168 9912
rect -41104 9848 -41084 9912
rect -47383 9832 -41084 9848
rect -47383 9768 -41168 9832
rect -41104 9768 -41084 9832
rect -47383 9752 -41084 9768
rect -47383 9688 -41168 9752
rect -41104 9688 -41084 9752
rect -47383 9672 -41084 9688
rect -47383 9608 -41168 9672
rect -41104 9608 -41084 9672
rect -47383 9592 -41084 9608
rect -47383 9528 -41168 9592
rect -41104 9528 -41084 9592
rect -47383 9500 -41084 9528
rect -41064 15672 -34765 15700
rect -41064 15608 -34849 15672
rect -34785 15608 -34765 15672
rect -41064 15592 -34765 15608
rect -41064 15528 -34849 15592
rect -34785 15528 -34765 15592
rect -41064 15512 -34765 15528
rect -41064 15448 -34849 15512
rect -34785 15448 -34765 15512
rect -41064 15432 -34765 15448
rect -41064 15368 -34849 15432
rect -34785 15368 -34765 15432
rect -41064 15352 -34765 15368
rect -41064 15288 -34849 15352
rect -34785 15288 -34765 15352
rect -41064 15272 -34765 15288
rect -41064 15208 -34849 15272
rect -34785 15208 -34765 15272
rect -41064 15192 -34765 15208
rect -41064 15128 -34849 15192
rect -34785 15128 -34765 15192
rect -41064 15112 -34765 15128
rect -41064 15048 -34849 15112
rect -34785 15048 -34765 15112
rect -41064 15032 -34765 15048
rect -41064 14968 -34849 15032
rect -34785 14968 -34765 15032
rect -41064 14952 -34765 14968
rect -41064 14888 -34849 14952
rect -34785 14888 -34765 14952
rect -41064 14872 -34765 14888
rect -41064 14808 -34849 14872
rect -34785 14808 -34765 14872
rect -41064 14792 -34765 14808
rect -41064 14728 -34849 14792
rect -34785 14728 -34765 14792
rect -41064 14712 -34765 14728
rect -41064 14648 -34849 14712
rect -34785 14648 -34765 14712
rect -41064 14632 -34765 14648
rect -41064 14568 -34849 14632
rect -34785 14568 -34765 14632
rect -41064 14552 -34765 14568
rect -41064 14488 -34849 14552
rect -34785 14488 -34765 14552
rect -41064 14472 -34765 14488
rect -41064 14408 -34849 14472
rect -34785 14408 -34765 14472
rect -41064 14392 -34765 14408
rect -41064 14328 -34849 14392
rect -34785 14328 -34765 14392
rect -41064 14312 -34765 14328
rect -41064 14248 -34849 14312
rect -34785 14248 -34765 14312
rect -41064 14232 -34765 14248
rect -41064 14168 -34849 14232
rect -34785 14168 -34765 14232
rect -41064 14152 -34765 14168
rect -41064 14088 -34849 14152
rect -34785 14088 -34765 14152
rect -41064 14072 -34765 14088
rect -41064 14008 -34849 14072
rect -34785 14008 -34765 14072
rect -41064 13992 -34765 14008
rect -41064 13928 -34849 13992
rect -34785 13928 -34765 13992
rect -41064 13912 -34765 13928
rect -41064 13848 -34849 13912
rect -34785 13848 -34765 13912
rect -41064 13832 -34765 13848
rect -41064 13768 -34849 13832
rect -34785 13768 -34765 13832
rect -41064 13752 -34765 13768
rect -41064 13688 -34849 13752
rect -34785 13688 -34765 13752
rect -41064 13672 -34765 13688
rect -41064 13608 -34849 13672
rect -34785 13608 -34765 13672
rect -41064 13592 -34765 13608
rect -41064 13528 -34849 13592
rect -34785 13528 -34765 13592
rect -41064 13512 -34765 13528
rect -41064 13448 -34849 13512
rect -34785 13448 -34765 13512
rect -41064 13432 -34765 13448
rect -41064 13368 -34849 13432
rect -34785 13368 -34765 13432
rect -41064 13352 -34765 13368
rect -41064 13288 -34849 13352
rect -34785 13288 -34765 13352
rect -41064 13272 -34765 13288
rect -41064 13208 -34849 13272
rect -34785 13208 -34765 13272
rect -41064 13192 -34765 13208
rect -41064 13128 -34849 13192
rect -34785 13128 -34765 13192
rect -41064 13112 -34765 13128
rect -41064 13048 -34849 13112
rect -34785 13048 -34765 13112
rect -41064 13032 -34765 13048
rect -41064 12968 -34849 13032
rect -34785 12968 -34765 13032
rect -41064 12952 -34765 12968
rect -41064 12888 -34849 12952
rect -34785 12888 -34765 12952
rect -41064 12872 -34765 12888
rect -41064 12808 -34849 12872
rect -34785 12808 -34765 12872
rect -41064 12792 -34765 12808
rect -41064 12728 -34849 12792
rect -34785 12728 -34765 12792
rect -41064 12712 -34765 12728
rect -41064 12648 -34849 12712
rect -34785 12648 -34765 12712
rect -41064 12632 -34765 12648
rect -41064 12568 -34849 12632
rect -34785 12568 -34765 12632
rect -41064 12552 -34765 12568
rect -41064 12488 -34849 12552
rect -34785 12488 -34765 12552
rect -41064 12472 -34765 12488
rect -41064 12408 -34849 12472
rect -34785 12408 -34765 12472
rect -41064 12392 -34765 12408
rect -41064 12328 -34849 12392
rect -34785 12328 -34765 12392
rect -41064 12312 -34765 12328
rect -41064 12248 -34849 12312
rect -34785 12248 -34765 12312
rect -41064 12232 -34765 12248
rect -41064 12168 -34849 12232
rect -34785 12168 -34765 12232
rect -41064 12152 -34765 12168
rect -41064 12088 -34849 12152
rect -34785 12088 -34765 12152
rect -41064 12072 -34765 12088
rect -41064 12008 -34849 12072
rect -34785 12008 -34765 12072
rect -41064 11992 -34765 12008
rect -41064 11928 -34849 11992
rect -34785 11928 -34765 11992
rect -41064 11912 -34765 11928
rect -41064 11848 -34849 11912
rect -34785 11848 -34765 11912
rect -41064 11832 -34765 11848
rect -41064 11768 -34849 11832
rect -34785 11768 -34765 11832
rect -41064 11752 -34765 11768
rect -41064 11688 -34849 11752
rect -34785 11688 -34765 11752
rect -41064 11672 -34765 11688
rect -41064 11608 -34849 11672
rect -34785 11608 -34765 11672
rect -41064 11592 -34765 11608
rect -41064 11528 -34849 11592
rect -34785 11528 -34765 11592
rect -41064 11512 -34765 11528
rect -41064 11448 -34849 11512
rect -34785 11448 -34765 11512
rect -41064 11432 -34765 11448
rect -41064 11368 -34849 11432
rect -34785 11368 -34765 11432
rect -41064 11352 -34765 11368
rect -41064 11288 -34849 11352
rect -34785 11288 -34765 11352
rect -41064 11272 -34765 11288
rect -41064 11208 -34849 11272
rect -34785 11208 -34765 11272
rect -41064 11192 -34765 11208
rect -41064 11128 -34849 11192
rect -34785 11128 -34765 11192
rect -41064 11112 -34765 11128
rect -41064 11048 -34849 11112
rect -34785 11048 -34765 11112
rect -41064 11032 -34765 11048
rect -41064 10968 -34849 11032
rect -34785 10968 -34765 11032
rect -41064 10952 -34765 10968
rect -41064 10888 -34849 10952
rect -34785 10888 -34765 10952
rect -41064 10872 -34765 10888
rect -41064 10808 -34849 10872
rect -34785 10808 -34765 10872
rect -41064 10792 -34765 10808
rect -41064 10728 -34849 10792
rect -34785 10728 -34765 10792
rect -41064 10712 -34765 10728
rect -41064 10648 -34849 10712
rect -34785 10648 -34765 10712
rect -41064 10632 -34765 10648
rect -41064 10568 -34849 10632
rect -34785 10568 -34765 10632
rect -41064 10552 -34765 10568
rect -41064 10488 -34849 10552
rect -34785 10488 -34765 10552
rect -41064 10472 -34765 10488
rect -41064 10408 -34849 10472
rect -34785 10408 -34765 10472
rect -41064 10392 -34765 10408
rect -41064 10328 -34849 10392
rect -34785 10328 -34765 10392
rect -41064 10312 -34765 10328
rect -41064 10248 -34849 10312
rect -34785 10248 -34765 10312
rect -41064 10232 -34765 10248
rect -41064 10168 -34849 10232
rect -34785 10168 -34765 10232
rect -41064 10152 -34765 10168
rect -41064 10088 -34849 10152
rect -34785 10088 -34765 10152
rect -41064 10072 -34765 10088
rect -41064 10008 -34849 10072
rect -34785 10008 -34765 10072
rect -41064 9992 -34765 10008
rect -41064 9928 -34849 9992
rect -34785 9928 -34765 9992
rect -41064 9912 -34765 9928
rect -41064 9848 -34849 9912
rect -34785 9848 -34765 9912
rect -41064 9832 -34765 9848
rect -41064 9768 -34849 9832
rect -34785 9768 -34765 9832
rect -41064 9752 -34765 9768
rect -41064 9688 -34849 9752
rect -34785 9688 -34765 9752
rect -41064 9672 -34765 9688
rect -41064 9608 -34849 9672
rect -34785 9608 -34765 9672
rect -41064 9592 -34765 9608
rect -41064 9528 -34849 9592
rect -34785 9528 -34765 9592
rect -41064 9500 -34765 9528
rect -34745 15672 -28446 15700
rect -34745 15608 -28530 15672
rect -28466 15608 -28446 15672
rect -34745 15592 -28446 15608
rect -34745 15528 -28530 15592
rect -28466 15528 -28446 15592
rect -34745 15512 -28446 15528
rect -34745 15448 -28530 15512
rect -28466 15448 -28446 15512
rect -34745 15432 -28446 15448
rect -34745 15368 -28530 15432
rect -28466 15368 -28446 15432
rect -34745 15352 -28446 15368
rect -34745 15288 -28530 15352
rect -28466 15288 -28446 15352
rect -34745 15272 -28446 15288
rect -34745 15208 -28530 15272
rect -28466 15208 -28446 15272
rect -34745 15192 -28446 15208
rect -34745 15128 -28530 15192
rect -28466 15128 -28446 15192
rect -34745 15112 -28446 15128
rect -34745 15048 -28530 15112
rect -28466 15048 -28446 15112
rect -34745 15032 -28446 15048
rect -34745 14968 -28530 15032
rect -28466 14968 -28446 15032
rect -34745 14952 -28446 14968
rect -34745 14888 -28530 14952
rect -28466 14888 -28446 14952
rect -34745 14872 -28446 14888
rect -34745 14808 -28530 14872
rect -28466 14808 -28446 14872
rect -34745 14792 -28446 14808
rect -34745 14728 -28530 14792
rect -28466 14728 -28446 14792
rect -34745 14712 -28446 14728
rect -34745 14648 -28530 14712
rect -28466 14648 -28446 14712
rect -34745 14632 -28446 14648
rect -34745 14568 -28530 14632
rect -28466 14568 -28446 14632
rect -34745 14552 -28446 14568
rect -34745 14488 -28530 14552
rect -28466 14488 -28446 14552
rect -34745 14472 -28446 14488
rect -34745 14408 -28530 14472
rect -28466 14408 -28446 14472
rect -34745 14392 -28446 14408
rect -34745 14328 -28530 14392
rect -28466 14328 -28446 14392
rect -34745 14312 -28446 14328
rect -34745 14248 -28530 14312
rect -28466 14248 -28446 14312
rect -34745 14232 -28446 14248
rect -34745 14168 -28530 14232
rect -28466 14168 -28446 14232
rect -34745 14152 -28446 14168
rect -34745 14088 -28530 14152
rect -28466 14088 -28446 14152
rect -34745 14072 -28446 14088
rect -34745 14008 -28530 14072
rect -28466 14008 -28446 14072
rect -34745 13992 -28446 14008
rect -34745 13928 -28530 13992
rect -28466 13928 -28446 13992
rect -34745 13912 -28446 13928
rect -34745 13848 -28530 13912
rect -28466 13848 -28446 13912
rect -34745 13832 -28446 13848
rect -34745 13768 -28530 13832
rect -28466 13768 -28446 13832
rect -34745 13752 -28446 13768
rect -34745 13688 -28530 13752
rect -28466 13688 -28446 13752
rect -34745 13672 -28446 13688
rect -34745 13608 -28530 13672
rect -28466 13608 -28446 13672
rect -34745 13592 -28446 13608
rect -34745 13528 -28530 13592
rect -28466 13528 -28446 13592
rect -34745 13512 -28446 13528
rect -34745 13448 -28530 13512
rect -28466 13448 -28446 13512
rect -34745 13432 -28446 13448
rect -34745 13368 -28530 13432
rect -28466 13368 -28446 13432
rect -34745 13352 -28446 13368
rect -34745 13288 -28530 13352
rect -28466 13288 -28446 13352
rect -34745 13272 -28446 13288
rect -34745 13208 -28530 13272
rect -28466 13208 -28446 13272
rect -34745 13192 -28446 13208
rect -34745 13128 -28530 13192
rect -28466 13128 -28446 13192
rect -34745 13112 -28446 13128
rect -34745 13048 -28530 13112
rect -28466 13048 -28446 13112
rect -34745 13032 -28446 13048
rect -34745 12968 -28530 13032
rect -28466 12968 -28446 13032
rect -34745 12952 -28446 12968
rect -34745 12888 -28530 12952
rect -28466 12888 -28446 12952
rect -34745 12872 -28446 12888
rect -34745 12808 -28530 12872
rect -28466 12808 -28446 12872
rect -34745 12792 -28446 12808
rect -34745 12728 -28530 12792
rect -28466 12728 -28446 12792
rect -34745 12712 -28446 12728
rect -34745 12648 -28530 12712
rect -28466 12648 -28446 12712
rect -34745 12632 -28446 12648
rect -34745 12568 -28530 12632
rect -28466 12568 -28446 12632
rect -34745 12552 -28446 12568
rect -34745 12488 -28530 12552
rect -28466 12488 -28446 12552
rect -34745 12472 -28446 12488
rect -34745 12408 -28530 12472
rect -28466 12408 -28446 12472
rect -34745 12392 -28446 12408
rect -34745 12328 -28530 12392
rect -28466 12328 -28446 12392
rect -34745 12312 -28446 12328
rect -34745 12248 -28530 12312
rect -28466 12248 -28446 12312
rect -34745 12232 -28446 12248
rect -34745 12168 -28530 12232
rect -28466 12168 -28446 12232
rect -34745 12152 -28446 12168
rect -34745 12088 -28530 12152
rect -28466 12088 -28446 12152
rect -34745 12072 -28446 12088
rect -34745 12008 -28530 12072
rect -28466 12008 -28446 12072
rect -34745 11992 -28446 12008
rect -34745 11928 -28530 11992
rect -28466 11928 -28446 11992
rect -34745 11912 -28446 11928
rect -34745 11848 -28530 11912
rect -28466 11848 -28446 11912
rect -34745 11832 -28446 11848
rect -34745 11768 -28530 11832
rect -28466 11768 -28446 11832
rect -34745 11752 -28446 11768
rect -34745 11688 -28530 11752
rect -28466 11688 -28446 11752
rect -34745 11672 -28446 11688
rect -34745 11608 -28530 11672
rect -28466 11608 -28446 11672
rect -34745 11592 -28446 11608
rect -34745 11528 -28530 11592
rect -28466 11528 -28446 11592
rect -34745 11512 -28446 11528
rect -34745 11448 -28530 11512
rect -28466 11448 -28446 11512
rect -34745 11432 -28446 11448
rect -34745 11368 -28530 11432
rect -28466 11368 -28446 11432
rect -34745 11352 -28446 11368
rect -34745 11288 -28530 11352
rect -28466 11288 -28446 11352
rect -34745 11272 -28446 11288
rect -34745 11208 -28530 11272
rect -28466 11208 -28446 11272
rect -34745 11192 -28446 11208
rect -34745 11128 -28530 11192
rect -28466 11128 -28446 11192
rect -34745 11112 -28446 11128
rect -34745 11048 -28530 11112
rect -28466 11048 -28446 11112
rect -34745 11032 -28446 11048
rect -34745 10968 -28530 11032
rect -28466 10968 -28446 11032
rect -34745 10952 -28446 10968
rect -34745 10888 -28530 10952
rect -28466 10888 -28446 10952
rect -34745 10872 -28446 10888
rect -34745 10808 -28530 10872
rect -28466 10808 -28446 10872
rect -34745 10792 -28446 10808
rect -34745 10728 -28530 10792
rect -28466 10728 -28446 10792
rect -34745 10712 -28446 10728
rect -34745 10648 -28530 10712
rect -28466 10648 -28446 10712
rect -34745 10632 -28446 10648
rect -34745 10568 -28530 10632
rect -28466 10568 -28446 10632
rect -34745 10552 -28446 10568
rect -34745 10488 -28530 10552
rect -28466 10488 -28446 10552
rect -34745 10472 -28446 10488
rect -34745 10408 -28530 10472
rect -28466 10408 -28446 10472
rect -34745 10392 -28446 10408
rect -34745 10328 -28530 10392
rect -28466 10328 -28446 10392
rect -34745 10312 -28446 10328
rect -34745 10248 -28530 10312
rect -28466 10248 -28446 10312
rect -34745 10232 -28446 10248
rect -34745 10168 -28530 10232
rect -28466 10168 -28446 10232
rect -34745 10152 -28446 10168
rect -34745 10088 -28530 10152
rect -28466 10088 -28446 10152
rect -34745 10072 -28446 10088
rect -34745 10008 -28530 10072
rect -28466 10008 -28446 10072
rect -34745 9992 -28446 10008
rect -34745 9928 -28530 9992
rect -28466 9928 -28446 9992
rect -34745 9912 -28446 9928
rect -34745 9848 -28530 9912
rect -28466 9848 -28446 9912
rect -34745 9832 -28446 9848
rect -34745 9768 -28530 9832
rect -28466 9768 -28446 9832
rect -34745 9752 -28446 9768
rect -34745 9688 -28530 9752
rect -28466 9688 -28446 9752
rect -34745 9672 -28446 9688
rect -34745 9608 -28530 9672
rect -28466 9608 -28446 9672
rect -34745 9592 -28446 9608
rect -34745 9528 -28530 9592
rect -28466 9528 -28446 9592
rect -34745 9500 -28446 9528
rect -28426 15672 -22127 15700
rect -28426 15608 -22211 15672
rect -22147 15608 -22127 15672
rect -28426 15592 -22127 15608
rect -28426 15528 -22211 15592
rect -22147 15528 -22127 15592
rect -28426 15512 -22127 15528
rect -28426 15448 -22211 15512
rect -22147 15448 -22127 15512
rect -28426 15432 -22127 15448
rect -28426 15368 -22211 15432
rect -22147 15368 -22127 15432
rect -28426 15352 -22127 15368
rect -28426 15288 -22211 15352
rect -22147 15288 -22127 15352
rect -28426 15272 -22127 15288
rect -28426 15208 -22211 15272
rect -22147 15208 -22127 15272
rect -28426 15192 -22127 15208
rect -28426 15128 -22211 15192
rect -22147 15128 -22127 15192
rect -28426 15112 -22127 15128
rect -28426 15048 -22211 15112
rect -22147 15048 -22127 15112
rect -28426 15032 -22127 15048
rect -28426 14968 -22211 15032
rect -22147 14968 -22127 15032
rect -28426 14952 -22127 14968
rect -28426 14888 -22211 14952
rect -22147 14888 -22127 14952
rect -28426 14872 -22127 14888
rect -28426 14808 -22211 14872
rect -22147 14808 -22127 14872
rect -28426 14792 -22127 14808
rect -28426 14728 -22211 14792
rect -22147 14728 -22127 14792
rect -28426 14712 -22127 14728
rect -28426 14648 -22211 14712
rect -22147 14648 -22127 14712
rect -28426 14632 -22127 14648
rect -28426 14568 -22211 14632
rect -22147 14568 -22127 14632
rect -28426 14552 -22127 14568
rect -28426 14488 -22211 14552
rect -22147 14488 -22127 14552
rect -28426 14472 -22127 14488
rect -28426 14408 -22211 14472
rect -22147 14408 -22127 14472
rect -28426 14392 -22127 14408
rect -28426 14328 -22211 14392
rect -22147 14328 -22127 14392
rect -28426 14312 -22127 14328
rect -28426 14248 -22211 14312
rect -22147 14248 -22127 14312
rect -28426 14232 -22127 14248
rect -28426 14168 -22211 14232
rect -22147 14168 -22127 14232
rect -28426 14152 -22127 14168
rect -28426 14088 -22211 14152
rect -22147 14088 -22127 14152
rect -28426 14072 -22127 14088
rect -28426 14008 -22211 14072
rect -22147 14008 -22127 14072
rect -28426 13992 -22127 14008
rect -28426 13928 -22211 13992
rect -22147 13928 -22127 13992
rect -28426 13912 -22127 13928
rect -28426 13848 -22211 13912
rect -22147 13848 -22127 13912
rect -28426 13832 -22127 13848
rect -28426 13768 -22211 13832
rect -22147 13768 -22127 13832
rect -28426 13752 -22127 13768
rect -28426 13688 -22211 13752
rect -22147 13688 -22127 13752
rect -28426 13672 -22127 13688
rect -28426 13608 -22211 13672
rect -22147 13608 -22127 13672
rect -28426 13592 -22127 13608
rect -28426 13528 -22211 13592
rect -22147 13528 -22127 13592
rect -28426 13512 -22127 13528
rect -28426 13448 -22211 13512
rect -22147 13448 -22127 13512
rect -28426 13432 -22127 13448
rect -28426 13368 -22211 13432
rect -22147 13368 -22127 13432
rect -28426 13352 -22127 13368
rect -28426 13288 -22211 13352
rect -22147 13288 -22127 13352
rect -28426 13272 -22127 13288
rect -28426 13208 -22211 13272
rect -22147 13208 -22127 13272
rect -28426 13192 -22127 13208
rect -28426 13128 -22211 13192
rect -22147 13128 -22127 13192
rect -28426 13112 -22127 13128
rect -28426 13048 -22211 13112
rect -22147 13048 -22127 13112
rect -28426 13032 -22127 13048
rect -28426 12968 -22211 13032
rect -22147 12968 -22127 13032
rect -28426 12952 -22127 12968
rect -28426 12888 -22211 12952
rect -22147 12888 -22127 12952
rect -28426 12872 -22127 12888
rect -28426 12808 -22211 12872
rect -22147 12808 -22127 12872
rect -28426 12792 -22127 12808
rect -28426 12728 -22211 12792
rect -22147 12728 -22127 12792
rect -28426 12712 -22127 12728
rect -28426 12648 -22211 12712
rect -22147 12648 -22127 12712
rect -28426 12632 -22127 12648
rect -28426 12568 -22211 12632
rect -22147 12568 -22127 12632
rect -28426 12552 -22127 12568
rect -28426 12488 -22211 12552
rect -22147 12488 -22127 12552
rect -28426 12472 -22127 12488
rect -28426 12408 -22211 12472
rect -22147 12408 -22127 12472
rect -28426 12392 -22127 12408
rect -28426 12328 -22211 12392
rect -22147 12328 -22127 12392
rect -28426 12312 -22127 12328
rect -28426 12248 -22211 12312
rect -22147 12248 -22127 12312
rect -28426 12232 -22127 12248
rect -28426 12168 -22211 12232
rect -22147 12168 -22127 12232
rect -28426 12152 -22127 12168
rect -28426 12088 -22211 12152
rect -22147 12088 -22127 12152
rect -28426 12072 -22127 12088
rect -28426 12008 -22211 12072
rect -22147 12008 -22127 12072
rect -28426 11992 -22127 12008
rect -28426 11928 -22211 11992
rect -22147 11928 -22127 11992
rect -28426 11912 -22127 11928
rect -28426 11848 -22211 11912
rect -22147 11848 -22127 11912
rect -28426 11832 -22127 11848
rect -28426 11768 -22211 11832
rect -22147 11768 -22127 11832
rect -28426 11752 -22127 11768
rect -28426 11688 -22211 11752
rect -22147 11688 -22127 11752
rect -28426 11672 -22127 11688
rect -28426 11608 -22211 11672
rect -22147 11608 -22127 11672
rect -28426 11592 -22127 11608
rect -28426 11528 -22211 11592
rect -22147 11528 -22127 11592
rect -28426 11512 -22127 11528
rect -28426 11448 -22211 11512
rect -22147 11448 -22127 11512
rect -28426 11432 -22127 11448
rect -28426 11368 -22211 11432
rect -22147 11368 -22127 11432
rect -28426 11352 -22127 11368
rect -28426 11288 -22211 11352
rect -22147 11288 -22127 11352
rect -28426 11272 -22127 11288
rect -28426 11208 -22211 11272
rect -22147 11208 -22127 11272
rect -28426 11192 -22127 11208
rect -28426 11128 -22211 11192
rect -22147 11128 -22127 11192
rect -28426 11112 -22127 11128
rect -28426 11048 -22211 11112
rect -22147 11048 -22127 11112
rect -28426 11032 -22127 11048
rect -28426 10968 -22211 11032
rect -22147 10968 -22127 11032
rect -28426 10952 -22127 10968
rect -28426 10888 -22211 10952
rect -22147 10888 -22127 10952
rect -28426 10872 -22127 10888
rect -28426 10808 -22211 10872
rect -22147 10808 -22127 10872
rect -28426 10792 -22127 10808
rect -28426 10728 -22211 10792
rect -22147 10728 -22127 10792
rect -28426 10712 -22127 10728
rect -28426 10648 -22211 10712
rect -22147 10648 -22127 10712
rect -28426 10632 -22127 10648
rect -28426 10568 -22211 10632
rect -22147 10568 -22127 10632
rect -28426 10552 -22127 10568
rect -28426 10488 -22211 10552
rect -22147 10488 -22127 10552
rect -28426 10472 -22127 10488
rect -28426 10408 -22211 10472
rect -22147 10408 -22127 10472
rect -28426 10392 -22127 10408
rect -28426 10328 -22211 10392
rect -22147 10328 -22127 10392
rect -28426 10312 -22127 10328
rect -28426 10248 -22211 10312
rect -22147 10248 -22127 10312
rect -28426 10232 -22127 10248
rect -28426 10168 -22211 10232
rect -22147 10168 -22127 10232
rect -28426 10152 -22127 10168
rect -28426 10088 -22211 10152
rect -22147 10088 -22127 10152
rect -28426 10072 -22127 10088
rect -28426 10008 -22211 10072
rect -22147 10008 -22127 10072
rect -28426 9992 -22127 10008
rect -28426 9928 -22211 9992
rect -22147 9928 -22127 9992
rect -28426 9912 -22127 9928
rect -28426 9848 -22211 9912
rect -22147 9848 -22127 9912
rect -28426 9832 -22127 9848
rect -28426 9768 -22211 9832
rect -22147 9768 -22127 9832
rect -28426 9752 -22127 9768
rect -28426 9688 -22211 9752
rect -22147 9688 -22127 9752
rect -28426 9672 -22127 9688
rect -28426 9608 -22211 9672
rect -22147 9608 -22127 9672
rect -28426 9592 -22127 9608
rect -28426 9528 -22211 9592
rect -22147 9528 -22127 9592
rect -28426 9500 -22127 9528
rect -22107 15672 -15808 15700
rect -22107 15608 -15892 15672
rect -15828 15608 -15808 15672
rect -22107 15592 -15808 15608
rect -22107 15528 -15892 15592
rect -15828 15528 -15808 15592
rect -22107 15512 -15808 15528
rect -22107 15448 -15892 15512
rect -15828 15448 -15808 15512
rect -22107 15432 -15808 15448
rect -22107 15368 -15892 15432
rect -15828 15368 -15808 15432
rect -22107 15352 -15808 15368
rect -22107 15288 -15892 15352
rect -15828 15288 -15808 15352
rect -22107 15272 -15808 15288
rect -22107 15208 -15892 15272
rect -15828 15208 -15808 15272
rect -22107 15192 -15808 15208
rect -22107 15128 -15892 15192
rect -15828 15128 -15808 15192
rect -22107 15112 -15808 15128
rect -22107 15048 -15892 15112
rect -15828 15048 -15808 15112
rect -22107 15032 -15808 15048
rect -22107 14968 -15892 15032
rect -15828 14968 -15808 15032
rect -22107 14952 -15808 14968
rect -22107 14888 -15892 14952
rect -15828 14888 -15808 14952
rect -22107 14872 -15808 14888
rect -22107 14808 -15892 14872
rect -15828 14808 -15808 14872
rect -22107 14792 -15808 14808
rect -22107 14728 -15892 14792
rect -15828 14728 -15808 14792
rect -22107 14712 -15808 14728
rect -22107 14648 -15892 14712
rect -15828 14648 -15808 14712
rect -22107 14632 -15808 14648
rect -22107 14568 -15892 14632
rect -15828 14568 -15808 14632
rect -22107 14552 -15808 14568
rect -22107 14488 -15892 14552
rect -15828 14488 -15808 14552
rect -22107 14472 -15808 14488
rect -22107 14408 -15892 14472
rect -15828 14408 -15808 14472
rect -22107 14392 -15808 14408
rect -22107 14328 -15892 14392
rect -15828 14328 -15808 14392
rect -22107 14312 -15808 14328
rect -22107 14248 -15892 14312
rect -15828 14248 -15808 14312
rect -22107 14232 -15808 14248
rect -22107 14168 -15892 14232
rect -15828 14168 -15808 14232
rect -22107 14152 -15808 14168
rect -22107 14088 -15892 14152
rect -15828 14088 -15808 14152
rect -22107 14072 -15808 14088
rect -22107 14008 -15892 14072
rect -15828 14008 -15808 14072
rect -22107 13992 -15808 14008
rect -22107 13928 -15892 13992
rect -15828 13928 -15808 13992
rect -22107 13912 -15808 13928
rect -22107 13848 -15892 13912
rect -15828 13848 -15808 13912
rect -22107 13832 -15808 13848
rect -22107 13768 -15892 13832
rect -15828 13768 -15808 13832
rect -22107 13752 -15808 13768
rect -22107 13688 -15892 13752
rect -15828 13688 -15808 13752
rect -22107 13672 -15808 13688
rect -22107 13608 -15892 13672
rect -15828 13608 -15808 13672
rect -22107 13592 -15808 13608
rect -22107 13528 -15892 13592
rect -15828 13528 -15808 13592
rect -22107 13512 -15808 13528
rect -22107 13448 -15892 13512
rect -15828 13448 -15808 13512
rect -22107 13432 -15808 13448
rect -22107 13368 -15892 13432
rect -15828 13368 -15808 13432
rect -22107 13352 -15808 13368
rect -22107 13288 -15892 13352
rect -15828 13288 -15808 13352
rect -22107 13272 -15808 13288
rect -22107 13208 -15892 13272
rect -15828 13208 -15808 13272
rect -22107 13192 -15808 13208
rect -22107 13128 -15892 13192
rect -15828 13128 -15808 13192
rect -22107 13112 -15808 13128
rect -22107 13048 -15892 13112
rect -15828 13048 -15808 13112
rect -22107 13032 -15808 13048
rect -22107 12968 -15892 13032
rect -15828 12968 -15808 13032
rect -22107 12952 -15808 12968
rect -22107 12888 -15892 12952
rect -15828 12888 -15808 12952
rect -22107 12872 -15808 12888
rect -22107 12808 -15892 12872
rect -15828 12808 -15808 12872
rect -22107 12792 -15808 12808
rect -22107 12728 -15892 12792
rect -15828 12728 -15808 12792
rect -22107 12712 -15808 12728
rect -22107 12648 -15892 12712
rect -15828 12648 -15808 12712
rect -22107 12632 -15808 12648
rect -22107 12568 -15892 12632
rect -15828 12568 -15808 12632
rect -22107 12552 -15808 12568
rect -22107 12488 -15892 12552
rect -15828 12488 -15808 12552
rect -22107 12472 -15808 12488
rect -22107 12408 -15892 12472
rect -15828 12408 -15808 12472
rect -22107 12392 -15808 12408
rect -22107 12328 -15892 12392
rect -15828 12328 -15808 12392
rect -22107 12312 -15808 12328
rect -22107 12248 -15892 12312
rect -15828 12248 -15808 12312
rect -22107 12232 -15808 12248
rect -22107 12168 -15892 12232
rect -15828 12168 -15808 12232
rect -22107 12152 -15808 12168
rect -22107 12088 -15892 12152
rect -15828 12088 -15808 12152
rect -22107 12072 -15808 12088
rect -22107 12008 -15892 12072
rect -15828 12008 -15808 12072
rect -22107 11992 -15808 12008
rect -22107 11928 -15892 11992
rect -15828 11928 -15808 11992
rect -22107 11912 -15808 11928
rect -22107 11848 -15892 11912
rect -15828 11848 -15808 11912
rect -22107 11832 -15808 11848
rect -22107 11768 -15892 11832
rect -15828 11768 -15808 11832
rect -22107 11752 -15808 11768
rect -22107 11688 -15892 11752
rect -15828 11688 -15808 11752
rect -22107 11672 -15808 11688
rect -22107 11608 -15892 11672
rect -15828 11608 -15808 11672
rect -22107 11592 -15808 11608
rect -22107 11528 -15892 11592
rect -15828 11528 -15808 11592
rect -22107 11512 -15808 11528
rect -22107 11448 -15892 11512
rect -15828 11448 -15808 11512
rect -22107 11432 -15808 11448
rect -22107 11368 -15892 11432
rect -15828 11368 -15808 11432
rect -22107 11352 -15808 11368
rect -22107 11288 -15892 11352
rect -15828 11288 -15808 11352
rect -22107 11272 -15808 11288
rect -22107 11208 -15892 11272
rect -15828 11208 -15808 11272
rect -22107 11192 -15808 11208
rect -22107 11128 -15892 11192
rect -15828 11128 -15808 11192
rect -22107 11112 -15808 11128
rect -22107 11048 -15892 11112
rect -15828 11048 -15808 11112
rect -22107 11032 -15808 11048
rect -22107 10968 -15892 11032
rect -15828 10968 -15808 11032
rect -22107 10952 -15808 10968
rect -22107 10888 -15892 10952
rect -15828 10888 -15808 10952
rect -22107 10872 -15808 10888
rect -22107 10808 -15892 10872
rect -15828 10808 -15808 10872
rect -22107 10792 -15808 10808
rect -22107 10728 -15892 10792
rect -15828 10728 -15808 10792
rect -22107 10712 -15808 10728
rect -22107 10648 -15892 10712
rect -15828 10648 -15808 10712
rect -22107 10632 -15808 10648
rect -22107 10568 -15892 10632
rect -15828 10568 -15808 10632
rect -22107 10552 -15808 10568
rect -22107 10488 -15892 10552
rect -15828 10488 -15808 10552
rect -22107 10472 -15808 10488
rect -22107 10408 -15892 10472
rect -15828 10408 -15808 10472
rect -22107 10392 -15808 10408
rect -22107 10328 -15892 10392
rect -15828 10328 -15808 10392
rect -22107 10312 -15808 10328
rect -22107 10248 -15892 10312
rect -15828 10248 -15808 10312
rect -22107 10232 -15808 10248
rect -22107 10168 -15892 10232
rect -15828 10168 -15808 10232
rect -22107 10152 -15808 10168
rect -22107 10088 -15892 10152
rect -15828 10088 -15808 10152
rect -22107 10072 -15808 10088
rect -22107 10008 -15892 10072
rect -15828 10008 -15808 10072
rect -22107 9992 -15808 10008
rect -22107 9928 -15892 9992
rect -15828 9928 -15808 9992
rect -22107 9912 -15808 9928
rect -22107 9848 -15892 9912
rect -15828 9848 -15808 9912
rect -22107 9832 -15808 9848
rect -22107 9768 -15892 9832
rect -15828 9768 -15808 9832
rect -22107 9752 -15808 9768
rect -22107 9688 -15892 9752
rect -15828 9688 -15808 9752
rect -22107 9672 -15808 9688
rect -22107 9608 -15892 9672
rect -15828 9608 -15808 9672
rect -22107 9592 -15808 9608
rect -22107 9528 -15892 9592
rect -15828 9528 -15808 9592
rect -22107 9500 -15808 9528
rect -15788 15672 -9489 15700
rect -15788 15608 -9573 15672
rect -9509 15608 -9489 15672
rect -15788 15592 -9489 15608
rect -15788 15528 -9573 15592
rect -9509 15528 -9489 15592
rect -15788 15512 -9489 15528
rect -15788 15448 -9573 15512
rect -9509 15448 -9489 15512
rect -15788 15432 -9489 15448
rect -15788 15368 -9573 15432
rect -9509 15368 -9489 15432
rect -15788 15352 -9489 15368
rect -15788 15288 -9573 15352
rect -9509 15288 -9489 15352
rect -15788 15272 -9489 15288
rect -15788 15208 -9573 15272
rect -9509 15208 -9489 15272
rect -15788 15192 -9489 15208
rect -15788 15128 -9573 15192
rect -9509 15128 -9489 15192
rect -15788 15112 -9489 15128
rect -15788 15048 -9573 15112
rect -9509 15048 -9489 15112
rect -15788 15032 -9489 15048
rect -15788 14968 -9573 15032
rect -9509 14968 -9489 15032
rect -15788 14952 -9489 14968
rect -15788 14888 -9573 14952
rect -9509 14888 -9489 14952
rect -15788 14872 -9489 14888
rect -15788 14808 -9573 14872
rect -9509 14808 -9489 14872
rect -15788 14792 -9489 14808
rect -15788 14728 -9573 14792
rect -9509 14728 -9489 14792
rect -15788 14712 -9489 14728
rect -15788 14648 -9573 14712
rect -9509 14648 -9489 14712
rect -15788 14632 -9489 14648
rect -15788 14568 -9573 14632
rect -9509 14568 -9489 14632
rect -15788 14552 -9489 14568
rect -15788 14488 -9573 14552
rect -9509 14488 -9489 14552
rect -15788 14472 -9489 14488
rect -15788 14408 -9573 14472
rect -9509 14408 -9489 14472
rect -15788 14392 -9489 14408
rect -15788 14328 -9573 14392
rect -9509 14328 -9489 14392
rect -15788 14312 -9489 14328
rect -15788 14248 -9573 14312
rect -9509 14248 -9489 14312
rect -15788 14232 -9489 14248
rect -15788 14168 -9573 14232
rect -9509 14168 -9489 14232
rect -15788 14152 -9489 14168
rect -15788 14088 -9573 14152
rect -9509 14088 -9489 14152
rect -15788 14072 -9489 14088
rect -15788 14008 -9573 14072
rect -9509 14008 -9489 14072
rect -15788 13992 -9489 14008
rect -15788 13928 -9573 13992
rect -9509 13928 -9489 13992
rect -15788 13912 -9489 13928
rect -15788 13848 -9573 13912
rect -9509 13848 -9489 13912
rect -15788 13832 -9489 13848
rect -15788 13768 -9573 13832
rect -9509 13768 -9489 13832
rect -15788 13752 -9489 13768
rect -15788 13688 -9573 13752
rect -9509 13688 -9489 13752
rect -15788 13672 -9489 13688
rect -15788 13608 -9573 13672
rect -9509 13608 -9489 13672
rect -15788 13592 -9489 13608
rect -15788 13528 -9573 13592
rect -9509 13528 -9489 13592
rect -15788 13512 -9489 13528
rect -15788 13448 -9573 13512
rect -9509 13448 -9489 13512
rect -15788 13432 -9489 13448
rect -15788 13368 -9573 13432
rect -9509 13368 -9489 13432
rect -15788 13352 -9489 13368
rect -15788 13288 -9573 13352
rect -9509 13288 -9489 13352
rect -15788 13272 -9489 13288
rect -15788 13208 -9573 13272
rect -9509 13208 -9489 13272
rect -15788 13192 -9489 13208
rect -15788 13128 -9573 13192
rect -9509 13128 -9489 13192
rect -15788 13112 -9489 13128
rect -15788 13048 -9573 13112
rect -9509 13048 -9489 13112
rect -15788 13032 -9489 13048
rect -15788 12968 -9573 13032
rect -9509 12968 -9489 13032
rect -15788 12952 -9489 12968
rect -15788 12888 -9573 12952
rect -9509 12888 -9489 12952
rect -15788 12872 -9489 12888
rect -15788 12808 -9573 12872
rect -9509 12808 -9489 12872
rect -15788 12792 -9489 12808
rect -15788 12728 -9573 12792
rect -9509 12728 -9489 12792
rect -15788 12712 -9489 12728
rect -15788 12648 -9573 12712
rect -9509 12648 -9489 12712
rect -15788 12632 -9489 12648
rect -15788 12568 -9573 12632
rect -9509 12568 -9489 12632
rect -15788 12552 -9489 12568
rect -15788 12488 -9573 12552
rect -9509 12488 -9489 12552
rect -15788 12472 -9489 12488
rect -15788 12408 -9573 12472
rect -9509 12408 -9489 12472
rect -15788 12392 -9489 12408
rect -15788 12328 -9573 12392
rect -9509 12328 -9489 12392
rect -15788 12312 -9489 12328
rect -15788 12248 -9573 12312
rect -9509 12248 -9489 12312
rect -15788 12232 -9489 12248
rect -15788 12168 -9573 12232
rect -9509 12168 -9489 12232
rect -15788 12152 -9489 12168
rect -15788 12088 -9573 12152
rect -9509 12088 -9489 12152
rect -15788 12072 -9489 12088
rect -15788 12008 -9573 12072
rect -9509 12008 -9489 12072
rect -15788 11992 -9489 12008
rect -15788 11928 -9573 11992
rect -9509 11928 -9489 11992
rect -15788 11912 -9489 11928
rect -15788 11848 -9573 11912
rect -9509 11848 -9489 11912
rect -15788 11832 -9489 11848
rect -15788 11768 -9573 11832
rect -9509 11768 -9489 11832
rect -15788 11752 -9489 11768
rect -15788 11688 -9573 11752
rect -9509 11688 -9489 11752
rect -15788 11672 -9489 11688
rect -15788 11608 -9573 11672
rect -9509 11608 -9489 11672
rect -15788 11592 -9489 11608
rect -15788 11528 -9573 11592
rect -9509 11528 -9489 11592
rect -15788 11512 -9489 11528
rect -15788 11448 -9573 11512
rect -9509 11448 -9489 11512
rect -15788 11432 -9489 11448
rect -15788 11368 -9573 11432
rect -9509 11368 -9489 11432
rect -15788 11352 -9489 11368
rect -15788 11288 -9573 11352
rect -9509 11288 -9489 11352
rect -15788 11272 -9489 11288
rect -15788 11208 -9573 11272
rect -9509 11208 -9489 11272
rect -15788 11192 -9489 11208
rect -15788 11128 -9573 11192
rect -9509 11128 -9489 11192
rect -15788 11112 -9489 11128
rect -15788 11048 -9573 11112
rect -9509 11048 -9489 11112
rect -15788 11032 -9489 11048
rect -15788 10968 -9573 11032
rect -9509 10968 -9489 11032
rect -15788 10952 -9489 10968
rect -15788 10888 -9573 10952
rect -9509 10888 -9489 10952
rect -15788 10872 -9489 10888
rect -15788 10808 -9573 10872
rect -9509 10808 -9489 10872
rect -15788 10792 -9489 10808
rect -15788 10728 -9573 10792
rect -9509 10728 -9489 10792
rect -15788 10712 -9489 10728
rect -15788 10648 -9573 10712
rect -9509 10648 -9489 10712
rect -15788 10632 -9489 10648
rect -15788 10568 -9573 10632
rect -9509 10568 -9489 10632
rect -15788 10552 -9489 10568
rect -15788 10488 -9573 10552
rect -9509 10488 -9489 10552
rect -15788 10472 -9489 10488
rect -15788 10408 -9573 10472
rect -9509 10408 -9489 10472
rect -15788 10392 -9489 10408
rect -15788 10328 -9573 10392
rect -9509 10328 -9489 10392
rect -15788 10312 -9489 10328
rect -15788 10248 -9573 10312
rect -9509 10248 -9489 10312
rect -15788 10232 -9489 10248
rect -15788 10168 -9573 10232
rect -9509 10168 -9489 10232
rect -15788 10152 -9489 10168
rect -15788 10088 -9573 10152
rect -9509 10088 -9489 10152
rect -15788 10072 -9489 10088
rect -15788 10008 -9573 10072
rect -9509 10008 -9489 10072
rect -15788 9992 -9489 10008
rect -15788 9928 -9573 9992
rect -9509 9928 -9489 9992
rect -15788 9912 -9489 9928
rect -15788 9848 -9573 9912
rect -9509 9848 -9489 9912
rect -15788 9832 -9489 9848
rect -15788 9768 -9573 9832
rect -9509 9768 -9489 9832
rect -15788 9752 -9489 9768
rect -15788 9688 -9573 9752
rect -9509 9688 -9489 9752
rect -15788 9672 -9489 9688
rect -15788 9608 -9573 9672
rect -9509 9608 -9489 9672
rect -15788 9592 -9489 9608
rect -15788 9528 -9573 9592
rect -9509 9528 -9489 9592
rect -15788 9500 -9489 9528
rect -9469 15672 -3170 15700
rect -9469 15608 -3254 15672
rect -3190 15608 -3170 15672
rect -9469 15592 -3170 15608
rect -9469 15528 -3254 15592
rect -3190 15528 -3170 15592
rect -9469 15512 -3170 15528
rect -9469 15448 -3254 15512
rect -3190 15448 -3170 15512
rect -9469 15432 -3170 15448
rect -9469 15368 -3254 15432
rect -3190 15368 -3170 15432
rect -9469 15352 -3170 15368
rect -9469 15288 -3254 15352
rect -3190 15288 -3170 15352
rect -9469 15272 -3170 15288
rect -9469 15208 -3254 15272
rect -3190 15208 -3170 15272
rect -9469 15192 -3170 15208
rect -9469 15128 -3254 15192
rect -3190 15128 -3170 15192
rect -9469 15112 -3170 15128
rect -9469 15048 -3254 15112
rect -3190 15048 -3170 15112
rect -9469 15032 -3170 15048
rect -9469 14968 -3254 15032
rect -3190 14968 -3170 15032
rect -9469 14952 -3170 14968
rect -9469 14888 -3254 14952
rect -3190 14888 -3170 14952
rect -9469 14872 -3170 14888
rect -9469 14808 -3254 14872
rect -3190 14808 -3170 14872
rect -9469 14792 -3170 14808
rect -9469 14728 -3254 14792
rect -3190 14728 -3170 14792
rect -9469 14712 -3170 14728
rect -9469 14648 -3254 14712
rect -3190 14648 -3170 14712
rect -9469 14632 -3170 14648
rect -9469 14568 -3254 14632
rect -3190 14568 -3170 14632
rect -9469 14552 -3170 14568
rect -9469 14488 -3254 14552
rect -3190 14488 -3170 14552
rect -9469 14472 -3170 14488
rect -9469 14408 -3254 14472
rect -3190 14408 -3170 14472
rect -9469 14392 -3170 14408
rect -9469 14328 -3254 14392
rect -3190 14328 -3170 14392
rect -9469 14312 -3170 14328
rect -9469 14248 -3254 14312
rect -3190 14248 -3170 14312
rect -9469 14232 -3170 14248
rect -9469 14168 -3254 14232
rect -3190 14168 -3170 14232
rect -9469 14152 -3170 14168
rect -9469 14088 -3254 14152
rect -3190 14088 -3170 14152
rect -9469 14072 -3170 14088
rect -9469 14008 -3254 14072
rect -3190 14008 -3170 14072
rect -9469 13992 -3170 14008
rect -9469 13928 -3254 13992
rect -3190 13928 -3170 13992
rect -9469 13912 -3170 13928
rect -9469 13848 -3254 13912
rect -3190 13848 -3170 13912
rect -9469 13832 -3170 13848
rect -9469 13768 -3254 13832
rect -3190 13768 -3170 13832
rect -9469 13752 -3170 13768
rect -9469 13688 -3254 13752
rect -3190 13688 -3170 13752
rect -9469 13672 -3170 13688
rect -9469 13608 -3254 13672
rect -3190 13608 -3170 13672
rect -9469 13592 -3170 13608
rect -9469 13528 -3254 13592
rect -3190 13528 -3170 13592
rect -9469 13512 -3170 13528
rect -9469 13448 -3254 13512
rect -3190 13448 -3170 13512
rect -9469 13432 -3170 13448
rect -9469 13368 -3254 13432
rect -3190 13368 -3170 13432
rect -9469 13352 -3170 13368
rect -9469 13288 -3254 13352
rect -3190 13288 -3170 13352
rect -9469 13272 -3170 13288
rect -9469 13208 -3254 13272
rect -3190 13208 -3170 13272
rect -9469 13192 -3170 13208
rect -9469 13128 -3254 13192
rect -3190 13128 -3170 13192
rect -9469 13112 -3170 13128
rect -9469 13048 -3254 13112
rect -3190 13048 -3170 13112
rect -9469 13032 -3170 13048
rect -9469 12968 -3254 13032
rect -3190 12968 -3170 13032
rect -9469 12952 -3170 12968
rect -9469 12888 -3254 12952
rect -3190 12888 -3170 12952
rect -9469 12872 -3170 12888
rect -9469 12808 -3254 12872
rect -3190 12808 -3170 12872
rect -9469 12792 -3170 12808
rect -9469 12728 -3254 12792
rect -3190 12728 -3170 12792
rect -9469 12712 -3170 12728
rect -9469 12648 -3254 12712
rect -3190 12648 -3170 12712
rect -9469 12632 -3170 12648
rect -9469 12568 -3254 12632
rect -3190 12568 -3170 12632
rect -9469 12552 -3170 12568
rect -9469 12488 -3254 12552
rect -3190 12488 -3170 12552
rect -9469 12472 -3170 12488
rect -9469 12408 -3254 12472
rect -3190 12408 -3170 12472
rect -9469 12392 -3170 12408
rect -9469 12328 -3254 12392
rect -3190 12328 -3170 12392
rect -9469 12312 -3170 12328
rect -9469 12248 -3254 12312
rect -3190 12248 -3170 12312
rect -9469 12232 -3170 12248
rect -9469 12168 -3254 12232
rect -3190 12168 -3170 12232
rect -9469 12152 -3170 12168
rect -9469 12088 -3254 12152
rect -3190 12088 -3170 12152
rect -9469 12072 -3170 12088
rect -9469 12008 -3254 12072
rect -3190 12008 -3170 12072
rect -9469 11992 -3170 12008
rect -9469 11928 -3254 11992
rect -3190 11928 -3170 11992
rect -9469 11912 -3170 11928
rect -9469 11848 -3254 11912
rect -3190 11848 -3170 11912
rect -9469 11832 -3170 11848
rect -9469 11768 -3254 11832
rect -3190 11768 -3170 11832
rect -9469 11752 -3170 11768
rect -9469 11688 -3254 11752
rect -3190 11688 -3170 11752
rect -9469 11672 -3170 11688
rect -9469 11608 -3254 11672
rect -3190 11608 -3170 11672
rect -9469 11592 -3170 11608
rect -9469 11528 -3254 11592
rect -3190 11528 -3170 11592
rect -9469 11512 -3170 11528
rect -9469 11448 -3254 11512
rect -3190 11448 -3170 11512
rect -9469 11432 -3170 11448
rect -9469 11368 -3254 11432
rect -3190 11368 -3170 11432
rect -9469 11352 -3170 11368
rect -9469 11288 -3254 11352
rect -3190 11288 -3170 11352
rect -9469 11272 -3170 11288
rect -9469 11208 -3254 11272
rect -3190 11208 -3170 11272
rect -9469 11192 -3170 11208
rect -9469 11128 -3254 11192
rect -3190 11128 -3170 11192
rect -9469 11112 -3170 11128
rect -9469 11048 -3254 11112
rect -3190 11048 -3170 11112
rect -9469 11032 -3170 11048
rect -9469 10968 -3254 11032
rect -3190 10968 -3170 11032
rect -9469 10952 -3170 10968
rect -9469 10888 -3254 10952
rect -3190 10888 -3170 10952
rect -9469 10872 -3170 10888
rect -9469 10808 -3254 10872
rect -3190 10808 -3170 10872
rect -9469 10792 -3170 10808
rect -9469 10728 -3254 10792
rect -3190 10728 -3170 10792
rect -9469 10712 -3170 10728
rect -9469 10648 -3254 10712
rect -3190 10648 -3170 10712
rect -9469 10632 -3170 10648
rect -9469 10568 -3254 10632
rect -3190 10568 -3170 10632
rect -9469 10552 -3170 10568
rect -9469 10488 -3254 10552
rect -3190 10488 -3170 10552
rect -9469 10472 -3170 10488
rect -9469 10408 -3254 10472
rect -3190 10408 -3170 10472
rect -9469 10392 -3170 10408
rect -9469 10328 -3254 10392
rect -3190 10328 -3170 10392
rect -9469 10312 -3170 10328
rect -9469 10248 -3254 10312
rect -3190 10248 -3170 10312
rect -9469 10232 -3170 10248
rect -9469 10168 -3254 10232
rect -3190 10168 -3170 10232
rect -9469 10152 -3170 10168
rect -9469 10088 -3254 10152
rect -3190 10088 -3170 10152
rect -9469 10072 -3170 10088
rect -9469 10008 -3254 10072
rect -3190 10008 -3170 10072
rect -9469 9992 -3170 10008
rect -9469 9928 -3254 9992
rect -3190 9928 -3170 9992
rect -9469 9912 -3170 9928
rect -9469 9848 -3254 9912
rect -3190 9848 -3170 9912
rect -9469 9832 -3170 9848
rect -9469 9768 -3254 9832
rect -3190 9768 -3170 9832
rect -9469 9752 -3170 9768
rect -9469 9688 -3254 9752
rect -3190 9688 -3170 9752
rect -9469 9672 -3170 9688
rect -9469 9608 -3254 9672
rect -3190 9608 -3170 9672
rect -9469 9592 -3170 9608
rect -9469 9528 -3254 9592
rect -3190 9528 -3170 9592
rect -9469 9500 -3170 9528
rect -3150 15672 3149 15700
rect -3150 15608 3065 15672
rect 3129 15608 3149 15672
rect -3150 15592 3149 15608
rect -3150 15528 3065 15592
rect 3129 15528 3149 15592
rect -3150 15512 3149 15528
rect -3150 15448 3065 15512
rect 3129 15448 3149 15512
rect -3150 15432 3149 15448
rect -3150 15368 3065 15432
rect 3129 15368 3149 15432
rect -3150 15352 3149 15368
rect -3150 15288 3065 15352
rect 3129 15288 3149 15352
rect -3150 15272 3149 15288
rect -3150 15208 3065 15272
rect 3129 15208 3149 15272
rect -3150 15192 3149 15208
rect -3150 15128 3065 15192
rect 3129 15128 3149 15192
rect -3150 15112 3149 15128
rect -3150 15048 3065 15112
rect 3129 15048 3149 15112
rect -3150 15032 3149 15048
rect -3150 14968 3065 15032
rect 3129 14968 3149 15032
rect -3150 14952 3149 14968
rect -3150 14888 3065 14952
rect 3129 14888 3149 14952
rect -3150 14872 3149 14888
rect -3150 14808 3065 14872
rect 3129 14808 3149 14872
rect -3150 14792 3149 14808
rect -3150 14728 3065 14792
rect 3129 14728 3149 14792
rect -3150 14712 3149 14728
rect -3150 14648 3065 14712
rect 3129 14648 3149 14712
rect -3150 14632 3149 14648
rect -3150 14568 3065 14632
rect 3129 14568 3149 14632
rect -3150 14552 3149 14568
rect -3150 14488 3065 14552
rect 3129 14488 3149 14552
rect -3150 14472 3149 14488
rect -3150 14408 3065 14472
rect 3129 14408 3149 14472
rect -3150 14392 3149 14408
rect -3150 14328 3065 14392
rect 3129 14328 3149 14392
rect -3150 14312 3149 14328
rect -3150 14248 3065 14312
rect 3129 14248 3149 14312
rect -3150 14232 3149 14248
rect -3150 14168 3065 14232
rect 3129 14168 3149 14232
rect -3150 14152 3149 14168
rect -3150 14088 3065 14152
rect 3129 14088 3149 14152
rect -3150 14072 3149 14088
rect -3150 14008 3065 14072
rect 3129 14008 3149 14072
rect -3150 13992 3149 14008
rect -3150 13928 3065 13992
rect 3129 13928 3149 13992
rect -3150 13912 3149 13928
rect -3150 13848 3065 13912
rect 3129 13848 3149 13912
rect -3150 13832 3149 13848
rect -3150 13768 3065 13832
rect 3129 13768 3149 13832
rect -3150 13752 3149 13768
rect -3150 13688 3065 13752
rect 3129 13688 3149 13752
rect -3150 13672 3149 13688
rect -3150 13608 3065 13672
rect 3129 13608 3149 13672
rect -3150 13592 3149 13608
rect -3150 13528 3065 13592
rect 3129 13528 3149 13592
rect -3150 13512 3149 13528
rect -3150 13448 3065 13512
rect 3129 13448 3149 13512
rect -3150 13432 3149 13448
rect -3150 13368 3065 13432
rect 3129 13368 3149 13432
rect -3150 13352 3149 13368
rect -3150 13288 3065 13352
rect 3129 13288 3149 13352
rect -3150 13272 3149 13288
rect -3150 13208 3065 13272
rect 3129 13208 3149 13272
rect -3150 13192 3149 13208
rect -3150 13128 3065 13192
rect 3129 13128 3149 13192
rect -3150 13112 3149 13128
rect -3150 13048 3065 13112
rect 3129 13048 3149 13112
rect -3150 13032 3149 13048
rect -3150 12968 3065 13032
rect 3129 12968 3149 13032
rect -3150 12952 3149 12968
rect -3150 12888 3065 12952
rect 3129 12888 3149 12952
rect -3150 12872 3149 12888
rect -3150 12808 3065 12872
rect 3129 12808 3149 12872
rect -3150 12792 3149 12808
rect -3150 12728 3065 12792
rect 3129 12728 3149 12792
rect -3150 12712 3149 12728
rect -3150 12648 3065 12712
rect 3129 12648 3149 12712
rect -3150 12632 3149 12648
rect -3150 12568 3065 12632
rect 3129 12568 3149 12632
rect -3150 12552 3149 12568
rect -3150 12488 3065 12552
rect 3129 12488 3149 12552
rect -3150 12472 3149 12488
rect -3150 12408 3065 12472
rect 3129 12408 3149 12472
rect -3150 12392 3149 12408
rect -3150 12328 3065 12392
rect 3129 12328 3149 12392
rect -3150 12312 3149 12328
rect -3150 12248 3065 12312
rect 3129 12248 3149 12312
rect -3150 12232 3149 12248
rect -3150 12168 3065 12232
rect 3129 12168 3149 12232
rect -3150 12152 3149 12168
rect -3150 12088 3065 12152
rect 3129 12088 3149 12152
rect -3150 12072 3149 12088
rect -3150 12008 3065 12072
rect 3129 12008 3149 12072
rect -3150 11992 3149 12008
rect -3150 11928 3065 11992
rect 3129 11928 3149 11992
rect -3150 11912 3149 11928
rect -3150 11848 3065 11912
rect 3129 11848 3149 11912
rect -3150 11832 3149 11848
rect -3150 11768 3065 11832
rect 3129 11768 3149 11832
rect -3150 11752 3149 11768
rect -3150 11688 3065 11752
rect 3129 11688 3149 11752
rect -3150 11672 3149 11688
rect -3150 11608 3065 11672
rect 3129 11608 3149 11672
rect -3150 11592 3149 11608
rect -3150 11528 3065 11592
rect 3129 11528 3149 11592
rect -3150 11512 3149 11528
rect -3150 11448 3065 11512
rect 3129 11448 3149 11512
rect -3150 11432 3149 11448
rect -3150 11368 3065 11432
rect 3129 11368 3149 11432
rect -3150 11352 3149 11368
rect -3150 11288 3065 11352
rect 3129 11288 3149 11352
rect -3150 11272 3149 11288
rect -3150 11208 3065 11272
rect 3129 11208 3149 11272
rect -3150 11192 3149 11208
rect -3150 11128 3065 11192
rect 3129 11128 3149 11192
rect -3150 11112 3149 11128
rect -3150 11048 3065 11112
rect 3129 11048 3149 11112
rect -3150 11032 3149 11048
rect -3150 10968 3065 11032
rect 3129 10968 3149 11032
rect -3150 10952 3149 10968
rect -3150 10888 3065 10952
rect 3129 10888 3149 10952
rect -3150 10872 3149 10888
rect -3150 10808 3065 10872
rect 3129 10808 3149 10872
rect -3150 10792 3149 10808
rect -3150 10728 3065 10792
rect 3129 10728 3149 10792
rect -3150 10712 3149 10728
rect -3150 10648 3065 10712
rect 3129 10648 3149 10712
rect -3150 10632 3149 10648
rect -3150 10568 3065 10632
rect 3129 10568 3149 10632
rect -3150 10552 3149 10568
rect -3150 10488 3065 10552
rect 3129 10488 3149 10552
rect -3150 10472 3149 10488
rect -3150 10408 3065 10472
rect 3129 10408 3149 10472
rect -3150 10392 3149 10408
rect -3150 10328 3065 10392
rect 3129 10328 3149 10392
rect -3150 10312 3149 10328
rect -3150 10248 3065 10312
rect 3129 10248 3149 10312
rect -3150 10232 3149 10248
rect -3150 10168 3065 10232
rect 3129 10168 3149 10232
rect -3150 10152 3149 10168
rect -3150 10088 3065 10152
rect 3129 10088 3149 10152
rect -3150 10072 3149 10088
rect -3150 10008 3065 10072
rect 3129 10008 3149 10072
rect -3150 9992 3149 10008
rect -3150 9928 3065 9992
rect 3129 9928 3149 9992
rect -3150 9912 3149 9928
rect -3150 9848 3065 9912
rect 3129 9848 3149 9912
rect -3150 9832 3149 9848
rect -3150 9768 3065 9832
rect 3129 9768 3149 9832
rect -3150 9752 3149 9768
rect -3150 9688 3065 9752
rect 3129 9688 3149 9752
rect -3150 9672 3149 9688
rect -3150 9608 3065 9672
rect 3129 9608 3149 9672
rect -3150 9592 3149 9608
rect -3150 9528 3065 9592
rect 3129 9528 3149 9592
rect -3150 9500 3149 9528
rect 3169 15672 9468 15700
rect 3169 15608 9384 15672
rect 9448 15608 9468 15672
rect 3169 15592 9468 15608
rect 3169 15528 9384 15592
rect 9448 15528 9468 15592
rect 3169 15512 9468 15528
rect 3169 15448 9384 15512
rect 9448 15448 9468 15512
rect 3169 15432 9468 15448
rect 3169 15368 9384 15432
rect 9448 15368 9468 15432
rect 3169 15352 9468 15368
rect 3169 15288 9384 15352
rect 9448 15288 9468 15352
rect 3169 15272 9468 15288
rect 3169 15208 9384 15272
rect 9448 15208 9468 15272
rect 3169 15192 9468 15208
rect 3169 15128 9384 15192
rect 9448 15128 9468 15192
rect 3169 15112 9468 15128
rect 3169 15048 9384 15112
rect 9448 15048 9468 15112
rect 3169 15032 9468 15048
rect 3169 14968 9384 15032
rect 9448 14968 9468 15032
rect 3169 14952 9468 14968
rect 3169 14888 9384 14952
rect 9448 14888 9468 14952
rect 3169 14872 9468 14888
rect 3169 14808 9384 14872
rect 9448 14808 9468 14872
rect 3169 14792 9468 14808
rect 3169 14728 9384 14792
rect 9448 14728 9468 14792
rect 3169 14712 9468 14728
rect 3169 14648 9384 14712
rect 9448 14648 9468 14712
rect 3169 14632 9468 14648
rect 3169 14568 9384 14632
rect 9448 14568 9468 14632
rect 3169 14552 9468 14568
rect 3169 14488 9384 14552
rect 9448 14488 9468 14552
rect 3169 14472 9468 14488
rect 3169 14408 9384 14472
rect 9448 14408 9468 14472
rect 3169 14392 9468 14408
rect 3169 14328 9384 14392
rect 9448 14328 9468 14392
rect 3169 14312 9468 14328
rect 3169 14248 9384 14312
rect 9448 14248 9468 14312
rect 3169 14232 9468 14248
rect 3169 14168 9384 14232
rect 9448 14168 9468 14232
rect 3169 14152 9468 14168
rect 3169 14088 9384 14152
rect 9448 14088 9468 14152
rect 3169 14072 9468 14088
rect 3169 14008 9384 14072
rect 9448 14008 9468 14072
rect 3169 13992 9468 14008
rect 3169 13928 9384 13992
rect 9448 13928 9468 13992
rect 3169 13912 9468 13928
rect 3169 13848 9384 13912
rect 9448 13848 9468 13912
rect 3169 13832 9468 13848
rect 3169 13768 9384 13832
rect 9448 13768 9468 13832
rect 3169 13752 9468 13768
rect 3169 13688 9384 13752
rect 9448 13688 9468 13752
rect 3169 13672 9468 13688
rect 3169 13608 9384 13672
rect 9448 13608 9468 13672
rect 3169 13592 9468 13608
rect 3169 13528 9384 13592
rect 9448 13528 9468 13592
rect 3169 13512 9468 13528
rect 3169 13448 9384 13512
rect 9448 13448 9468 13512
rect 3169 13432 9468 13448
rect 3169 13368 9384 13432
rect 9448 13368 9468 13432
rect 3169 13352 9468 13368
rect 3169 13288 9384 13352
rect 9448 13288 9468 13352
rect 3169 13272 9468 13288
rect 3169 13208 9384 13272
rect 9448 13208 9468 13272
rect 3169 13192 9468 13208
rect 3169 13128 9384 13192
rect 9448 13128 9468 13192
rect 3169 13112 9468 13128
rect 3169 13048 9384 13112
rect 9448 13048 9468 13112
rect 3169 13032 9468 13048
rect 3169 12968 9384 13032
rect 9448 12968 9468 13032
rect 3169 12952 9468 12968
rect 3169 12888 9384 12952
rect 9448 12888 9468 12952
rect 3169 12872 9468 12888
rect 3169 12808 9384 12872
rect 9448 12808 9468 12872
rect 3169 12792 9468 12808
rect 3169 12728 9384 12792
rect 9448 12728 9468 12792
rect 3169 12712 9468 12728
rect 3169 12648 9384 12712
rect 9448 12648 9468 12712
rect 3169 12632 9468 12648
rect 3169 12568 9384 12632
rect 9448 12568 9468 12632
rect 3169 12552 9468 12568
rect 3169 12488 9384 12552
rect 9448 12488 9468 12552
rect 3169 12472 9468 12488
rect 3169 12408 9384 12472
rect 9448 12408 9468 12472
rect 3169 12392 9468 12408
rect 3169 12328 9384 12392
rect 9448 12328 9468 12392
rect 3169 12312 9468 12328
rect 3169 12248 9384 12312
rect 9448 12248 9468 12312
rect 3169 12232 9468 12248
rect 3169 12168 9384 12232
rect 9448 12168 9468 12232
rect 3169 12152 9468 12168
rect 3169 12088 9384 12152
rect 9448 12088 9468 12152
rect 3169 12072 9468 12088
rect 3169 12008 9384 12072
rect 9448 12008 9468 12072
rect 3169 11992 9468 12008
rect 3169 11928 9384 11992
rect 9448 11928 9468 11992
rect 3169 11912 9468 11928
rect 3169 11848 9384 11912
rect 9448 11848 9468 11912
rect 3169 11832 9468 11848
rect 3169 11768 9384 11832
rect 9448 11768 9468 11832
rect 3169 11752 9468 11768
rect 3169 11688 9384 11752
rect 9448 11688 9468 11752
rect 3169 11672 9468 11688
rect 3169 11608 9384 11672
rect 9448 11608 9468 11672
rect 3169 11592 9468 11608
rect 3169 11528 9384 11592
rect 9448 11528 9468 11592
rect 3169 11512 9468 11528
rect 3169 11448 9384 11512
rect 9448 11448 9468 11512
rect 3169 11432 9468 11448
rect 3169 11368 9384 11432
rect 9448 11368 9468 11432
rect 3169 11352 9468 11368
rect 3169 11288 9384 11352
rect 9448 11288 9468 11352
rect 3169 11272 9468 11288
rect 3169 11208 9384 11272
rect 9448 11208 9468 11272
rect 3169 11192 9468 11208
rect 3169 11128 9384 11192
rect 9448 11128 9468 11192
rect 3169 11112 9468 11128
rect 3169 11048 9384 11112
rect 9448 11048 9468 11112
rect 3169 11032 9468 11048
rect 3169 10968 9384 11032
rect 9448 10968 9468 11032
rect 3169 10952 9468 10968
rect 3169 10888 9384 10952
rect 9448 10888 9468 10952
rect 3169 10872 9468 10888
rect 3169 10808 9384 10872
rect 9448 10808 9468 10872
rect 3169 10792 9468 10808
rect 3169 10728 9384 10792
rect 9448 10728 9468 10792
rect 3169 10712 9468 10728
rect 3169 10648 9384 10712
rect 9448 10648 9468 10712
rect 3169 10632 9468 10648
rect 3169 10568 9384 10632
rect 9448 10568 9468 10632
rect 3169 10552 9468 10568
rect 3169 10488 9384 10552
rect 9448 10488 9468 10552
rect 3169 10472 9468 10488
rect 3169 10408 9384 10472
rect 9448 10408 9468 10472
rect 3169 10392 9468 10408
rect 3169 10328 9384 10392
rect 9448 10328 9468 10392
rect 3169 10312 9468 10328
rect 3169 10248 9384 10312
rect 9448 10248 9468 10312
rect 3169 10232 9468 10248
rect 3169 10168 9384 10232
rect 9448 10168 9468 10232
rect 3169 10152 9468 10168
rect 3169 10088 9384 10152
rect 9448 10088 9468 10152
rect 3169 10072 9468 10088
rect 3169 10008 9384 10072
rect 9448 10008 9468 10072
rect 3169 9992 9468 10008
rect 3169 9928 9384 9992
rect 9448 9928 9468 9992
rect 3169 9912 9468 9928
rect 3169 9848 9384 9912
rect 9448 9848 9468 9912
rect 3169 9832 9468 9848
rect 3169 9768 9384 9832
rect 9448 9768 9468 9832
rect 3169 9752 9468 9768
rect 3169 9688 9384 9752
rect 9448 9688 9468 9752
rect 3169 9672 9468 9688
rect 3169 9608 9384 9672
rect 9448 9608 9468 9672
rect 3169 9592 9468 9608
rect 3169 9528 9384 9592
rect 9448 9528 9468 9592
rect 3169 9500 9468 9528
rect 9488 15672 15787 15700
rect 9488 15608 15703 15672
rect 15767 15608 15787 15672
rect 9488 15592 15787 15608
rect 9488 15528 15703 15592
rect 15767 15528 15787 15592
rect 9488 15512 15787 15528
rect 9488 15448 15703 15512
rect 15767 15448 15787 15512
rect 9488 15432 15787 15448
rect 9488 15368 15703 15432
rect 15767 15368 15787 15432
rect 9488 15352 15787 15368
rect 9488 15288 15703 15352
rect 15767 15288 15787 15352
rect 9488 15272 15787 15288
rect 9488 15208 15703 15272
rect 15767 15208 15787 15272
rect 9488 15192 15787 15208
rect 9488 15128 15703 15192
rect 15767 15128 15787 15192
rect 9488 15112 15787 15128
rect 9488 15048 15703 15112
rect 15767 15048 15787 15112
rect 9488 15032 15787 15048
rect 9488 14968 15703 15032
rect 15767 14968 15787 15032
rect 9488 14952 15787 14968
rect 9488 14888 15703 14952
rect 15767 14888 15787 14952
rect 9488 14872 15787 14888
rect 9488 14808 15703 14872
rect 15767 14808 15787 14872
rect 9488 14792 15787 14808
rect 9488 14728 15703 14792
rect 15767 14728 15787 14792
rect 9488 14712 15787 14728
rect 9488 14648 15703 14712
rect 15767 14648 15787 14712
rect 9488 14632 15787 14648
rect 9488 14568 15703 14632
rect 15767 14568 15787 14632
rect 9488 14552 15787 14568
rect 9488 14488 15703 14552
rect 15767 14488 15787 14552
rect 9488 14472 15787 14488
rect 9488 14408 15703 14472
rect 15767 14408 15787 14472
rect 9488 14392 15787 14408
rect 9488 14328 15703 14392
rect 15767 14328 15787 14392
rect 9488 14312 15787 14328
rect 9488 14248 15703 14312
rect 15767 14248 15787 14312
rect 9488 14232 15787 14248
rect 9488 14168 15703 14232
rect 15767 14168 15787 14232
rect 9488 14152 15787 14168
rect 9488 14088 15703 14152
rect 15767 14088 15787 14152
rect 9488 14072 15787 14088
rect 9488 14008 15703 14072
rect 15767 14008 15787 14072
rect 9488 13992 15787 14008
rect 9488 13928 15703 13992
rect 15767 13928 15787 13992
rect 9488 13912 15787 13928
rect 9488 13848 15703 13912
rect 15767 13848 15787 13912
rect 9488 13832 15787 13848
rect 9488 13768 15703 13832
rect 15767 13768 15787 13832
rect 9488 13752 15787 13768
rect 9488 13688 15703 13752
rect 15767 13688 15787 13752
rect 9488 13672 15787 13688
rect 9488 13608 15703 13672
rect 15767 13608 15787 13672
rect 9488 13592 15787 13608
rect 9488 13528 15703 13592
rect 15767 13528 15787 13592
rect 9488 13512 15787 13528
rect 9488 13448 15703 13512
rect 15767 13448 15787 13512
rect 9488 13432 15787 13448
rect 9488 13368 15703 13432
rect 15767 13368 15787 13432
rect 9488 13352 15787 13368
rect 9488 13288 15703 13352
rect 15767 13288 15787 13352
rect 9488 13272 15787 13288
rect 9488 13208 15703 13272
rect 15767 13208 15787 13272
rect 9488 13192 15787 13208
rect 9488 13128 15703 13192
rect 15767 13128 15787 13192
rect 9488 13112 15787 13128
rect 9488 13048 15703 13112
rect 15767 13048 15787 13112
rect 9488 13032 15787 13048
rect 9488 12968 15703 13032
rect 15767 12968 15787 13032
rect 9488 12952 15787 12968
rect 9488 12888 15703 12952
rect 15767 12888 15787 12952
rect 9488 12872 15787 12888
rect 9488 12808 15703 12872
rect 15767 12808 15787 12872
rect 9488 12792 15787 12808
rect 9488 12728 15703 12792
rect 15767 12728 15787 12792
rect 9488 12712 15787 12728
rect 9488 12648 15703 12712
rect 15767 12648 15787 12712
rect 9488 12632 15787 12648
rect 9488 12568 15703 12632
rect 15767 12568 15787 12632
rect 9488 12552 15787 12568
rect 9488 12488 15703 12552
rect 15767 12488 15787 12552
rect 9488 12472 15787 12488
rect 9488 12408 15703 12472
rect 15767 12408 15787 12472
rect 9488 12392 15787 12408
rect 9488 12328 15703 12392
rect 15767 12328 15787 12392
rect 9488 12312 15787 12328
rect 9488 12248 15703 12312
rect 15767 12248 15787 12312
rect 9488 12232 15787 12248
rect 9488 12168 15703 12232
rect 15767 12168 15787 12232
rect 9488 12152 15787 12168
rect 9488 12088 15703 12152
rect 15767 12088 15787 12152
rect 9488 12072 15787 12088
rect 9488 12008 15703 12072
rect 15767 12008 15787 12072
rect 9488 11992 15787 12008
rect 9488 11928 15703 11992
rect 15767 11928 15787 11992
rect 9488 11912 15787 11928
rect 9488 11848 15703 11912
rect 15767 11848 15787 11912
rect 9488 11832 15787 11848
rect 9488 11768 15703 11832
rect 15767 11768 15787 11832
rect 9488 11752 15787 11768
rect 9488 11688 15703 11752
rect 15767 11688 15787 11752
rect 9488 11672 15787 11688
rect 9488 11608 15703 11672
rect 15767 11608 15787 11672
rect 9488 11592 15787 11608
rect 9488 11528 15703 11592
rect 15767 11528 15787 11592
rect 9488 11512 15787 11528
rect 9488 11448 15703 11512
rect 15767 11448 15787 11512
rect 9488 11432 15787 11448
rect 9488 11368 15703 11432
rect 15767 11368 15787 11432
rect 9488 11352 15787 11368
rect 9488 11288 15703 11352
rect 15767 11288 15787 11352
rect 9488 11272 15787 11288
rect 9488 11208 15703 11272
rect 15767 11208 15787 11272
rect 9488 11192 15787 11208
rect 9488 11128 15703 11192
rect 15767 11128 15787 11192
rect 9488 11112 15787 11128
rect 9488 11048 15703 11112
rect 15767 11048 15787 11112
rect 9488 11032 15787 11048
rect 9488 10968 15703 11032
rect 15767 10968 15787 11032
rect 9488 10952 15787 10968
rect 9488 10888 15703 10952
rect 15767 10888 15787 10952
rect 9488 10872 15787 10888
rect 9488 10808 15703 10872
rect 15767 10808 15787 10872
rect 9488 10792 15787 10808
rect 9488 10728 15703 10792
rect 15767 10728 15787 10792
rect 9488 10712 15787 10728
rect 9488 10648 15703 10712
rect 15767 10648 15787 10712
rect 9488 10632 15787 10648
rect 9488 10568 15703 10632
rect 15767 10568 15787 10632
rect 9488 10552 15787 10568
rect 9488 10488 15703 10552
rect 15767 10488 15787 10552
rect 9488 10472 15787 10488
rect 9488 10408 15703 10472
rect 15767 10408 15787 10472
rect 9488 10392 15787 10408
rect 9488 10328 15703 10392
rect 15767 10328 15787 10392
rect 9488 10312 15787 10328
rect 9488 10248 15703 10312
rect 15767 10248 15787 10312
rect 9488 10232 15787 10248
rect 9488 10168 15703 10232
rect 15767 10168 15787 10232
rect 9488 10152 15787 10168
rect 9488 10088 15703 10152
rect 15767 10088 15787 10152
rect 9488 10072 15787 10088
rect 9488 10008 15703 10072
rect 15767 10008 15787 10072
rect 9488 9992 15787 10008
rect 9488 9928 15703 9992
rect 15767 9928 15787 9992
rect 9488 9912 15787 9928
rect 9488 9848 15703 9912
rect 15767 9848 15787 9912
rect 9488 9832 15787 9848
rect 9488 9768 15703 9832
rect 15767 9768 15787 9832
rect 9488 9752 15787 9768
rect 9488 9688 15703 9752
rect 15767 9688 15787 9752
rect 9488 9672 15787 9688
rect 9488 9608 15703 9672
rect 15767 9608 15787 9672
rect 9488 9592 15787 9608
rect 9488 9528 15703 9592
rect 15767 9528 15787 9592
rect 9488 9500 15787 9528
rect 15807 15672 22106 15700
rect 15807 15608 22022 15672
rect 22086 15608 22106 15672
rect 15807 15592 22106 15608
rect 15807 15528 22022 15592
rect 22086 15528 22106 15592
rect 15807 15512 22106 15528
rect 15807 15448 22022 15512
rect 22086 15448 22106 15512
rect 15807 15432 22106 15448
rect 15807 15368 22022 15432
rect 22086 15368 22106 15432
rect 15807 15352 22106 15368
rect 15807 15288 22022 15352
rect 22086 15288 22106 15352
rect 15807 15272 22106 15288
rect 15807 15208 22022 15272
rect 22086 15208 22106 15272
rect 15807 15192 22106 15208
rect 15807 15128 22022 15192
rect 22086 15128 22106 15192
rect 15807 15112 22106 15128
rect 15807 15048 22022 15112
rect 22086 15048 22106 15112
rect 15807 15032 22106 15048
rect 15807 14968 22022 15032
rect 22086 14968 22106 15032
rect 15807 14952 22106 14968
rect 15807 14888 22022 14952
rect 22086 14888 22106 14952
rect 15807 14872 22106 14888
rect 15807 14808 22022 14872
rect 22086 14808 22106 14872
rect 15807 14792 22106 14808
rect 15807 14728 22022 14792
rect 22086 14728 22106 14792
rect 15807 14712 22106 14728
rect 15807 14648 22022 14712
rect 22086 14648 22106 14712
rect 15807 14632 22106 14648
rect 15807 14568 22022 14632
rect 22086 14568 22106 14632
rect 15807 14552 22106 14568
rect 15807 14488 22022 14552
rect 22086 14488 22106 14552
rect 15807 14472 22106 14488
rect 15807 14408 22022 14472
rect 22086 14408 22106 14472
rect 15807 14392 22106 14408
rect 15807 14328 22022 14392
rect 22086 14328 22106 14392
rect 15807 14312 22106 14328
rect 15807 14248 22022 14312
rect 22086 14248 22106 14312
rect 15807 14232 22106 14248
rect 15807 14168 22022 14232
rect 22086 14168 22106 14232
rect 15807 14152 22106 14168
rect 15807 14088 22022 14152
rect 22086 14088 22106 14152
rect 15807 14072 22106 14088
rect 15807 14008 22022 14072
rect 22086 14008 22106 14072
rect 15807 13992 22106 14008
rect 15807 13928 22022 13992
rect 22086 13928 22106 13992
rect 15807 13912 22106 13928
rect 15807 13848 22022 13912
rect 22086 13848 22106 13912
rect 15807 13832 22106 13848
rect 15807 13768 22022 13832
rect 22086 13768 22106 13832
rect 15807 13752 22106 13768
rect 15807 13688 22022 13752
rect 22086 13688 22106 13752
rect 15807 13672 22106 13688
rect 15807 13608 22022 13672
rect 22086 13608 22106 13672
rect 15807 13592 22106 13608
rect 15807 13528 22022 13592
rect 22086 13528 22106 13592
rect 15807 13512 22106 13528
rect 15807 13448 22022 13512
rect 22086 13448 22106 13512
rect 15807 13432 22106 13448
rect 15807 13368 22022 13432
rect 22086 13368 22106 13432
rect 15807 13352 22106 13368
rect 15807 13288 22022 13352
rect 22086 13288 22106 13352
rect 15807 13272 22106 13288
rect 15807 13208 22022 13272
rect 22086 13208 22106 13272
rect 15807 13192 22106 13208
rect 15807 13128 22022 13192
rect 22086 13128 22106 13192
rect 15807 13112 22106 13128
rect 15807 13048 22022 13112
rect 22086 13048 22106 13112
rect 15807 13032 22106 13048
rect 15807 12968 22022 13032
rect 22086 12968 22106 13032
rect 15807 12952 22106 12968
rect 15807 12888 22022 12952
rect 22086 12888 22106 12952
rect 15807 12872 22106 12888
rect 15807 12808 22022 12872
rect 22086 12808 22106 12872
rect 15807 12792 22106 12808
rect 15807 12728 22022 12792
rect 22086 12728 22106 12792
rect 15807 12712 22106 12728
rect 15807 12648 22022 12712
rect 22086 12648 22106 12712
rect 15807 12632 22106 12648
rect 15807 12568 22022 12632
rect 22086 12568 22106 12632
rect 15807 12552 22106 12568
rect 15807 12488 22022 12552
rect 22086 12488 22106 12552
rect 15807 12472 22106 12488
rect 15807 12408 22022 12472
rect 22086 12408 22106 12472
rect 15807 12392 22106 12408
rect 15807 12328 22022 12392
rect 22086 12328 22106 12392
rect 15807 12312 22106 12328
rect 15807 12248 22022 12312
rect 22086 12248 22106 12312
rect 15807 12232 22106 12248
rect 15807 12168 22022 12232
rect 22086 12168 22106 12232
rect 15807 12152 22106 12168
rect 15807 12088 22022 12152
rect 22086 12088 22106 12152
rect 15807 12072 22106 12088
rect 15807 12008 22022 12072
rect 22086 12008 22106 12072
rect 15807 11992 22106 12008
rect 15807 11928 22022 11992
rect 22086 11928 22106 11992
rect 15807 11912 22106 11928
rect 15807 11848 22022 11912
rect 22086 11848 22106 11912
rect 15807 11832 22106 11848
rect 15807 11768 22022 11832
rect 22086 11768 22106 11832
rect 15807 11752 22106 11768
rect 15807 11688 22022 11752
rect 22086 11688 22106 11752
rect 15807 11672 22106 11688
rect 15807 11608 22022 11672
rect 22086 11608 22106 11672
rect 15807 11592 22106 11608
rect 15807 11528 22022 11592
rect 22086 11528 22106 11592
rect 15807 11512 22106 11528
rect 15807 11448 22022 11512
rect 22086 11448 22106 11512
rect 15807 11432 22106 11448
rect 15807 11368 22022 11432
rect 22086 11368 22106 11432
rect 15807 11352 22106 11368
rect 15807 11288 22022 11352
rect 22086 11288 22106 11352
rect 15807 11272 22106 11288
rect 15807 11208 22022 11272
rect 22086 11208 22106 11272
rect 15807 11192 22106 11208
rect 15807 11128 22022 11192
rect 22086 11128 22106 11192
rect 15807 11112 22106 11128
rect 15807 11048 22022 11112
rect 22086 11048 22106 11112
rect 15807 11032 22106 11048
rect 15807 10968 22022 11032
rect 22086 10968 22106 11032
rect 15807 10952 22106 10968
rect 15807 10888 22022 10952
rect 22086 10888 22106 10952
rect 15807 10872 22106 10888
rect 15807 10808 22022 10872
rect 22086 10808 22106 10872
rect 15807 10792 22106 10808
rect 15807 10728 22022 10792
rect 22086 10728 22106 10792
rect 15807 10712 22106 10728
rect 15807 10648 22022 10712
rect 22086 10648 22106 10712
rect 15807 10632 22106 10648
rect 15807 10568 22022 10632
rect 22086 10568 22106 10632
rect 15807 10552 22106 10568
rect 15807 10488 22022 10552
rect 22086 10488 22106 10552
rect 15807 10472 22106 10488
rect 15807 10408 22022 10472
rect 22086 10408 22106 10472
rect 15807 10392 22106 10408
rect 15807 10328 22022 10392
rect 22086 10328 22106 10392
rect 15807 10312 22106 10328
rect 15807 10248 22022 10312
rect 22086 10248 22106 10312
rect 15807 10232 22106 10248
rect 15807 10168 22022 10232
rect 22086 10168 22106 10232
rect 15807 10152 22106 10168
rect 15807 10088 22022 10152
rect 22086 10088 22106 10152
rect 15807 10072 22106 10088
rect 15807 10008 22022 10072
rect 22086 10008 22106 10072
rect 15807 9992 22106 10008
rect 15807 9928 22022 9992
rect 22086 9928 22106 9992
rect 15807 9912 22106 9928
rect 15807 9848 22022 9912
rect 22086 9848 22106 9912
rect 15807 9832 22106 9848
rect 15807 9768 22022 9832
rect 22086 9768 22106 9832
rect 15807 9752 22106 9768
rect 15807 9688 22022 9752
rect 22086 9688 22106 9752
rect 15807 9672 22106 9688
rect 15807 9608 22022 9672
rect 22086 9608 22106 9672
rect 15807 9592 22106 9608
rect 15807 9528 22022 9592
rect 22086 9528 22106 9592
rect 15807 9500 22106 9528
rect 22126 15672 28425 15700
rect 22126 15608 28341 15672
rect 28405 15608 28425 15672
rect 22126 15592 28425 15608
rect 22126 15528 28341 15592
rect 28405 15528 28425 15592
rect 22126 15512 28425 15528
rect 22126 15448 28341 15512
rect 28405 15448 28425 15512
rect 22126 15432 28425 15448
rect 22126 15368 28341 15432
rect 28405 15368 28425 15432
rect 22126 15352 28425 15368
rect 22126 15288 28341 15352
rect 28405 15288 28425 15352
rect 22126 15272 28425 15288
rect 22126 15208 28341 15272
rect 28405 15208 28425 15272
rect 22126 15192 28425 15208
rect 22126 15128 28341 15192
rect 28405 15128 28425 15192
rect 22126 15112 28425 15128
rect 22126 15048 28341 15112
rect 28405 15048 28425 15112
rect 22126 15032 28425 15048
rect 22126 14968 28341 15032
rect 28405 14968 28425 15032
rect 22126 14952 28425 14968
rect 22126 14888 28341 14952
rect 28405 14888 28425 14952
rect 22126 14872 28425 14888
rect 22126 14808 28341 14872
rect 28405 14808 28425 14872
rect 22126 14792 28425 14808
rect 22126 14728 28341 14792
rect 28405 14728 28425 14792
rect 22126 14712 28425 14728
rect 22126 14648 28341 14712
rect 28405 14648 28425 14712
rect 22126 14632 28425 14648
rect 22126 14568 28341 14632
rect 28405 14568 28425 14632
rect 22126 14552 28425 14568
rect 22126 14488 28341 14552
rect 28405 14488 28425 14552
rect 22126 14472 28425 14488
rect 22126 14408 28341 14472
rect 28405 14408 28425 14472
rect 22126 14392 28425 14408
rect 22126 14328 28341 14392
rect 28405 14328 28425 14392
rect 22126 14312 28425 14328
rect 22126 14248 28341 14312
rect 28405 14248 28425 14312
rect 22126 14232 28425 14248
rect 22126 14168 28341 14232
rect 28405 14168 28425 14232
rect 22126 14152 28425 14168
rect 22126 14088 28341 14152
rect 28405 14088 28425 14152
rect 22126 14072 28425 14088
rect 22126 14008 28341 14072
rect 28405 14008 28425 14072
rect 22126 13992 28425 14008
rect 22126 13928 28341 13992
rect 28405 13928 28425 13992
rect 22126 13912 28425 13928
rect 22126 13848 28341 13912
rect 28405 13848 28425 13912
rect 22126 13832 28425 13848
rect 22126 13768 28341 13832
rect 28405 13768 28425 13832
rect 22126 13752 28425 13768
rect 22126 13688 28341 13752
rect 28405 13688 28425 13752
rect 22126 13672 28425 13688
rect 22126 13608 28341 13672
rect 28405 13608 28425 13672
rect 22126 13592 28425 13608
rect 22126 13528 28341 13592
rect 28405 13528 28425 13592
rect 22126 13512 28425 13528
rect 22126 13448 28341 13512
rect 28405 13448 28425 13512
rect 22126 13432 28425 13448
rect 22126 13368 28341 13432
rect 28405 13368 28425 13432
rect 22126 13352 28425 13368
rect 22126 13288 28341 13352
rect 28405 13288 28425 13352
rect 22126 13272 28425 13288
rect 22126 13208 28341 13272
rect 28405 13208 28425 13272
rect 22126 13192 28425 13208
rect 22126 13128 28341 13192
rect 28405 13128 28425 13192
rect 22126 13112 28425 13128
rect 22126 13048 28341 13112
rect 28405 13048 28425 13112
rect 22126 13032 28425 13048
rect 22126 12968 28341 13032
rect 28405 12968 28425 13032
rect 22126 12952 28425 12968
rect 22126 12888 28341 12952
rect 28405 12888 28425 12952
rect 22126 12872 28425 12888
rect 22126 12808 28341 12872
rect 28405 12808 28425 12872
rect 22126 12792 28425 12808
rect 22126 12728 28341 12792
rect 28405 12728 28425 12792
rect 22126 12712 28425 12728
rect 22126 12648 28341 12712
rect 28405 12648 28425 12712
rect 22126 12632 28425 12648
rect 22126 12568 28341 12632
rect 28405 12568 28425 12632
rect 22126 12552 28425 12568
rect 22126 12488 28341 12552
rect 28405 12488 28425 12552
rect 22126 12472 28425 12488
rect 22126 12408 28341 12472
rect 28405 12408 28425 12472
rect 22126 12392 28425 12408
rect 22126 12328 28341 12392
rect 28405 12328 28425 12392
rect 22126 12312 28425 12328
rect 22126 12248 28341 12312
rect 28405 12248 28425 12312
rect 22126 12232 28425 12248
rect 22126 12168 28341 12232
rect 28405 12168 28425 12232
rect 22126 12152 28425 12168
rect 22126 12088 28341 12152
rect 28405 12088 28425 12152
rect 22126 12072 28425 12088
rect 22126 12008 28341 12072
rect 28405 12008 28425 12072
rect 22126 11992 28425 12008
rect 22126 11928 28341 11992
rect 28405 11928 28425 11992
rect 22126 11912 28425 11928
rect 22126 11848 28341 11912
rect 28405 11848 28425 11912
rect 22126 11832 28425 11848
rect 22126 11768 28341 11832
rect 28405 11768 28425 11832
rect 22126 11752 28425 11768
rect 22126 11688 28341 11752
rect 28405 11688 28425 11752
rect 22126 11672 28425 11688
rect 22126 11608 28341 11672
rect 28405 11608 28425 11672
rect 22126 11592 28425 11608
rect 22126 11528 28341 11592
rect 28405 11528 28425 11592
rect 22126 11512 28425 11528
rect 22126 11448 28341 11512
rect 28405 11448 28425 11512
rect 22126 11432 28425 11448
rect 22126 11368 28341 11432
rect 28405 11368 28425 11432
rect 22126 11352 28425 11368
rect 22126 11288 28341 11352
rect 28405 11288 28425 11352
rect 22126 11272 28425 11288
rect 22126 11208 28341 11272
rect 28405 11208 28425 11272
rect 22126 11192 28425 11208
rect 22126 11128 28341 11192
rect 28405 11128 28425 11192
rect 22126 11112 28425 11128
rect 22126 11048 28341 11112
rect 28405 11048 28425 11112
rect 22126 11032 28425 11048
rect 22126 10968 28341 11032
rect 28405 10968 28425 11032
rect 22126 10952 28425 10968
rect 22126 10888 28341 10952
rect 28405 10888 28425 10952
rect 22126 10872 28425 10888
rect 22126 10808 28341 10872
rect 28405 10808 28425 10872
rect 22126 10792 28425 10808
rect 22126 10728 28341 10792
rect 28405 10728 28425 10792
rect 22126 10712 28425 10728
rect 22126 10648 28341 10712
rect 28405 10648 28425 10712
rect 22126 10632 28425 10648
rect 22126 10568 28341 10632
rect 28405 10568 28425 10632
rect 22126 10552 28425 10568
rect 22126 10488 28341 10552
rect 28405 10488 28425 10552
rect 22126 10472 28425 10488
rect 22126 10408 28341 10472
rect 28405 10408 28425 10472
rect 22126 10392 28425 10408
rect 22126 10328 28341 10392
rect 28405 10328 28425 10392
rect 22126 10312 28425 10328
rect 22126 10248 28341 10312
rect 28405 10248 28425 10312
rect 22126 10232 28425 10248
rect 22126 10168 28341 10232
rect 28405 10168 28425 10232
rect 22126 10152 28425 10168
rect 22126 10088 28341 10152
rect 28405 10088 28425 10152
rect 22126 10072 28425 10088
rect 22126 10008 28341 10072
rect 28405 10008 28425 10072
rect 22126 9992 28425 10008
rect 22126 9928 28341 9992
rect 28405 9928 28425 9992
rect 22126 9912 28425 9928
rect 22126 9848 28341 9912
rect 28405 9848 28425 9912
rect 22126 9832 28425 9848
rect 22126 9768 28341 9832
rect 28405 9768 28425 9832
rect 22126 9752 28425 9768
rect 22126 9688 28341 9752
rect 28405 9688 28425 9752
rect 22126 9672 28425 9688
rect 22126 9608 28341 9672
rect 28405 9608 28425 9672
rect 22126 9592 28425 9608
rect 22126 9528 28341 9592
rect 28405 9528 28425 9592
rect 22126 9500 28425 9528
rect 28445 15672 34744 15700
rect 28445 15608 34660 15672
rect 34724 15608 34744 15672
rect 28445 15592 34744 15608
rect 28445 15528 34660 15592
rect 34724 15528 34744 15592
rect 28445 15512 34744 15528
rect 28445 15448 34660 15512
rect 34724 15448 34744 15512
rect 28445 15432 34744 15448
rect 28445 15368 34660 15432
rect 34724 15368 34744 15432
rect 28445 15352 34744 15368
rect 28445 15288 34660 15352
rect 34724 15288 34744 15352
rect 28445 15272 34744 15288
rect 28445 15208 34660 15272
rect 34724 15208 34744 15272
rect 28445 15192 34744 15208
rect 28445 15128 34660 15192
rect 34724 15128 34744 15192
rect 28445 15112 34744 15128
rect 28445 15048 34660 15112
rect 34724 15048 34744 15112
rect 28445 15032 34744 15048
rect 28445 14968 34660 15032
rect 34724 14968 34744 15032
rect 28445 14952 34744 14968
rect 28445 14888 34660 14952
rect 34724 14888 34744 14952
rect 28445 14872 34744 14888
rect 28445 14808 34660 14872
rect 34724 14808 34744 14872
rect 28445 14792 34744 14808
rect 28445 14728 34660 14792
rect 34724 14728 34744 14792
rect 28445 14712 34744 14728
rect 28445 14648 34660 14712
rect 34724 14648 34744 14712
rect 28445 14632 34744 14648
rect 28445 14568 34660 14632
rect 34724 14568 34744 14632
rect 28445 14552 34744 14568
rect 28445 14488 34660 14552
rect 34724 14488 34744 14552
rect 28445 14472 34744 14488
rect 28445 14408 34660 14472
rect 34724 14408 34744 14472
rect 28445 14392 34744 14408
rect 28445 14328 34660 14392
rect 34724 14328 34744 14392
rect 28445 14312 34744 14328
rect 28445 14248 34660 14312
rect 34724 14248 34744 14312
rect 28445 14232 34744 14248
rect 28445 14168 34660 14232
rect 34724 14168 34744 14232
rect 28445 14152 34744 14168
rect 28445 14088 34660 14152
rect 34724 14088 34744 14152
rect 28445 14072 34744 14088
rect 28445 14008 34660 14072
rect 34724 14008 34744 14072
rect 28445 13992 34744 14008
rect 28445 13928 34660 13992
rect 34724 13928 34744 13992
rect 28445 13912 34744 13928
rect 28445 13848 34660 13912
rect 34724 13848 34744 13912
rect 28445 13832 34744 13848
rect 28445 13768 34660 13832
rect 34724 13768 34744 13832
rect 28445 13752 34744 13768
rect 28445 13688 34660 13752
rect 34724 13688 34744 13752
rect 28445 13672 34744 13688
rect 28445 13608 34660 13672
rect 34724 13608 34744 13672
rect 28445 13592 34744 13608
rect 28445 13528 34660 13592
rect 34724 13528 34744 13592
rect 28445 13512 34744 13528
rect 28445 13448 34660 13512
rect 34724 13448 34744 13512
rect 28445 13432 34744 13448
rect 28445 13368 34660 13432
rect 34724 13368 34744 13432
rect 28445 13352 34744 13368
rect 28445 13288 34660 13352
rect 34724 13288 34744 13352
rect 28445 13272 34744 13288
rect 28445 13208 34660 13272
rect 34724 13208 34744 13272
rect 28445 13192 34744 13208
rect 28445 13128 34660 13192
rect 34724 13128 34744 13192
rect 28445 13112 34744 13128
rect 28445 13048 34660 13112
rect 34724 13048 34744 13112
rect 28445 13032 34744 13048
rect 28445 12968 34660 13032
rect 34724 12968 34744 13032
rect 28445 12952 34744 12968
rect 28445 12888 34660 12952
rect 34724 12888 34744 12952
rect 28445 12872 34744 12888
rect 28445 12808 34660 12872
rect 34724 12808 34744 12872
rect 28445 12792 34744 12808
rect 28445 12728 34660 12792
rect 34724 12728 34744 12792
rect 28445 12712 34744 12728
rect 28445 12648 34660 12712
rect 34724 12648 34744 12712
rect 28445 12632 34744 12648
rect 28445 12568 34660 12632
rect 34724 12568 34744 12632
rect 28445 12552 34744 12568
rect 28445 12488 34660 12552
rect 34724 12488 34744 12552
rect 28445 12472 34744 12488
rect 28445 12408 34660 12472
rect 34724 12408 34744 12472
rect 28445 12392 34744 12408
rect 28445 12328 34660 12392
rect 34724 12328 34744 12392
rect 28445 12312 34744 12328
rect 28445 12248 34660 12312
rect 34724 12248 34744 12312
rect 28445 12232 34744 12248
rect 28445 12168 34660 12232
rect 34724 12168 34744 12232
rect 28445 12152 34744 12168
rect 28445 12088 34660 12152
rect 34724 12088 34744 12152
rect 28445 12072 34744 12088
rect 28445 12008 34660 12072
rect 34724 12008 34744 12072
rect 28445 11992 34744 12008
rect 28445 11928 34660 11992
rect 34724 11928 34744 11992
rect 28445 11912 34744 11928
rect 28445 11848 34660 11912
rect 34724 11848 34744 11912
rect 28445 11832 34744 11848
rect 28445 11768 34660 11832
rect 34724 11768 34744 11832
rect 28445 11752 34744 11768
rect 28445 11688 34660 11752
rect 34724 11688 34744 11752
rect 28445 11672 34744 11688
rect 28445 11608 34660 11672
rect 34724 11608 34744 11672
rect 28445 11592 34744 11608
rect 28445 11528 34660 11592
rect 34724 11528 34744 11592
rect 28445 11512 34744 11528
rect 28445 11448 34660 11512
rect 34724 11448 34744 11512
rect 28445 11432 34744 11448
rect 28445 11368 34660 11432
rect 34724 11368 34744 11432
rect 28445 11352 34744 11368
rect 28445 11288 34660 11352
rect 34724 11288 34744 11352
rect 28445 11272 34744 11288
rect 28445 11208 34660 11272
rect 34724 11208 34744 11272
rect 28445 11192 34744 11208
rect 28445 11128 34660 11192
rect 34724 11128 34744 11192
rect 28445 11112 34744 11128
rect 28445 11048 34660 11112
rect 34724 11048 34744 11112
rect 28445 11032 34744 11048
rect 28445 10968 34660 11032
rect 34724 10968 34744 11032
rect 28445 10952 34744 10968
rect 28445 10888 34660 10952
rect 34724 10888 34744 10952
rect 28445 10872 34744 10888
rect 28445 10808 34660 10872
rect 34724 10808 34744 10872
rect 28445 10792 34744 10808
rect 28445 10728 34660 10792
rect 34724 10728 34744 10792
rect 28445 10712 34744 10728
rect 28445 10648 34660 10712
rect 34724 10648 34744 10712
rect 28445 10632 34744 10648
rect 28445 10568 34660 10632
rect 34724 10568 34744 10632
rect 28445 10552 34744 10568
rect 28445 10488 34660 10552
rect 34724 10488 34744 10552
rect 28445 10472 34744 10488
rect 28445 10408 34660 10472
rect 34724 10408 34744 10472
rect 28445 10392 34744 10408
rect 28445 10328 34660 10392
rect 34724 10328 34744 10392
rect 28445 10312 34744 10328
rect 28445 10248 34660 10312
rect 34724 10248 34744 10312
rect 28445 10232 34744 10248
rect 28445 10168 34660 10232
rect 34724 10168 34744 10232
rect 28445 10152 34744 10168
rect 28445 10088 34660 10152
rect 34724 10088 34744 10152
rect 28445 10072 34744 10088
rect 28445 10008 34660 10072
rect 34724 10008 34744 10072
rect 28445 9992 34744 10008
rect 28445 9928 34660 9992
rect 34724 9928 34744 9992
rect 28445 9912 34744 9928
rect 28445 9848 34660 9912
rect 34724 9848 34744 9912
rect 28445 9832 34744 9848
rect 28445 9768 34660 9832
rect 34724 9768 34744 9832
rect 28445 9752 34744 9768
rect 28445 9688 34660 9752
rect 34724 9688 34744 9752
rect 28445 9672 34744 9688
rect 28445 9608 34660 9672
rect 34724 9608 34744 9672
rect 28445 9592 34744 9608
rect 28445 9528 34660 9592
rect 34724 9528 34744 9592
rect 28445 9500 34744 9528
rect 34764 15672 41063 15700
rect 34764 15608 40979 15672
rect 41043 15608 41063 15672
rect 34764 15592 41063 15608
rect 34764 15528 40979 15592
rect 41043 15528 41063 15592
rect 34764 15512 41063 15528
rect 34764 15448 40979 15512
rect 41043 15448 41063 15512
rect 34764 15432 41063 15448
rect 34764 15368 40979 15432
rect 41043 15368 41063 15432
rect 34764 15352 41063 15368
rect 34764 15288 40979 15352
rect 41043 15288 41063 15352
rect 34764 15272 41063 15288
rect 34764 15208 40979 15272
rect 41043 15208 41063 15272
rect 34764 15192 41063 15208
rect 34764 15128 40979 15192
rect 41043 15128 41063 15192
rect 34764 15112 41063 15128
rect 34764 15048 40979 15112
rect 41043 15048 41063 15112
rect 34764 15032 41063 15048
rect 34764 14968 40979 15032
rect 41043 14968 41063 15032
rect 34764 14952 41063 14968
rect 34764 14888 40979 14952
rect 41043 14888 41063 14952
rect 34764 14872 41063 14888
rect 34764 14808 40979 14872
rect 41043 14808 41063 14872
rect 34764 14792 41063 14808
rect 34764 14728 40979 14792
rect 41043 14728 41063 14792
rect 34764 14712 41063 14728
rect 34764 14648 40979 14712
rect 41043 14648 41063 14712
rect 34764 14632 41063 14648
rect 34764 14568 40979 14632
rect 41043 14568 41063 14632
rect 34764 14552 41063 14568
rect 34764 14488 40979 14552
rect 41043 14488 41063 14552
rect 34764 14472 41063 14488
rect 34764 14408 40979 14472
rect 41043 14408 41063 14472
rect 34764 14392 41063 14408
rect 34764 14328 40979 14392
rect 41043 14328 41063 14392
rect 34764 14312 41063 14328
rect 34764 14248 40979 14312
rect 41043 14248 41063 14312
rect 34764 14232 41063 14248
rect 34764 14168 40979 14232
rect 41043 14168 41063 14232
rect 34764 14152 41063 14168
rect 34764 14088 40979 14152
rect 41043 14088 41063 14152
rect 34764 14072 41063 14088
rect 34764 14008 40979 14072
rect 41043 14008 41063 14072
rect 34764 13992 41063 14008
rect 34764 13928 40979 13992
rect 41043 13928 41063 13992
rect 34764 13912 41063 13928
rect 34764 13848 40979 13912
rect 41043 13848 41063 13912
rect 34764 13832 41063 13848
rect 34764 13768 40979 13832
rect 41043 13768 41063 13832
rect 34764 13752 41063 13768
rect 34764 13688 40979 13752
rect 41043 13688 41063 13752
rect 34764 13672 41063 13688
rect 34764 13608 40979 13672
rect 41043 13608 41063 13672
rect 34764 13592 41063 13608
rect 34764 13528 40979 13592
rect 41043 13528 41063 13592
rect 34764 13512 41063 13528
rect 34764 13448 40979 13512
rect 41043 13448 41063 13512
rect 34764 13432 41063 13448
rect 34764 13368 40979 13432
rect 41043 13368 41063 13432
rect 34764 13352 41063 13368
rect 34764 13288 40979 13352
rect 41043 13288 41063 13352
rect 34764 13272 41063 13288
rect 34764 13208 40979 13272
rect 41043 13208 41063 13272
rect 34764 13192 41063 13208
rect 34764 13128 40979 13192
rect 41043 13128 41063 13192
rect 34764 13112 41063 13128
rect 34764 13048 40979 13112
rect 41043 13048 41063 13112
rect 34764 13032 41063 13048
rect 34764 12968 40979 13032
rect 41043 12968 41063 13032
rect 34764 12952 41063 12968
rect 34764 12888 40979 12952
rect 41043 12888 41063 12952
rect 34764 12872 41063 12888
rect 34764 12808 40979 12872
rect 41043 12808 41063 12872
rect 34764 12792 41063 12808
rect 34764 12728 40979 12792
rect 41043 12728 41063 12792
rect 34764 12712 41063 12728
rect 34764 12648 40979 12712
rect 41043 12648 41063 12712
rect 34764 12632 41063 12648
rect 34764 12568 40979 12632
rect 41043 12568 41063 12632
rect 34764 12552 41063 12568
rect 34764 12488 40979 12552
rect 41043 12488 41063 12552
rect 34764 12472 41063 12488
rect 34764 12408 40979 12472
rect 41043 12408 41063 12472
rect 34764 12392 41063 12408
rect 34764 12328 40979 12392
rect 41043 12328 41063 12392
rect 34764 12312 41063 12328
rect 34764 12248 40979 12312
rect 41043 12248 41063 12312
rect 34764 12232 41063 12248
rect 34764 12168 40979 12232
rect 41043 12168 41063 12232
rect 34764 12152 41063 12168
rect 34764 12088 40979 12152
rect 41043 12088 41063 12152
rect 34764 12072 41063 12088
rect 34764 12008 40979 12072
rect 41043 12008 41063 12072
rect 34764 11992 41063 12008
rect 34764 11928 40979 11992
rect 41043 11928 41063 11992
rect 34764 11912 41063 11928
rect 34764 11848 40979 11912
rect 41043 11848 41063 11912
rect 34764 11832 41063 11848
rect 34764 11768 40979 11832
rect 41043 11768 41063 11832
rect 34764 11752 41063 11768
rect 34764 11688 40979 11752
rect 41043 11688 41063 11752
rect 34764 11672 41063 11688
rect 34764 11608 40979 11672
rect 41043 11608 41063 11672
rect 34764 11592 41063 11608
rect 34764 11528 40979 11592
rect 41043 11528 41063 11592
rect 34764 11512 41063 11528
rect 34764 11448 40979 11512
rect 41043 11448 41063 11512
rect 34764 11432 41063 11448
rect 34764 11368 40979 11432
rect 41043 11368 41063 11432
rect 34764 11352 41063 11368
rect 34764 11288 40979 11352
rect 41043 11288 41063 11352
rect 34764 11272 41063 11288
rect 34764 11208 40979 11272
rect 41043 11208 41063 11272
rect 34764 11192 41063 11208
rect 34764 11128 40979 11192
rect 41043 11128 41063 11192
rect 34764 11112 41063 11128
rect 34764 11048 40979 11112
rect 41043 11048 41063 11112
rect 34764 11032 41063 11048
rect 34764 10968 40979 11032
rect 41043 10968 41063 11032
rect 34764 10952 41063 10968
rect 34764 10888 40979 10952
rect 41043 10888 41063 10952
rect 34764 10872 41063 10888
rect 34764 10808 40979 10872
rect 41043 10808 41063 10872
rect 34764 10792 41063 10808
rect 34764 10728 40979 10792
rect 41043 10728 41063 10792
rect 34764 10712 41063 10728
rect 34764 10648 40979 10712
rect 41043 10648 41063 10712
rect 34764 10632 41063 10648
rect 34764 10568 40979 10632
rect 41043 10568 41063 10632
rect 34764 10552 41063 10568
rect 34764 10488 40979 10552
rect 41043 10488 41063 10552
rect 34764 10472 41063 10488
rect 34764 10408 40979 10472
rect 41043 10408 41063 10472
rect 34764 10392 41063 10408
rect 34764 10328 40979 10392
rect 41043 10328 41063 10392
rect 34764 10312 41063 10328
rect 34764 10248 40979 10312
rect 41043 10248 41063 10312
rect 34764 10232 41063 10248
rect 34764 10168 40979 10232
rect 41043 10168 41063 10232
rect 34764 10152 41063 10168
rect 34764 10088 40979 10152
rect 41043 10088 41063 10152
rect 34764 10072 41063 10088
rect 34764 10008 40979 10072
rect 41043 10008 41063 10072
rect 34764 9992 41063 10008
rect 34764 9928 40979 9992
rect 41043 9928 41063 9992
rect 34764 9912 41063 9928
rect 34764 9848 40979 9912
rect 41043 9848 41063 9912
rect 34764 9832 41063 9848
rect 34764 9768 40979 9832
rect 41043 9768 41063 9832
rect 34764 9752 41063 9768
rect 34764 9688 40979 9752
rect 41043 9688 41063 9752
rect 34764 9672 41063 9688
rect 34764 9608 40979 9672
rect 41043 9608 41063 9672
rect 34764 9592 41063 9608
rect 34764 9528 40979 9592
rect 41043 9528 41063 9592
rect 34764 9500 41063 9528
rect 41083 15672 47382 15700
rect 41083 15608 47298 15672
rect 47362 15608 47382 15672
rect 41083 15592 47382 15608
rect 41083 15528 47298 15592
rect 47362 15528 47382 15592
rect 41083 15512 47382 15528
rect 41083 15448 47298 15512
rect 47362 15448 47382 15512
rect 41083 15432 47382 15448
rect 41083 15368 47298 15432
rect 47362 15368 47382 15432
rect 41083 15352 47382 15368
rect 41083 15288 47298 15352
rect 47362 15288 47382 15352
rect 41083 15272 47382 15288
rect 41083 15208 47298 15272
rect 47362 15208 47382 15272
rect 41083 15192 47382 15208
rect 41083 15128 47298 15192
rect 47362 15128 47382 15192
rect 41083 15112 47382 15128
rect 41083 15048 47298 15112
rect 47362 15048 47382 15112
rect 41083 15032 47382 15048
rect 41083 14968 47298 15032
rect 47362 14968 47382 15032
rect 41083 14952 47382 14968
rect 41083 14888 47298 14952
rect 47362 14888 47382 14952
rect 41083 14872 47382 14888
rect 41083 14808 47298 14872
rect 47362 14808 47382 14872
rect 41083 14792 47382 14808
rect 41083 14728 47298 14792
rect 47362 14728 47382 14792
rect 41083 14712 47382 14728
rect 41083 14648 47298 14712
rect 47362 14648 47382 14712
rect 41083 14632 47382 14648
rect 41083 14568 47298 14632
rect 47362 14568 47382 14632
rect 41083 14552 47382 14568
rect 41083 14488 47298 14552
rect 47362 14488 47382 14552
rect 41083 14472 47382 14488
rect 41083 14408 47298 14472
rect 47362 14408 47382 14472
rect 41083 14392 47382 14408
rect 41083 14328 47298 14392
rect 47362 14328 47382 14392
rect 41083 14312 47382 14328
rect 41083 14248 47298 14312
rect 47362 14248 47382 14312
rect 41083 14232 47382 14248
rect 41083 14168 47298 14232
rect 47362 14168 47382 14232
rect 41083 14152 47382 14168
rect 41083 14088 47298 14152
rect 47362 14088 47382 14152
rect 41083 14072 47382 14088
rect 41083 14008 47298 14072
rect 47362 14008 47382 14072
rect 41083 13992 47382 14008
rect 41083 13928 47298 13992
rect 47362 13928 47382 13992
rect 41083 13912 47382 13928
rect 41083 13848 47298 13912
rect 47362 13848 47382 13912
rect 41083 13832 47382 13848
rect 41083 13768 47298 13832
rect 47362 13768 47382 13832
rect 41083 13752 47382 13768
rect 41083 13688 47298 13752
rect 47362 13688 47382 13752
rect 41083 13672 47382 13688
rect 41083 13608 47298 13672
rect 47362 13608 47382 13672
rect 41083 13592 47382 13608
rect 41083 13528 47298 13592
rect 47362 13528 47382 13592
rect 41083 13512 47382 13528
rect 41083 13448 47298 13512
rect 47362 13448 47382 13512
rect 41083 13432 47382 13448
rect 41083 13368 47298 13432
rect 47362 13368 47382 13432
rect 41083 13352 47382 13368
rect 41083 13288 47298 13352
rect 47362 13288 47382 13352
rect 41083 13272 47382 13288
rect 41083 13208 47298 13272
rect 47362 13208 47382 13272
rect 41083 13192 47382 13208
rect 41083 13128 47298 13192
rect 47362 13128 47382 13192
rect 41083 13112 47382 13128
rect 41083 13048 47298 13112
rect 47362 13048 47382 13112
rect 41083 13032 47382 13048
rect 41083 12968 47298 13032
rect 47362 12968 47382 13032
rect 41083 12952 47382 12968
rect 41083 12888 47298 12952
rect 47362 12888 47382 12952
rect 41083 12872 47382 12888
rect 41083 12808 47298 12872
rect 47362 12808 47382 12872
rect 41083 12792 47382 12808
rect 41083 12728 47298 12792
rect 47362 12728 47382 12792
rect 41083 12712 47382 12728
rect 41083 12648 47298 12712
rect 47362 12648 47382 12712
rect 41083 12632 47382 12648
rect 41083 12568 47298 12632
rect 47362 12568 47382 12632
rect 41083 12552 47382 12568
rect 41083 12488 47298 12552
rect 47362 12488 47382 12552
rect 41083 12472 47382 12488
rect 41083 12408 47298 12472
rect 47362 12408 47382 12472
rect 41083 12392 47382 12408
rect 41083 12328 47298 12392
rect 47362 12328 47382 12392
rect 41083 12312 47382 12328
rect 41083 12248 47298 12312
rect 47362 12248 47382 12312
rect 41083 12232 47382 12248
rect 41083 12168 47298 12232
rect 47362 12168 47382 12232
rect 41083 12152 47382 12168
rect 41083 12088 47298 12152
rect 47362 12088 47382 12152
rect 41083 12072 47382 12088
rect 41083 12008 47298 12072
rect 47362 12008 47382 12072
rect 41083 11992 47382 12008
rect 41083 11928 47298 11992
rect 47362 11928 47382 11992
rect 41083 11912 47382 11928
rect 41083 11848 47298 11912
rect 47362 11848 47382 11912
rect 41083 11832 47382 11848
rect 41083 11768 47298 11832
rect 47362 11768 47382 11832
rect 41083 11752 47382 11768
rect 41083 11688 47298 11752
rect 47362 11688 47382 11752
rect 41083 11672 47382 11688
rect 41083 11608 47298 11672
rect 47362 11608 47382 11672
rect 41083 11592 47382 11608
rect 41083 11528 47298 11592
rect 47362 11528 47382 11592
rect 41083 11512 47382 11528
rect 41083 11448 47298 11512
rect 47362 11448 47382 11512
rect 41083 11432 47382 11448
rect 41083 11368 47298 11432
rect 47362 11368 47382 11432
rect 41083 11352 47382 11368
rect 41083 11288 47298 11352
rect 47362 11288 47382 11352
rect 41083 11272 47382 11288
rect 41083 11208 47298 11272
rect 47362 11208 47382 11272
rect 41083 11192 47382 11208
rect 41083 11128 47298 11192
rect 47362 11128 47382 11192
rect 41083 11112 47382 11128
rect 41083 11048 47298 11112
rect 47362 11048 47382 11112
rect 41083 11032 47382 11048
rect 41083 10968 47298 11032
rect 47362 10968 47382 11032
rect 41083 10952 47382 10968
rect 41083 10888 47298 10952
rect 47362 10888 47382 10952
rect 41083 10872 47382 10888
rect 41083 10808 47298 10872
rect 47362 10808 47382 10872
rect 41083 10792 47382 10808
rect 41083 10728 47298 10792
rect 47362 10728 47382 10792
rect 41083 10712 47382 10728
rect 41083 10648 47298 10712
rect 47362 10648 47382 10712
rect 41083 10632 47382 10648
rect 41083 10568 47298 10632
rect 47362 10568 47382 10632
rect 41083 10552 47382 10568
rect 41083 10488 47298 10552
rect 47362 10488 47382 10552
rect 41083 10472 47382 10488
rect 41083 10408 47298 10472
rect 47362 10408 47382 10472
rect 41083 10392 47382 10408
rect 41083 10328 47298 10392
rect 47362 10328 47382 10392
rect 41083 10312 47382 10328
rect 41083 10248 47298 10312
rect 47362 10248 47382 10312
rect 41083 10232 47382 10248
rect 41083 10168 47298 10232
rect 47362 10168 47382 10232
rect 41083 10152 47382 10168
rect 41083 10088 47298 10152
rect 47362 10088 47382 10152
rect 41083 10072 47382 10088
rect 41083 10008 47298 10072
rect 47362 10008 47382 10072
rect 41083 9992 47382 10008
rect 41083 9928 47298 9992
rect 47362 9928 47382 9992
rect 41083 9912 47382 9928
rect 41083 9848 47298 9912
rect 47362 9848 47382 9912
rect 41083 9832 47382 9848
rect 41083 9768 47298 9832
rect 47362 9768 47382 9832
rect 41083 9752 47382 9768
rect 41083 9688 47298 9752
rect 47362 9688 47382 9752
rect 41083 9672 47382 9688
rect 41083 9608 47298 9672
rect 47362 9608 47382 9672
rect 41083 9592 47382 9608
rect 41083 9528 47298 9592
rect 47362 9528 47382 9592
rect 41083 9500 47382 9528
rect -47383 9372 -41084 9400
rect -47383 9308 -41168 9372
rect -41104 9308 -41084 9372
rect -47383 9292 -41084 9308
rect -47383 9228 -41168 9292
rect -41104 9228 -41084 9292
rect -47383 9212 -41084 9228
rect -47383 9148 -41168 9212
rect -41104 9148 -41084 9212
rect -47383 9132 -41084 9148
rect -47383 9068 -41168 9132
rect -41104 9068 -41084 9132
rect -47383 9052 -41084 9068
rect -47383 8988 -41168 9052
rect -41104 8988 -41084 9052
rect -47383 8972 -41084 8988
rect -47383 8908 -41168 8972
rect -41104 8908 -41084 8972
rect -47383 8892 -41084 8908
rect -47383 8828 -41168 8892
rect -41104 8828 -41084 8892
rect -47383 8812 -41084 8828
rect -47383 8748 -41168 8812
rect -41104 8748 -41084 8812
rect -47383 8732 -41084 8748
rect -47383 8668 -41168 8732
rect -41104 8668 -41084 8732
rect -47383 8652 -41084 8668
rect -47383 8588 -41168 8652
rect -41104 8588 -41084 8652
rect -47383 8572 -41084 8588
rect -47383 8508 -41168 8572
rect -41104 8508 -41084 8572
rect -47383 8492 -41084 8508
rect -47383 8428 -41168 8492
rect -41104 8428 -41084 8492
rect -47383 8412 -41084 8428
rect -47383 8348 -41168 8412
rect -41104 8348 -41084 8412
rect -47383 8332 -41084 8348
rect -47383 8268 -41168 8332
rect -41104 8268 -41084 8332
rect -47383 8252 -41084 8268
rect -47383 8188 -41168 8252
rect -41104 8188 -41084 8252
rect -47383 8172 -41084 8188
rect -47383 8108 -41168 8172
rect -41104 8108 -41084 8172
rect -47383 8092 -41084 8108
rect -47383 8028 -41168 8092
rect -41104 8028 -41084 8092
rect -47383 8012 -41084 8028
rect -47383 7948 -41168 8012
rect -41104 7948 -41084 8012
rect -47383 7932 -41084 7948
rect -47383 7868 -41168 7932
rect -41104 7868 -41084 7932
rect -47383 7852 -41084 7868
rect -47383 7788 -41168 7852
rect -41104 7788 -41084 7852
rect -47383 7772 -41084 7788
rect -47383 7708 -41168 7772
rect -41104 7708 -41084 7772
rect -47383 7692 -41084 7708
rect -47383 7628 -41168 7692
rect -41104 7628 -41084 7692
rect -47383 7612 -41084 7628
rect -47383 7548 -41168 7612
rect -41104 7548 -41084 7612
rect -47383 7532 -41084 7548
rect -47383 7468 -41168 7532
rect -41104 7468 -41084 7532
rect -47383 7452 -41084 7468
rect -47383 7388 -41168 7452
rect -41104 7388 -41084 7452
rect -47383 7372 -41084 7388
rect -47383 7308 -41168 7372
rect -41104 7308 -41084 7372
rect -47383 7292 -41084 7308
rect -47383 7228 -41168 7292
rect -41104 7228 -41084 7292
rect -47383 7212 -41084 7228
rect -47383 7148 -41168 7212
rect -41104 7148 -41084 7212
rect -47383 7132 -41084 7148
rect -47383 7068 -41168 7132
rect -41104 7068 -41084 7132
rect -47383 7052 -41084 7068
rect -47383 6988 -41168 7052
rect -41104 6988 -41084 7052
rect -47383 6972 -41084 6988
rect -47383 6908 -41168 6972
rect -41104 6908 -41084 6972
rect -47383 6892 -41084 6908
rect -47383 6828 -41168 6892
rect -41104 6828 -41084 6892
rect -47383 6812 -41084 6828
rect -47383 6748 -41168 6812
rect -41104 6748 -41084 6812
rect -47383 6732 -41084 6748
rect -47383 6668 -41168 6732
rect -41104 6668 -41084 6732
rect -47383 6652 -41084 6668
rect -47383 6588 -41168 6652
rect -41104 6588 -41084 6652
rect -47383 6572 -41084 6588
rect -47383 6508 -41168 6572
rect -41104 6508 -41084 6572
rect -47383 6492 -41084 6508
rect -47383 6428 -41168 6492
rect -41104 6428 -41084 6492
rect -47383 6412 -41084 6428
rect -47383 6348 -41168 6412
rect -41104 6348 -41084 6412
rect -47383 6332 -41084 6348
rect -47383 6268 -41168 6332
rect -41104 6268 -41084 6332
rect -47383 6252 -41084 6268
rect -47383 6188 -41168 6252
rect -41104 6188 -41084 6252
rect -47383 6172 -41084 6188
rect -47383 6108 -41168 6172
rect -41104 6108 -41084 6172
rect -47383 6092 -41084 6108
rect -47383 6028 -41168 6092
rect -41104 6028 -41084 6092
rect -47383 6012 -41084 6028
rect -47383 5948 -41168 6012
rect -41104 5948 -41084 6012
rect -47383 5932 -41084 5948
rect -47383 5868 -41168 5932
rect -41104 5868 -41084 5932
rect -47383 5852 -41084 5868
rect -47383 5788 -41168 5852
rect -41104 5788 -41084 5852
rect -47383 5772 -41084 5788
rect -47383 5708 -41168 5772
rect -41104 5708 -41084 5772
rect -47383 5692 -41084 5708
rect -47383 5628 -41168 5692
rect -41104 5628 -41084 5692
rect -47383 5612 -41084 5628
rect -47383 5548 -41168 5612
rect -41104 5548 -41084 5612
rect -47383 5532 -41084 5548
rect -47383 5468 -41168 5532
rect -41104 5468 -41084 5532
rect -47383 5452 -41084 5468
rect -47383 5388 -41168 5452
rect -41104 5388 -41084 5452
rect -47383 5372 -41084 5388
rect -47383 5308 -41168 5372
rect -41104 5308 -41084 5372
rect -47383 5292 -41084 5308
rect -47383 5228 -41168 5292
rect -41104 5228 -41084 5292
rect -47383 5212 -41084 5228
rect -47383 5148 -41168 5212
rect -41104 5148 -41084 5212
rect -47383 5132 -41084 5148
rect -47383 5068 -41168 5132
rect -41104 5068 -41084 5132
rect -47383 5052 -41084 5068
rect -47383 4988 -41168 5052
rect -41104 4988 -41084 5052
rect -47383 4972 -41084 4988
rect -47383 4908 -41168 4972
rect -41104 4908 -41084 4972
rect -47383 4892 -41084 4908
rect -47383 4828 -41168 4892
rect -41104 4828 -41084 4892
rect -47383 4812 -41084 4828
rect -47383 4748 -41168 4812
rect -41104 4748 -41084 4812
rect -47383 4732 -41084 4748
rect -47383 4668 -41168 4732
rect -41104 4668 -41084 4732
rect -47383 4652 -41084 4668
rect -47383 4588 -41168 4652
rect -41104 4588 -41084 4652
rect -47383 4572 -41084 4588
rect -47383 4508 -41168 4572
rect -41104 4508 -41084 4572
rect -47383 4492 -41084 4508
rect -47383 4428 -41168 4492
rect -41104 4428 -41084 4492
rect -47383 4412 -41084 4428
rect -47383 4348 -41168 4412
rect -41104 4348 -41084 4412
rect -47383 4332 -41084 4348
rect -47383 4268 -41168 4332
rect -41104 4268 -41084 4332
rect -47383 4252 -41084 4268
rect -47383 4188 -41168 4252
rect -41104 4188 -41084 4252
rect -47383 4172 -41084 4188
rect -47383 4108 -41168 4172
rect -41104 4108 -41084 4172
rect -47383 4092 -41084 4108
rect -47383 4028 -41168 4092
rect -41104 4028 -41084 4092
rect -47383 4012 -41084 4028
rect -47383 3948 -41168 4012
rect -41104 3948 -41084 4012
rect -47383 3932 -41084 3948
rect -47383 3868 -41168 3932
rect -41104 3868 -41084 3932
rect -47383 3852 -41084 3868
rect -47383 3788 -41168 3852
rect -41104 3788 -41084 3852
rect -47383 3772 -41084 3788
rect -47383 3708 -41168 3772
rect -41104 3708 -41084 3772
rect -47383 3692 -41084 3708
rect -47383 3628 -41168 3692
rect -41104 3628 -41084 3692
rect -47383 3612 -41084 3628
rect -47383 3548 -41168 3612
rect -41104 3548 -41084 3612
rect -47383 3532 -41084 3548
rect -47383 3468 -41168 3532
rect -41104 3468 -41084 3532
rect -47383 3452 -41084 3468
rect -47383 3388 -41168 3452
rect -41104 3388 -41084 3452
rect -47383 3372 -41084 3388
rect -47383 3308 -41168 3372
rect -41104 3308 -41084 3372
rect -47383 3292 -41084 3308
rect -47383 3228 -41168 3292
rect -41104 3228 -41084 3292
rect -47383 3200 -41084 3228
rect -41064 9372 -34765 9400
rect -41064 9308 -34849 9372
rect -34785 9308 -34765 9372
rect -41064 9292 -34765 9308
rect -41064 9228 -34849 9292
rect -34785 9228 -34765 9292
rect -41064 9212 -34765 9228
rect -41064 9148 -34849 9212
rect -34785 9148 -34765 9212
rect -41064 9132 -34765 9148
rect -41064 9068 -34849 9132
rect -34785 9068 -34765 9132
rect -41064 9052 -34765 9068
rect -41064 8988 -34849 9052
rect -34785 8988 -34765 9052
rect -41064 8972 -34765 8988
rect -41064 8908 -34849 8972
rect -34785 8908 -34765 8972
rect -41064 8892 -34765 8908
rect -41064 8828 -34849 8892
rect -34785 8828 -34765 8892
rect -41064 8812 -34765 8828
rect -41064 8748 -34849 8812
rect -34785 8748 -34765 8812
rect -41064 8732 -34765 8748
rect -41064 8668 -34849 8732
rect -34785 8668 -34765 8732
rect -41064 8652 -34765 8668
rect -41064 8588 -34849 8652
rect -34785 8588 -34765 8652
rect -41064 8572 -34765 8588
rect -41064 8508 -34849 8572
rect -34785 8508 -34765 8572
rect -41064 8492 -34765 8508
rect -41064 8428 -34849 8492
rect -34785 8428 -34765 8492
rect -41064 8412 -34765 8428
rect -41064 8348 -34849 8412
rect -34785 8348 -34765 8412
rect -41064 8332 -34765 8348
rect -41064 8268 -34849 8332
rect -34785 8268 -34765 8332
rect -41064 8252 -34765 8268
rect -41064 8188 -34849 8252
rect -34785 8188 -34765 8252
rect -41064 8172 -34765 8188
rect -41064 8108 -34849 8172
rect -34785 8108 -34765 8172
rect -41064 8092 -34765 8108
rect -41064 8028 -34849 8092
rect -34785 8028 -34765 8092
rect -41064 8012 -34765 8028
rect -41064 7948 -34849 8012
rect -34785 7948 -34765 8012
rect -41064 7932 -34765 7948
rect -41064 7868 -34849 7932
rect -34785 7868 -34765 7932
rect -41064 7852 -34765 7868
rect -41064 7788 -34849 7852
rect -34785 7788 -34765 7852
rect -41064 7772 -34765 7788
rect -41064 7708 -34849 7772
rect -34785 7708 -34765 7772
rect -41064 7692 -34765 7708
rect -41064 7628 -34849 7692
rect -34785 7628 -34765 7692
rect -41064 7612 -34765 7628
rect -41064 7548 -34849 7612
rect -34785 7548 -34765 7612
rect -41064 7532 -34765 7548
rect -41064 7468 -34849 7532
rect -34785 7468 -34765 7532
rect -41064 7452 -34765 7468
rect -41064 7388 -34849 7452
rect -34785 7388 -34765 7452
rect -41064 7372 -34765 7388
rect -41064 7308 -34849 7372
rect -34785 7308 -34765 7372
rect -41064 7292 -34765 7308
rect -41064 7228 -34849 7292
rect -34785 7228 -34765 7292
rect -41064 7212 -34765 7228
rect -41064 7148 -34849 7212
rect -34785 7148 -34765 7212
rect -41064 7132 -34765 7148
rect -41064 7068 -34849 7132
rect -34785 7068 -34765 7132
rect -41064 7052 -34765 7068
rect -41064 6988 -34849 7052
rect -34785 6988 -34765 7052
rect -41064 6972 -34765 6988
rect -41064 6908 -34849 6972
rect -34785 6908 -34765 6972
rect -41064 6892 -34765 6908
rect -41064 6828 -34849 6892
rect -34785 6828 -34765 6892
rect -41064 6812 -34765 6828
rect -41064 6748 -34849 6812
rect -34785 6748 -34765 6812
rect -41064 6732 -34765 6748
rect -41064 6668 -34849 6732
rect -34785 6668 -34765 6732
rect -41064 6652 -34765 6668
rect -41064 6588 -34849 6652
rect -34785 6588 -34765 6652
rect -41064 6572 -34765 6588
rect -41064 6508 -34849 6572
rect -34785 6508 -34765 6572
rect -41064 6492 -34765 6508
rect -41064 6428 -34849 6492
rect -34785 6428 -34765 6492
rect -41064 6412 -34765 6428
rect -41064 6348 -34849 6412
rect -34785 6348 -34765 6412
rect -41064 6332 -34765 6348
rect -41064 6268 -34849 6332
rect -34785 6268 -34765 6332
rect -41064 6252 -34765 6268
rect -41064 6188 -34849 6252
rect -34785 6188 -34765 6252
rect -41064 6172 -34765 6188
rect -41064 6108 -34849 6172
rect -34785 6108 -34765 6172
rect -41064 6092 -34765 6108
rect -41064 6028 -34849 6092
rect -34785 6028 -34765 6092
rect -41064 6012 -34765 6028
rect -41064 5948 -34849 6012
rect -34785 5948 -34765 6012
rect -41064 5932 -34765 5948
rect -41064 5868 -34849 5932
rect -34785 5868 -34765 5932
rect -41064 5852 -34765 5868
rect -41064 5788 -34849 5852
rect -34785 5788 -34765 5852
rect -41064 5772 -34765 5788
rect -41064 5708 -34849 5772
rect -34785 5708 -34765 5772
rect -41064 5692 -34765 5708
rect -41064 5628 -34849 5692
rect -34785 5628 -34765 5692
rect -41064 5612 -34765 5628
rect -41064 5548 -34849 5612
rect -34785 5548 -34765 5612
rect -41064 5532 -34765 5548
rect -41064 5468 -34849 5532
rect -34785 5468 -34765 5532
rect -41064 5452 -34765 5468
rect -41064 5388 -34849 5452
rect -34785 5388 -34765 5452
rect -41064 5372 -34765 5388
rect -41064 5308 -34849 5372
rect -34785 5308 -34765 5372
rect -41064 5292 -34765 5308
rect -41064 5228 -34849 5292
rect -34785 5228 -34765 5292
rect -41064 5212 -34765 5228
rect -41064 5148 -34849 5212
rect -34785 5148 -34765 5212
rect -41064 5132 -34765 5148
rect -41064 5068 -34849 5132
rect -34785 5068 -34765 5132
rect -41064 5052 -34765 5068
rect -41064 4988 -34849 5052
rect -34785 4988 -34765 5052
rect -41064 4972 -34765 4988
rect -41064 4908 -34849 4972
rect -34785 4908 -34765 4972
rect -41064 4892 -34765 4908
rect -41064 4828 -34849 4892
rect -34785 4828 -34765 4892
rect -41064 4812 -34765 4828
rect -41064 4748 -34849 4812
rect -34785 4748 -34765 4812
rect -41064 4732 -34765 4748
rect -41064 4668 -34849 4732
rect -34785 4668 -34765 4732
rect -41064 4652 -34765 4668
rect -41064 4588 -34849 4652
rect -34785 4588 -34765 4652
rect -41064 4572 -34765 4588
rect -41064 4508 -34849 4572
rect -34785 4508 -34765 4572
rect -41064 4492 -34765 4508
rect -41064 4428 -34849 4492
rect -34785 4428 -34765 4492
rect -41064 4412 -34765 4428
rect -41064 4348 -34849 4412
rect -34785 4348 -34765 4412
rect -41064 4332 -34765 4348
rect -41064 4268 -34849 4332
rect -34785 4268 -34765 4332
rect -41064 4252 -34765 4268
rect -41064 4188 -34849 4252
rect -34785 4188 -34765 4252
rect -41064 4172 -34765 4188
rect -41064 4108 -34849 4172
rect -34785 4108 -34765 4172
rect -41064 4092 -34765 4108
rect -41064 4028 -34849 4092
rect -34785 4028 -34765 4092
rect -41064 4012 -34765 4028
rect -41064 3948 -34849 4012
rect -34785 3948 -34765 4012
rect -41064 3932 -34765 3948
rect -41064 3868 -34849 3932
rect -34785 3868 -34765 3932
rect -41064 3852 -34765 3868
rect -41064 3788 -34849 3852
rect -34785 3788 -34765 3852
rect -41064 3772 -34765 3788
rect -41064 3708 -34849 3772
rect -34785 3708 -34765 3772
rect -41064 3692 -34765 3708
rect -41064 3628 -34849 3692
rect -34785 3628 -34765 3692
rect -41064 3612 -34765 3628
rect -41064 3548 -34849 3612
rect -34785 3548 -34765 3612
rect -41064 3532 -34765 3548
rect -41064 3468 -34849 3532
rect -34785 3468 -34765 3532
rect -41064 3452 -34765 3468
rect -41064 3388 -34849 3452
rect -34785 3388 -34765 3452
rect -41064 3372 -34765 3388
rect -41064 3308 -34849 3372
rect -34785 3308 -34765 3372
rect -41064 3292 -34765 3308
rect -41064 3228 -34849 3292
rect -34785 3228 -34765 3292
rect -41064 3200 -34765 3228
rect -34745 9372 -28446 9400
rect -34745 9308 -28530 9372
rect -28466 9308 -28446 9372
rect -34745 9292 -28446 9308
rect -34745 9228 -28530 9292
rect -28466 9228 -28446 9292
rect -34745 9212 -28446 9228
rect -34745 9148 -28530 9212
rect -28466 9148 -28446 9212
rect -34745 9132 -28446 9148
rect -34745 9068 -28530 9132
rect -28466 9068 -28446 9132
rect -34745 9052 -28446 9068
rect -34745 8988 -28530 9052
rect -28466 8988 -28446 9052
rect -34745 8972 -28446 8988
rect -34745 8908 -28530 8972
rect -28466 8908 -28446 8972
rect -34745 8892 -28446 8908
rect -34745 8828 -28530 8892
rect -28466 8828 -28446 8892
rect -34745 8812 -28446 8828
rect -34745 8748 -28530 8812
rect -28466 8748 -28446 8812
rect -34745 8732 -28446 8748
rect -34745 8668 -28530 8732
rect -28466 8668 -28446 8732
rect -34745 8652 -28446 8668
rect -34745 8588 -28530 8652
rect -28466 8588 -28446 8652
rect -34745 8572 -28446 8588
rect -34745 8508 -28530 8572
rect -28466 8508 -28446 8572
rect -34745 8492 -28446 8508
rect -34745 8428 -28530 8492
rect -28466 8428 -28446 8492
rect -34745 8412 -28446 8428
rect -34745 8348 -28530 8412
rect -28466 8348 -28446 8412
rect -34745 8332 -28446 8348
rect -34745 8268 -28530 8332
rect -28466 8268 -28446 8332
rect -34745 8252 -28446 8268
rect -34745 8188 -28530 8252
rect -28466 8188 -28446 8252
rect -34745 8172 -28446 8188
rect -34745 8108 -28530 8172
rect -28466 8108 -28446 8172
rect -34745 8092 -28446 8108
rect -34745 8028 -28530 8092
rect -28466 8028 -28446 8092
rect -34745 8012 -28446 8028
rect -34745 7948 -28530 8012
rect -28466 7948 -28446 8012
rect -34745 7932 -28446 7948
rect -34745 7868 -28530 7932
rect -28466 7868 -28446 7932
rect -34745 7852 -28446 7868
rect -34745 7788 -28530 7852
rect -28466 7788 -28446 7852
rect -34745 7772 -28446 7788
rect -34745 7708 -28530 7772
rect -28466 7708 -28446 7772
rect -34745 7692 -28446 7708
rect -34745 7628 -28530 7692
rect -28466 7628 -28446 7692
rect -34745 7612 -28446 7628
rect -34745 7548 -28530 7612
rect -28466 7548 -28446 7612
rect -34745 7532 -28446 7548
rect -34745 7468 -28530 7532
rect -28466 7468 -28446 7532
rect -34745 7452 -28446 7468
rect -34745 7388 -28530 7452
rect -28466 7388 -28446 7452
rect -34745 7372 -28446 7388
rect -34745 7308 -28530 7372
rect -28466 7308 -28446 7372
rect -34745 7292 -28446 7308
rect -34745 7228 -28530 7292
rect -28466 7228 -28446 7292
rect -34745 7212 -28446 7228
rect -34745 7148 -28530 7212
rect -28466 7148 -28446 7212
rect -34745 7132 -28446 7148
rect -34745 7068 -28530 7132
rect -28466 7068 -28446 7132
rect -34745 7052 -28446 7068
rect -34745 6988 -28530 7052
rect -28466 6988 -28446 7052
rect -34745 6972 -28446 6988
rect -34745 6908 -28530 6972
rect -28466 6908 -28446 6972
rect -34745 6892 -28446 6908
rect -34745 6828 -28530 6892
rect -28466 6828 -28446 6892
rect -34745 6812 -28446 6828
rect -34745 6748 -28530 6812
rect -28466 6748 -28446 6812
rect -34745 6732 -28446 6748
rect -34745 6668 -28530 6732
rect -28466 6668 -28446 6732
rect -34745 6652 -28446 6668
rect -34745 6588 -28530 6652
rect -28466 6588 -28446 6652
rect -34745 6572 -28446 6588
rect -34745 6508 -28530 6572
rect -28466 6508 -28446 6572
rect -34745 6492 -28446 6508
rect -34745 6428 -28530 6492
rect -28466 6428 -28446 6492
rect -34745 6412 -28446 6428
rect -34745 6348 -28530 6412
rect -28466 6348 -28446 6412
rect -34745 6332 -28446 6348
rect -34745 6268 -28530 6332
rect -28466 6268 -28446 6332
rect -34745 6252 -28446 6268
rect -34745 6188 -28530 6252
rect -28466 6188 -28446 6252
rect -34745 6172 -28446 6188
rect -34745 6108 -28530 6172
rect -28466 6108 -28446 6172
rect -34745 6092 -28446 6108
rect -34745 6028 -28530 6092
rect -28466 6028 -28446 6092
rect -34745 6012 -28446 6028
rect -34745 5948 -28530 6012
rect -28466 5948 -28446 6012
rect -34745 5932 -28446 5948
rect -34745 5868 -28530 5932
rect -28466 5868 -28446 5932
rect -34745 5852 -28446 5868
rect -34745 5788 -28530 5852
rect -28466 5788 -28446 5852
rect -34745 5772 -28446 5788
rect -34745 5708 -28530 5772
rect -28466 5708 -28446 5772
rect -34745 5692 -28446 5708
rect -34745 5628 -28530 5692
rect -28466 5628 -28446 5692
rect -34745 5612 -28446 5628
rect -34745 5548 -28530 5612
rect -28466 5548 -28446 5612
rect -34745 5532 -28446 5548
rect -34745 5468 -28530 5532
rect -28466 5468 -28446 5532
rect -34745 5452 -28446 5468
rect -34745 5388 -28530 5452
rect -28466 5388 -28446 5452
rect -34745 5372 -28446 5388
rect -34745 5308 -28530 5372
rect -28466 5308 -28446 5372
rect -34745 5292 -28446 5308
rect -34745 5228 -28530 5292
rect -28466 5228 -28446 5292
rect -34745 5212 -28446 5228
rect -34745 5148 -28530 5212
rect -28466 5148 -28446 5212
rect -34745 5132 -28446 5148
rect -34745 5068 -28530 5132
rect -28466 5068 -28446 5132
rect -34745 5052 -28446 5068
rect -34745 4988 -28530 5052
rect -28466 4988 -28446 5052
rect -34745 4972 -28446 4988
rect -34745 4908 -28530 4972
rect -28466 4908 -28446 4972
rect -34745 4892 -28446 4908
rect -34745 4828 -28530 4892
rect -28466 4828 -28446 4892
rect -34745 4812 -28446 4828
rect -34745 4748 -28530 4812
rect -28466 4748 -28446 4812
rect -34745 4732 -28446 4748
rect -34745 4668 -28530 4732
rect -28466 4668 -28446 4732
rect -34745 4652 -28446 4668
rect -34745 4588 -28530 4652
rect -28466 4588 -28446 4652
rect -34745 4572 -28446 4588
rect -34745 4508 -28530 4572
rect -28466 4508 -28446 4572
rect -34745 4492 -28446 4508
rect -34745 4428 -28530 4492
rect -28466 4428 -28446 4492
rect -34745 4412 -28446 4428
rect -34745 4348 -28530 4412
rect -28466 4348 -28446 4412
rect -34745 4332 -28446 4348
rect -34745 4268 -28530 4332
rect -28466 4268 -28446 4332
rect -34745 4252 -28446 4268
rect -34745 4188 -28530 4252
rect -28466 4188 -28446 4252
rect -34745 4172 -28446 4188
rect -34745 4108 -28530 4172
rect -28466 4108 -28446 4172
rect -34745 4092 -28446 4108
rect -34745 4028 -28530 4092
rect -28466 4028 -28446 4092
rect -34745 4012 -28446 4028
rect -34745 3948 -28530 4012
rect -28466 3948 -28446 4012
rect -34745 3932 -28446 3948
rect -34745 3868 -28530 3932
rect -28466 3868 -28446 3932
rect -34745 3852 -28446 3868
rect -34745 3788 -28530 3852
rect -28466 3788 -28446 3852
rect -34745 3772 -28446 3788
rect -34745 3708 -28530 3772
rect -28466 3708 -28446 3772
rect -34745 3692 -28446 3708
rect -34745 3628 -28530 3692
rect -28466 3628 -28446 3692
rect -34745 3612 -28446 3628
rect -34745 3548 -28530 3612
rect -28466 3548 -28446 3612
rect -34745 3532 -28446 3548
rect -34745 3468 -28530 3532
rect -28466 3468 -28446 3532
rect -34745 3452 -28446 3468
rect -34745 3388 -28530 3452
rect -28466 3388 -28446 3452
rect -34745 3372 -28446 3388
rect -34745 3308 -28530 3372
rect -28466 3308 -28446 3372
rect -34745 3292 -28446 3308
rect -34745 3228 -28530 3292
rect -28466 3228 -28446 3292
rect -34745 3200 -28446 3228
rect -28426 9372 -22127 9400
rect -28426 9308 -22211 9372
rect -22147 9308 -22127 9372
rect -28426 9292 -22127 9308
rect -28426 9228 -22211 9292
rect -22147 9228 -22127 9292
rect -28426 9212 -22127 9228
rect -28426 9148 -22211 9212
rect -22147 9148 -22127 9212
rect -28426 9132 -22127 9148
rect -28426 9068 -22211 9132
rect -22147 9068 -22127 9132
rect -28426 9052 -22127 9068
rect -28426 8988 -22211 9052
rect -22147 8988 -22127 9052
rect -28426 8972 -22127 8988
rect -28426 8908 -22211 8972
rect -22147 8908 -22127 8972
rect -28426 8892 -22127 8908
rect -28426 8828 -22211 8892
rect -22147 8828 -22127 8892
rect -28426 8812 -22127 8828
rect -28426 8748 -22211 8812
rect -22147 8748 -22127 8812
rect -28426 8732 -22127 8748
rect -28426 8668 -22211 8732
rect -22147 8668 -22127 8732
rect -28426 8652 -22127 8668
rect -28426 8588 -22211 8652
rect -22147 8588 -22127 8652
rect -28426 8572 -22127 8588
rect -28426 8508 -22211 8572
rect -22147 8508 -22127 8572
rect -28426 8492 -22127 8508
rect -28426 8428 -22211 8492
rect -22147 8428 -22127 8492
rect -28426 8412 -22127 8428
rect -28426 8348 -22211 8412
rect -22147 8348 -22127 8412
rect -28426 8332 -22127 8348
rect -28426 8268 -22211 8332
rect -22147 8268 -22127 8332
rect -28426 8252 -22127 8268
rect -28426 8188 -22211 8252
rect -22147 8188 -22127 8252
rect -28426 8172 -22127 8188
rect -28426 8108 -22211 8172
rect -22147 8108 -22127 8172
rect -28426 8092 -22127 8108
rect -28426 8028 -22211 8092
rect -22147 8028 -22127 8092
rect -28426 8012 -22127 8028
rect -28426 7948 -22211 8012
rect -22147 7948 -22127 8012
rect -28426 7932 -22127 7948
rect -28426 7868 -22211 7932
rect -22147 7868 -22127 7932
rect -28426 7852 -22127 7868
rect -28426 7788 -22211 7852
rect -22147 7788 -22127 7852
rect -28426 7772 -22127 7788
rect -28426 7708 -22211 7772
rect -22147 7708 -22127 7772
rect -28426 7692 -22127 7708
rect -28426 7628 -22211 7692
rect -22147 7628 -22127 7692
rect -28426 7612 -22127 7628
rect -28426 7548 -22211 7612
rect -22147 7548 -22127 7612
rect -28426 7532 -22127 7548
rect -28426 7468 -22211 7532
rect -22147 7468 -22127 7532
rect -28426 7452 -22127 7468
rect -28426 7388 -22211 7452
rect -22147 7388 -22127 7452
rect -28426 7372 -22127 7388
rect -28426 7308 -22211 7372
rect -22147 7308 -22127 7372
rect -28426 7292 -22127 7308
rect -28426 7228 -22211 7292
rect -22147 7228 -22127 7292
rect -28426 7212 -22127 7228
rect -28426 7148 -22211 7212
rect -22147 7148 -22127 7212
rect -28426 7132 -22127 7148
rect -28426 7068 -22211 7132
rect -22147 7068 -22127 7132
rect -28426 7052 -22127 7068
rect -28426 6988 -22211 7052
rect -22147 6988 -22127 7052
rect -28426 6972 -22127 6988
rect -28426 6908 -22211 6972
rect -22147 6908 -22127 6972
rect -28426 6892 -22127 6908
rect -28426 6828 -22211 6892
rect -22147 6828 -22127 6892
rect -28426 6812 -22127 6828
rect -28426 6748 -22211 6812
rect -22147 6748 -22127 6812
rect -28426 6732 -22127 6748
rect -28426 6668 -22211 6732
rect -22147 6668 -22127 6732
rect -28426 6652 -22127 6668
rect -28426 6588 -22211 6652
rect -22147 6588 -22127 6652
rect -28426 6572 -22127 6588
rect -28426 6508 -22211 6572
rect -22147 6508 -22127 6572
rect -28426 6492 -22127 6508
rect -28426 6428 -22211 6492
rect -22147 6428 -22127 6492
rect -28426 6412 -22127 6428
rect -28426 6348 -22211 6412
rect -22147 6348 -22127 6412
rect -28426 6332 -22127 6348
rect -28426 6268 -22211 6332
rect -22147 6268 -22127 6332
rect -28426 6252 -22127 6268
rect -28426 6188 -22211 6252
rect -22147 6188 -22127 6252
rect -28426 6172 -22127 6188
rect -28426 6108 -22211 6172
rect -22147 6108 -22127 6172
rect -28426 6092 -22127 6108
rect -28426 6028 -22211 6092
rect -22147 6028 -22127 6092
rect -28426 6012 -22127 6028
rect -28426 5948 -22211 6012
rect -22147 5948 -22127 6012
rect -28426 5932 -22127 5948
rect -28426 5868 -22211 5932
rect -22147 5868 -22127 5932
rect -28426 5852 -22127 5868
rect -28426 5788 -22211 5852
rect -22147 5788 -22127 5852
rect -28426 5772 -22127 5788
rect -28426 5708 -22211 5772
rect -22147 5708 -22127 5772
rect -28426 5692 -22127 5708
rect -28426 5628 -22211 5692
rect -22147 5628 -22127 5692
rect -28426 5612 -22127 5628
rect -28426 5548 -22211 5612
rect -22147 5548 -22127 5612
rect -28426 5532 -22127 5548
rect -28426 5468 -22211 5532
rect -22147 5468 -22127 5532
rect -28426 5452 -22127 5468
rect -28426 5388 -22211 5452
rect -22147 5388 -22127 5452
rect -28426 5372 -22127 5388
rect -28426 5308 -22211 5372
rect -22147 5308 -22127 5372
rect -28426 5292 -22127 5308
rect -28426 5228 -22211 5292
rect -22147 5228 -22127 5292
rect -28426 5212 -22127 5228
rect -28426 5148 -22211 5212
rect -22147 5148 -22127 5212
rect -28426 5132 -22127 5148
rect -28426 5068 -22211 5132
rect -22147 5068 -22127 5132
rect -28426 5052 -22127 5068
rect -28426 4988 -22211 5052
rect -22147 4988 -22127 5052
rect -28426 4972 -22127 4988
rect -28426 4908 -22211 4972
rect -22147 4908 -22127 4972
rect -28426 4892 -22127 4908
rect -28426 4828 -22211 4892
rect -22147 4828 -22127 4892
rect -28426 4812 -22127 4828
rect -28426 4748 -22211 4812
rect -22147 4748 -22127 4812
rect -28426 4732 -22127 4748
rect -28426 4668 -22211 4732
rect -22147 4668 -22127 4732
rect -28426 4652 -22127 4668
rect -28426 4588 -22211 4652
rect -22147 4588 -22127 4652
rect -28426 4572 -22127 4588
rect -28426 4508 -22211 4572
rect -22147 4508 -22127 4572
rect -28426 4492 -22127 4508
rect -28426 4428 -22211 4492
rect -22147 4428 -22127 4492
rect -28426 4412 -22127 4428
rect -28426 4348 -22211 4412
rect -22147 4348 -22127 4412
rect -28426 4332 -22127 4348
rect -28426 4268 -22211 4332
rect -22147 4268 -22127 4332
rect -28426 4252 -22127 4268
rect -28426 4188 -22211 4252
rect -22147 4188 -22127 4252
rect -28426 4172 -22127 4188
rect -28426 4108 -22211 4172
rect -22147 4108 -22127 4172
rect -28426 4092 -22127 4108
rect -28426 4028 -22211 4092
rect -22147 4028 -22127 4092
rect -28426 4012 -22127 4028
rect -28426 3948 -22211 4012
rect -22147 3948 -22127 4012
rect -28426 3932 -22127 3948
rect -28426 3868 -22211 3932
rect -22147 3868 -22127 3932
rect -28426 3852 -22127 3868
rect -28426 3788 -22211 3852
rect -22147 3788 -22127 3852
rect -28426 3772 -22127 3788
rect -28426 3708 -22211 3772
rect -22147 3708 -22127 3772
rect -28426 3692 -22127 3708
rect -28426 3628 -22211 3692
rect -22147 3628 -22127 3692
rect -28426 3612 -22127 3628
rect -28426 3548 -22211 3612
rect -22147 3548 -22127 3612
rect -28426 3532 -22127 3548
rect -28426 3468 -22211 3532
rect -22147 3468 -22127 3532
rect -28426 3452 -22127 3468
rect -28426 3388 -22211 3452
rect -22147 3388 -22127 3452
rect -28426 3372 -22127 3388
rect -28426 3308 -22211 3372
rect -22147 3308 -22127 3372
rect -28426 3292 -22127 3308
rect -28426 3228 -22211 3292
rect -22147 3228 -22127 3292
rect -28426 3200 -22127 3228
rect -22107 9372 -15808 9400
rect -22107 9308 -15892 9372
rect -15828 9308 -15808 9372
rect -22107 9292 -15808 9308
rect -22107 9228 -15892 9292
rect -15828 9228 -15808 9292
rect -22107 9212 -15808 9228
rect -22107 9148 -15892 9212
rect -15828 9148 -15808 9212
rect -22107 9132 -15808 9148
rect -22107 9068 -15892 9132
rect -15828 9068 -15808 9132
rect -22107 9052 -15808 9068
rect -22107 8988 -15892 9052
rect -15828 8988 -15808 9052
rect -22107 8972 -15808 8988
rect -22107 8908 -15892 8972
rect -15828 8908 -15808 8972
rect -22107 8892 -15808 8908
rect -22107 8828 -15892 8892
rect -15828 8828 -15808 8892
rect -22107 8812 -15808 8828
rect -22107 8748 -15892 8812
rect -15828 8748 -15808 8812
rect -22107 8732 -15808 8748
rect -22107 8668 -15892 8732
rect -15828 8668 -15808 8732
rect -22107 8652 -15808 8668
rect -22107 8588 -15892 8652
rect -15828 8588 -15808 8652
rect -22107 8572 -15808 8588
rect -22107 8508 -15892 8572
rect -15828 8508 -15808 8572
rect -22107 8492 -15808 8508
rect -22107 8428 -15892 8492
rect -15828 8428 -15808 8492
rect -22107 8412 -15808 8428
rect -22107 8348 -15892 8412
rect -15828 8348 -15808 8412
rect -22107 8332 -15808 8348
rect -22107 8268 -15892 8332
rect -15828 8268 -15808 8332
rect -22107 8252 -15808 8268
rect -22107 8188 -15892 8252
rect -15828 8188 -15808 8252
rect -22107 8172 -15808 8188
rect -22107 8108 -15892 8172
rect -15828 8108 -15808 8172
rect -22107 8092 -15808 8108
rect -22107 8028 -15892 8092
rect -15828 8028 -15808 8092
rect -22107 8012 -15808 8028
rect -22107 7948 -15892 8012
rect -15828 7948 -15808 8012
rect -22107 7932 -15808 7948
rect -22107 7868 -15892 7932
rect -15828 7868 -15808 7932
rect -22107 7852 -15808 7868
rect -22107 7788 -15892 7852
rect -15828 7788 -15808 7852
rect -22107 7772 -15808 7788
rect -22107 7708 -15892 7772
rect -15828 7708 -15808 7772
rect -22107 7692 -15808 7708
rect -22107 7628 -15892 7692
rect -15828 7628 -15808 7692
rect -22107 7612 -15808 7628
rect -22107 7548 -15892 7612
rect -15828 7548 -15808 7612
rect -22107 7532 -15808 7548
rect -22107 7468 -15892 7532
rect -15828 7468 -15808 7532
rect -22107 7452 -15808 7468
rect -22107 7388 -15892 7452
rect -15828 7388 -15808 7452
rect -22107 7372 -15808 7388
rect -22107 7308 -15892 7372
rect -15828 7308 -15808 7372
rect -22107 7292 -15808 7308
rect -22107 7228 -15892 7292
rect -15828 7228 -15808 7292
rect -22107 7212 -15808 7228
rect -22107 7148 -15892 7212
rect -15828 7148 -15808 7212
rect -22107 7132 -15808 7148
rect -22107 7068 -15892 7132
rect -15828 7068 -15808 7132
rect -22107 7052 -15808 7068
rect -22107 6988 -15892 7052
rect -15828 6988 -15808 7052
rect -22107 6972 -15808 6988
rect -22107 6908 -15892 6972
rect -15828 6908 -15808 6972
rect -22107 6892 -15808 6908
rect -22107 6828 -15892 6892
rect -15828 6828 -15808 6892
rect -22107 6812 -15808 6828
rect -22107 6748 -15892 6812
rect -15828 6748 -15808 6812
rect -22107 6732 -15808 6748
rect -22107 6668 -15892 6732
rect -15828 6668 -15808 6732
rect -22107 6652 -15808 6668
rect -22107 6588 -15892 6652
rect -15828 6588 -15808 6652
rect -22107 6572 -15808 6588
rect -22107 6508 -15892 6572
rect -15828 6508 -15808 6572
rect -22107 6492 -15808 6508
rect -22107 6428 -15892 6492
rect -15828 6428 -15808 6492
rect -22107 6412 -15808 6428
rect -22107 6348 -15892 6412
rect -15828 6348 -15808 6412
rect -22107 6332 -15808 6348
rect -22107 6268 -15892 6332
rect -15828 6268 -15808 6332
rect -22107 6252 -15808 6268
rect -22107 6188 -15892 6252
rect -15828 6188 -15808 6252
rect -22107 6172 -15808 6188
rect -22107 6108 -15892 6172
rect -15828 6108 -15808 6172
rect -22107 6092 -15808 6108
rect -22107 6028 -15892 6092
rect -15828 6028 -15808 6092
rect -22107 6012 -15808 6028
rect -22107 5948 -15892 6012
rect -15828 5948 -15808 6012
rect -22107 5932 -15808 5948
rect -22107 5868 -15892 5932
rect -15828 5868 -15808 5932
rect -22107 5852 -15808 5868
rect -22107 5788 -15892 5852
rect -15828 5788 -15808 5852
rect -22107 5772 -15808 5788
rect -22107 5708 -15892 5772
rect -15828 5708 -15808 5772
rect -22107 5692 -15808 5708
rect -22107 5628 -15892 5692
rect -15828 5628 -15808 5692
rect -22107 5612 -15808 5628
rect -22107 5548 -15892 5612
rect -15828 5548 -15808 5612
rect -22107 5532 -15808 5548
rect -22107 5468 -15892 5532
rect -15828 5468 -15808 5532
rect -22107 5452 -15808 5468
rect -22107 5388 -15892 5452
rect -15828 5388 -15808 5452
rect -22107 5372 -15808 5388
rect -22107 5308 -15892 5372
rect -15828 5308 -15808 5372
rect -22107 5292 -15808 5308
rect -22107 5228 -15892 5292
rect -15828 5228 -15808 5292
rect -22107 5212 -15808 5228
rect -22107 5148 -15892 5212
rect -15828 5148 -15808 5212
rect -22107 5132 -15808 5148
rect -22107 5068 -15892 5132
rect -15828 5068 -15808 5132
rect -22107 5052 -15808 5068
rect -22107 4988 -15892 5052
rect -15828 4988 -15808 5052
rect -22107 4972 -15808 4988
rect -22107 4908 -15892 4972
rect -15828 4908 -15808 4972
rect -22107 4892 -15808 4908
rect -22107 4828 -15892 4892
rect -15828 4828 -15808 4892
rect -22107 4812 -15808 4828
rect -22107 4748 -15892 4812
rect -15828 4748 -15808 4812
rect -22107 4732 -15808 4748
rect -22107 4668 -15892 4732
rect -15828 4668 -15808 4732
rect -22107 4652 -15808 4668
rect -22107 4588 -15892 4652
rect -15828 4588 -15808 4652
rect -22107 4572 -15808 4588
rect -22107 4508 -15892 4572
rect -15828 4508 -15808 4572
rect -22107 4492 -15808 4508
rect -22107 4428 -15892 4492
rect -15828 4428 -15808 4492
rect -22107 4412 -15808 4428
rect -22107 4348 -15892 4412
rect -15828 4348 -15808 4412
rect -22107 4332 -15808 4348
rect -22107 4268 -15892 4332
rect -15828 4268 -15808 4332
rect -22107 4252 -15808 4268
rect -22107 4188 -15892 4252
rect -15828 4188 -15808 4252
rect -22107 4172 -15808 4188
rect -22107 4108 -15892 4172
rect -15828 4108 -15808 4172
rect -22107 4092 -15808 4108
rect -22107 4028 -15892 4092
rect -15828 4028 -15808 4092
rect -22107 4012 -15808 4028
rect -22107 3948 -15892 4012
rect -15828 3948 -15808 4012
rect -22107 3932 -15808 3948
rect -22107 3868 -15892 3932
rect -15828 3868 -15808 3932
rect -22107 3852 -15808 3868
rect -22107 3788 -15892 3852
rect -15828 3788 -15808 3852
rect -22107 3772 -15808 3788
rect -22107 3708 -15892 3772
rect -15828 3708 -15808 3772
rect -22107 3692 -15808 3708
rect -22107 3628 -15892 3692
rect -15828 3628 -15808 3692
rect -22107 3612 -15808 3628
rect -22107 3548 -15892 3612
rect -15828 3548 -15808 3612
rect -22107 3532 -15808 3548
rect -22107 3468 -15892 3532
rect -15828 3468 -15808 3532
rect -22107 3452 -15808 3468
rect -22107 3388 -15892 3452
rect -15828 3388 -15808 3452
rect -22107 3372 -15808 3388
rect -22107 3308 -15892 3372
rect -15828 3308 -15808 3372
rect -22107 3292 -15808 3308
rect -22107 3228 -15892 3292
rect -15828 3228 -15808 3292
rect -22107 3200 -15808 3228
rect -15788 9372 -9489 9400
rect -15788 9308 -9573 9372
rect -9509 9308 -9489 9372
rect -15788 9292 -9489 9308
rect -15788 9228 -9573 9292
rect -9509 9228 -9489 9292
rect -15788 9212 -9489 9228
rect -15788 9148 -9573 9212
rect -9509 9148 -9489 9212
rect -15788 9132 -9489 9148
rect -15788 9068 -9573 9132
rect -9509 9068 -9489 9132
rect -15788 9052 -9489 9068
rect -15788 8988 -9573 9052
rect -9509 8988 -9489 9052
rect -15788 8972 -9489 8988
rect -15788 8908 -9573 8972
rect -9509 8908 -9489 8972
rect -15788 8892 -9489 8908
rect -15788 8828 -9573 8892
rect -9509 8828 -9489 8892
rect -15788 8812 -9489 8828
rect -15788 8748 -9573 8812
rect -9509 8748 -9489 8812
rect -15788 8732 -9489 8748
rect -15788 8668 -9573 8732
rect -9509 8668 -9489 8732
rect -15788 8652 -9489 8668
rect -15788 8588 -9573 8652
rect -9509 8588 -9489 8652
rect -15788 8572 -9489 8588
rect -15788 8508 -9573 8572
rect -9509 8508 -9489 8572
rect -15788 8492 -9489 8508
rect -15788 8428 -9573 8492
rect -9509 8428 -9489 8492
rect -15788 8412 -9489 8428
rect -15788 8348 -9573 8412
rect -9509 8348 -9489 8412
rect -15788 8332 -9489 8348
rect -15788 8268 -9573 8332
rect -9509 8268 -9489 8332
rect -15788 8252 -9489 8268
rect -15788 8188 -9573 8252
rect -9509 8188 -9489 8252
rect -15788 8172 -9489 8188
rect -15788 8108 -9573 8172
rect -9509 8108 -9489 8172
rect -15788 8092 -9489 8108
rect -15788 8028 -9573 8092
rect -9509 8028 -9489 8092
rect -15788 8012 -9489 8028
rect -15788 7948 -9573 8012
rect -9509 7948 -9489 8012
rect -15788 7932 -9489 7948
rect -15788 7868 -9573 7932
rect -9509 7868 -9489 7932
rect -15788 7852 -9489 7868
rect -15788 7788 -9573 7852
rect -9509 7788 -9489 7852
rect -15788 7772 -9489 7788
rect -15788 7708 -9573 7772
rect -9509 7708 -9489 7772
rect -15788 7692 -9489 7708
rect -15788 7628 -9573 7692
rect -9509 7628 -9489 7692
rect -15788 7612 -9489 7628
rect -15788 7548 -9573 7612
rect -9509 7548 -9489 7612
rect -15788 7532 -9489 7548
rect -15788 7468 -9573 7532
rect -9509 7468 -9489 7532
rect -15788 7452 -9489 7468
rect -15788 7388 -9573 7452
rect -9509 7388 -9489 7452
rect -15788 7372 -9489 7388
rect -15788 7308 -9573 7372
rect -9509 7308 -9489 7372
rect -15788 7292 -9489 7308
rect -15788 7228 -9573 7292
rect -9509 7228 -9489 7292
rect -15788 7212 -9489 7228
rect -15788 7148 -9573 7212
rect -9509 7148 -9489 7212
rect -15788 7132 -9489 7148
rect -15788 7068 -9573 7132
rect -9509 7068 -9489 7132
rect -15788 7052 -9489 7068
rect -15788 6988 -9573 7052
rect -9509 6988 -9489 7052
rect -15788 6972 -9489 6988
rect -15788 6908 -9573 6972
rect -9509 6908 -9489 6972
rect -15788 6892 -9489 6908
rect -15788 6828 -9573 6892
rect -9509 6828 -9489 6892
rect -15788 6812 -9489 6828
rect -15788 6748 -9573 6812
rect -9509 6748 -9489 6812
rect -15788 6732 -9489 6748
rect -15788 6668 -9573 6732
rect -9509 6668 -9489 6732
rect -15788 6652 -9489 6668
rect -15788 6588 -9573 6652
rect -9509 6588 -9489 6652
rect -15788 6572 -9489 6588
rect -15788 6508 -9573 6572
rect -9509 6508 -9489 6572
rect -15788 6492 -9489 6508
rect -15788 6428 -9573 6492
rect -9509 6428 -9489 6492
rect -15788 6412 -9489 6428
rect -15788 6348 -9573 6412
rect -9509 6348 -9489 6412
rect -15788 6332 -9489 6348
rect -15788 6268 -9573 6332
rect -9509 6268 -9489 6332
rect -15788 6252 -9489 6268
rect -15788 6188 -9573 6252
rect -9509 6188 -9489 6252
rect -15788 6172 -9489 6188
rect -15788 6108 -9573 6172
rect -9509 6108 -9489 6172
rect -15788 6092 -9489 6108
rect -15788 6028 -9573 6092
rect -9509 6028 -9489 6092
rect -15788 6012 -9489 6028
rect -15788 5948 -9573 6012
rect -9509 5948 -9489 6012
rect -15788 5932 -9489 5948
rect -15788 5868 -9573 5932
rect -9509 5868 -9489 5932
rect -15788 5852 -9489 5868
rect -15788 5788 -9573 5852
rect -9509 5788 -9489 5852
rect -15788 5772 -9489 5788
rect -15788 5708 -9573 5772
rect -9509 5708 -9489 5772
rect -15788 5692 -9489 5708
rect -15788 5628 -9573 5692
rect -9509 5628 -9489 5692
rect -15788 5612 -9489 5628
rect -15788 5548 -9573 5612
rect -9509 5548 -9489 5612
rect -15788 5532 -9489 5548
rect -15788 5468 -9573 5532
rect -9509 5468 -9489 5532
rect -15788 5452 -9489 5468
rect -15788 5388 -9573 5452
rect -9509 5388 -9489 5452
rect -15788 5372 -9489 5388
rect -15788 5308 -9573 5372
rect -9509 5308 -9489 5372
rect -15788 5292 -9489 5308
rect -15788 5228 -9573 5292
rect -9509 5228 -9489 5292
rect -15788 5212 -9489 5228
rect -15788 5148 -9573 5212
rect -9509 5148 -9489 5212
rect -15788 5132 -9489 5148
rect -15788 5068 -9573 5132
rect -9509 5068 -9489 5132
rect -15788 5052 -9489 5068
rect -15788 4988 -9573 5052
rect -9509 4988 -9489 5052
rect -15788 4972 -9489 4988
rect -15788 4908 -9573 4972
rect -9509 4908 -9489 4972
rect -15788 4892 -9489 4908
rect -15788 4828 -9573 4892
rect -9509 4828 -9489 4892
rect -15788 4812 -9489 4828
rect -15788 4748 -9573 4812
rect -9509 4748 -9489 4812
rect -15788 4732 -9489 4748
rect -15788 4668 -9573 4732
rect -9509 4668 -9489 4732
rect -15788 4652 -9489 4668
rect -15788 4588 -9573 4652
rect -9509 4588 -9489 4652
rect -15788 4572 -9489 4588
rect -15788 4508 -9573 4572
rect -9509 4508 -9489 4572
rect -15788 4492 -9489 4508
rect -15788 4428 -9573 4492
rect -9509 4428 -9489 4492
rect -15788 4412 -9489 4428
rect -15788 4348 -9573 4412
rect -9509 4348 -9489 4412
rect -15788 4332 -9489 4348
rect -15788 4268 -9573 4332
rect -9509 4268 -9489 4332
rect -15788 4252 -9489 4268
rect -15788 4188 -9573 4252
rect -9509 4188 -9489 4252
rect -15788 4172 -9489 4188
rect -15788 4108 -9573 4172
rect -9509 4108 -9489 4172
rect -15788 4092 -9489 4108
rect -15788 4028 -9573 4092
rect -9509 4028 -9489 4092
rect -15788 4012 -9489 4028
rect -15788 3948 -9573 4012
rect -9509 3948 -9489 4012
rect -15788 3932 -9489 3948
rect -15788 3868 -9573 3932
rect -9509 3868 -9489 3932
rect -15788 3852 -9489 3868
rect -15788 3788 -9573 3852
rect -9509 3788 -9489 3852
rect -15788 3772 -9489 3788
rect -15788 3708 -9573 3772
rect -9509 3708 -9489 3772
rect -15788 3692 -9489 3708
rect -15788 3628 -9573 3692
rect -9509 3628 -9489 3692
rect -15788 3612 -9489 3628
rect -15788 3548 -9573 3612
rect -9509 3548 -9489 3612
rect -15788 3532 -9489 3548
rect -15788 3468 -9573 3532
rect -9509 3468 -9489 3532
rect -15788 3452 -9489 3468
rect -15788 3388 -9573 3452
rect -9509 3388 -9489 3452
rect -15788 3372 -9489 3388
rect -15788 3308 -9573 3372
rect -9509 3308 -9489 3372
rect -15788 3292 -9489 3308
rect -15788 3228 -9573 3292
rect -9509 3228 -9489 3292
rect -15788 3200 -9489 3228
rect -9469 9372 -3170 9400
rect -9469 9308 -3254 9372
rect -3190 9308 -3170 9372
rect -9469 9292 -3170 9308
rect -9469 9228 -3254 9292
rect -3190 9228 -3170 9292
rect -9469 9212 -3170 9228
rect -9469 9148 -3254 9212
rect -3190 9148 -3170 9212
rect -9469 9132 -3170 9148
rect -9469 9068 -3254 9132
rect -3190 9068 -3170 9132
rect -9469 9052 -3170 9068
rect -9469 8988 -3254 9052
rect -3190 8988 -3170 9052
rect -9469 8972 -3170 8988
rect -9469 8908 -3254 8972
rect -3190 8908 -3170 8972
rect -9469 8892 -3170 8908
rect -9469 8828 -3254 8892
rect -3190 8828 -3170 8892
rect -9469 8812 -3170 8828
rect -9469 8748 -3254 8812
rect -3190 8748 -3170 8812
rect -9469 8732 -3170 8748
rect -9469 8668 -3254 8732
rect -3190 8668 -3170 8732
rect -9469 8652 -3170 8668
rect -9469 8588 -3254 8652
rect -3190 8588 -3170 8652
rect -9469 8572 -3170 8588
rect -9469 8508 -3254 8572
rect -3190 8508 -3170 8572
rect -9469 8492 -3170 8508
rect -9469 8428 -3254 8492
rect -3190 8428 -3170 8492
rect -9469 8412 -3170 8428
rect -9469 8348 -3254 8412
rect -3190 8348 -3170 8412
rect -9469 8332 -3170 8348
rect -9469 8268 -3254 8332
rect -3190 8268 -3170 8332
rect -9469 8252 -3170 8268
rect -9469 8188 -3254 8252
rect -3190 8188 -3170 8252
rect -9469 8172 -3170 8188
rect -9469 8108 -3254 8172
rect -3190 8108 -3170 8172
rect -9469 8092 -3170 8108
rect -9469 8028 -3254 8092
rect -3190 8028 -3170 8092
rect -9469 8012 -3170 8028
rect -9469 7948 -3254 8012
rect -3190 7948 -3170 8012
rect -9469 7932 -3170 7948
rect -9469 7868 -3254 7932
rect -3190 7868 -3170 7932
rect -9469 7852 -3170 7868
rect -9469 7788 -3254 7852
rect -3190 7788 -3170 7852
rect -9469 7772 -3170 7788
rect -9469 7708 -3254 7772
rect -3190 7708 -3170 7772
rect -9469 7692 -3170 7708
rect -9469 7628 -3254 7692
rect -3190 7628 -3170 7692
rect -9469 7612 -3170 7628
rect -9469 7548 -3254 7612
rect -3190 7548 -3170 7612
rect -9469 7532 -3170 7548
rect -9469 7468 -3254 7532
rect -3190 7468 -3170 7532
rect -9469 7452 -3170 7468
rect -9469 7388 -3254 7452
rect -3190 7388 -3170 7452
rect -9469 7372 -3170 7388
rect -9469 7308 -3254 7372
rect -3190 7308 -3170 7372
rect -9469 7292 -3170 7308
rect -9469 7228 -3254 7292
rect -3190 7228 -3170 7292
rect -9469 7212 -3170 7228
rect -9469 7148 -3254 7212
rect -3190 7148 -3170 7212
rect -9469 7132 -3170 7148
rect -9469 7068 -3254 7132
rect -3190 7068 -3170 7132
rect -9469 7052 -3170 7068
rect -9469 6988 -3254 7052
rect -3190 6988 -3170 7052
rect -9469 6972 -3170 6988
rect -9469 6908 -3254 6972
rect -3190 6908 -3170 6972
rect -9469 6892 -3170 6908
rect -9469 6828 -3254 6892
rect -3190 6828 -3170 6892
rect -9469 6812 -3170 6828
rect -9469 6748 -3254 6812
rect -3190 6748 -3170 6812
rect -9469 6732 -3170 6748
rect -9469 6668 -3254 6732
rect -3190 6668 -3170 6732
rect -9469 6652 -3170 6668
rect -9469 6588 -3254 6652
rect -3190 6588 -3170 6652
rect -9469 6572 -3170 6588
rect -9469 6508 -3254 6572
rect -3190 6508 -3170 6572
rect -9469 6492 -3170 6508
rect -9469 6428 -3254 6492
rect -3190 6428 -3170 6492
rect -9469 6412 -3170 6428
rect -9469 6348 -3254 6412
rect -3190 6348 -3170 6412
rect -9469 6332 -3170 6348
rect -9469 6268 -3254 6332
rect -3190 6268 -3170 6332
rect -9469 6252 -3170 6268
rect -9469 6188 -3254 6252
rect -3190 6188 -3170 6252
rect -9469 6172 -3170 6188
rect -9469 6108 -3254 6172
rect -3190 6108 -3170 6172
rect -9469 6092 -3170 6108
rect -9469 6028 -3254 6092
rect -3190 6028 -3170 6092
rect -9469 6012 -3170 6028
rect -9469 5948 -3254 6012
rect -3190 5948 -3170 6012
rect -9469 5932 -3170 5948
rect -9469 5868 -3254 5932
rect -3190 5868 -3170 5932
rect -9469 5852 -3170 5868
rect -9469 5788 -3254 5852
rect -3190 5788 -3170 5852
rect -9469 5772 -3170 5788
rect -9469 5708 -3254 5772
rect -3190 5708 -3170 5772
rect -9469 5692 -3170 5708
rect -9469 5628 -3254 5692
rect -3190 5628 -3170 5692
rect -9469 5612 -3170 5628
rect -9469 5548 -3254 5612
rect -3190 5548 -3170 5612
rect -9469 5532 -3170 5548
rect -9469 5468 -3254 5532
rect -3190 5468 -3170 5532
rect -9469 5452 -3170 5468
rect -9469 5388 -3254 5452
rect -3190 5388 -3170 5452
rect -9469 5372 -3170 5388
rect -9469 5308 -3254 5372
rect -3190 5308 -3170 5372
rect -9469 5292 -3170 5308
rect -9469 5228 -3254 5292
rect -3190 5228 -3170 5292
rect -9469 5212 -3170 5228
rect -9469 5148 -3254 5212
rect -3190 5148 -3170 5212
rect -9469 5132 -3170 5148
rect -9469 5068 -3254 5132
rect -3190 5068 -3170 5132
rect -9469 5052 -3170 5068
rect -9469 4988 -3254 5052
rect -3190 4988 -3170 5052
rect -9469 4972 -3170 4988
rect -9469 4908 -3254 4972
rect -3190 4908 -3170 4972
rect -9469 4892 -3170 4908
rect -9469 4828 -3254 4892
rect -3190 4828 -3170 4892
rect -9469 4812 -3170 4828
rect -9469 4748 -3254 4812
rect -3190 4748 -3170 4812
rect -9469 4732 -3170 4748
rect -9469 4668 -3254 4732
rect -3190 4668 -3170 4732
rect -9469 4652 -3170 4668
rect -9469 4588 -3254 4652
rect -3190 4588 -3170 4652
rect -9469 4572 -3170 4588
rect -9469 4508 -3254 4572
rect -3190 4508 -3170 4572
rect -9469 4492 -3170 4508
rect -9469 4428 -3254 4492
rect -3190 4428 -3170 4492
rect -9469 4412 -3170 4428
rect -9469 4348 -3254 4412
rect -3190 4348 -3170 4412
rect -9469 4332 -3170 4348
rect -9469 4268 -3254 4332
rect -3190 4268 -3170 4332
rect -9469 4252 -3170 4268
rect -9469 4188 -3254 4252
rect -3190 4188 -3170 4252
rect -9469 4172 -3170 4188
rect -9469 4108 -3254 4172
rect -3190 4108 -3170 4172
rect -9469 4092 -3170 4108
rect -9469 4028 -3254 4092
rect -3190 4028 -3170 4092
rect -9469 4012 -3170 4028
rect -9469 3948 -3254 4012
rect -3190 3948 -3170 4012
rect -9469 3932 -3170 3948
rect -9469 3868 -3254 3932
rect -3190 3868 -3170 3932
rect -9469 3852 -3170 3868
rect -9469 3788 -3254 3852
rect -3190 3788 -3170 3852
rect -9469 3772 -3170 3788
rect -9469 3708 -3254 3772
rect -3190 3708 -3170 3772
rect -9469 3692 -3170 3708
rect -9469 3628 -3254 3692
rect -3190 3628 -3170 3692
rect -9469 3612 -3170 3628
rect -9469 3548 -3254 3612
rect -3190 3548 -3170 3612
rect -9469 3532 -3170 3548
rect -9469 3468 -3254 3532
rect -3190 3468 -3170 3532
rect -9469 3452 -3170 3468
rect -9469 3388 -3254 3452
rect -3190 3388 -3170 3452
rect -9469 3372 -3170 3388
rect -9469 3308 -3254 3372
rect -3190 3308 -3170 3372
rect -9469 3292 -3170 3308
rect -9469 3228 -3254 3292
rect -3190 3228 -3170 3292
rect -9469 3200 -3170 3228
rect -3150 9372 3149 9400
rect -3150 9308 3065 9372
rect 3129 9308 3149 9372
rect -3150 9292 3149 9308
rect -3150 9228 3065 9292
rect 3129 9228 3149 9292
rect -3150 9212 3149 9228
rect -3150 9148 3065 9212
rect 3129 9148 3149 9212
rect -3150 9132 3149 9148
rect -3150 9068 3065 9132
rect 3129 9068 3149 9132
rect -3150 9052 3149 9068
rect -3150 8988 3065 9052
rect 3129 8988 3149 9052
rect -3150 8972 3149 8988
rect -3150 8908 3065 8972
rect 3129 8908 3149 8972
rect -3150 8892 3149 8908
rect -3150 8828 3065 8892
rect 3129 8828 3149 8892
rect -3150 8812 3149 8828
rect -3150 8748 3065 8812
rect 3129 8748 3149 8812
rect -3150 8732 3149 8748
rect -3150 8668 3065 8732
rect 3129 8668 3149 8732
rect -3150 8652 3149 8668
rect -3150 8588 3065 8652
rect 3129 8588 3149 8652
rect -3150 8572 3149 8588
rect -3150 8508 3065 8572
rect 3129 8508 3149 8572
rect -3150 8492 3149 8508
rect -3150 8428 3065 8492
rect 3129 8428 3149 8492
rect -3150 8412 3149 8428
rect -3150 8348 3065 8412
rect 3129 8348 3149 8412
rect -3150 8332 3149 8348
rect -3150 8268 3065 8332
rect 3129 8268 3149 8332
rect -3150 8252 3149 8268
rect -3150 8188 3065 8252
rect 3129 8188 3149 8252
rect -3150 8172 3149 8188
rect -3150 8108 3065 8172
rect 3129 8108 3149 8172
rect -3150 8092 3149 8108
rect -3150 8028 3065 8092
rect 3129 8028 3149 8092
rect -3150 8012 3149 8028
rect -3150 7948 3065 8012
rect 3129 7948 3149 8012
rect -3150 7932 3149 7948
rect -3150 7868 3065 7932
rect 3129 7868 3149 7932
rect -3150 7852 3149 7868
rect -3150 7788 3065 7852
rect 3129 7788 3149 7852
rect -3150 7772 3149 7788
rect -3150 7708 3065 7772
rect 3129 7708 3149 7772
rect -3150 7692 3149 7708
rect -3150 7628 3065 7692
rect 3129 7628 3149 7692
rect -3150 7612 3149 7628
rect -3150 7548 3065 7612
rect 3129 7548 3149 7612
rect -3150 7532 3149 7548
rect -3150 7468 3065 7532
rect 3129 7468 3149 7532
rect -3150 7452 3149 7468
rect -3150 7388 3065 7452
rect 3129 7388 3149 7452
rect -3150 7372 3149 7388
rect -3150 7308 3065 7372
rect 3129 7308 3149 7372
rect -3150 7292 3149 7308
rect -3150 7228 3065 7292
rect 3129 7228 3149 7292
rect -3150 7212 3149 7228
rect -3150 7148 3065 7212
rect 3129 7148 3149 7212
rect -3150 7132 3149 7148
rect -3150 7068 3065 7132
rect 3129 7068 3149 7132
rect -3150 7052 3149 7068
rect -3150 6988 3065 7052
rect 3129 6988 3149 7052
rect -3150 6972 3149 6988
rect -3150 6908 3065 6972
rect 3129 6908 3149 6972
rect -3150 6892 3149 6908
rect -3150 6828 3065 6892
rect 3129 6828 3149 6892
rect -3150 6812 3149 6828
rect -3150 6748 3065 6812
rect 3129 6748 3149 6812
rect -3150 6732 3149 6748
rect -3150 6668 3065 6732
rect 3129 6668 3149 6732
rect -3150 6652 3149 6668
rect -3150 6588 3065 6652
rect 3129 6588 3149 6652
rect -3150 6572 3149 6588
rect -3150 6508 3065 6572
rect 3129 6508 3149 6572
rect -3150 6492 3149 6508
rect -3150 6428 3065 6492
rect 3129 6428 3149 6492
rect -3150 6412 3149 6428
rect -3150 6348 3065 6412
rect 3129 6348 3149 6412
rect -3150 6332 3149 6348
rect -3150 6268 3065 6332
rect 3129 6268 3149 6332
rect -3150 6252 3149 6268
rect -3150 6188 3065 6252
rect 3129 6188 3149 6252
rect -3150 6172 3149 6188
rect -3150 6108 3065 6172
rect 3129 6108 3149 6172
rect -3150 6092 3149 6108
rect -3150 6028 3065 6092
rect 3129 6028 3149 6092
rect -3150 6012 3149 6028
rect -3150 5948 3065 6012
rect 3129 5948 3149 6012
rect -3150 5932 3149 5948
rect -3150 5868 3065 5932
rect 3129 5868 3149 5932
rect -3150 5852 3149 5868
rect -3150 5788 3065 5852
rect 3129 5788 3149 5852
rect -3150 5772 3149 5788
rect -3150 5708 3065 5772
rect 3129 5708 3149 5772
rect -3150 5692 3149 5708
rect -3150 5628 3065 5692
rect 3129 5628 3149 5692
rect -3150 5612 3149 5628
rect -3150 5548 3065 5612
rect 3129 5548 3149 5612
rect -3150 5532 3149 5548
rect -3150 5468 3065 5532
rect 3129 5468 3149 5532
rect -3150 5452 3149 5468
rect -3150 5388 3065 5452
rect 3129 5388 3149 5452
rect -3150 5372 3149 5388
rect -3150 5308 3065 5372
rect 3129 5308 3149 5372
rect -3150 5292 3149 5308
rect -3150 5228 3065 5292
rect 3129 5228 3149 5292
rect -3150 5212 3149 5228
rect -3150 5148 3065 5212
rect 3129 5148 3149 5212
rect -3150 5132 3149 5148
rect -3150 5068 3065 5132
rect 3129 5068 3149 5132
rect -3150 5052 3149 5068
rect -3150 4988 3065 5052
rect 3129 4988 3149 5052
rect -3150 4972 3149 4988
rect -3150 4908 3065 4972
rect 3129 4908 3149 4972
rect -3150 4892 3149 4908
rect -3150 4828 3065 4892
rect 3129 4828 3149 4892
rect -3150 4812 3149 4828
rect -3150 4748 3065 4812
rect 3129 4748 3149 4812
rect -3150 4732 3149 4748
rect -3150 4668 3065 4732
rect 3129 4668 3149 4732
rect -3150 4652 3149 4668
rect -3150 4588 3065 4652
rect 3129 4588 3149 4652
rect -3150 4572 3149 4588
rect -3150 4508 3065 4572
rect 3129 4508 3149 4572
rect -3150 4492 3149 4508
rect -3150 4428 3065 4492
rect 3129 4428 3149 4492
rect -3150 4412 3149 4428
rect -3150 4348 3065 4412
rect 3129 4348 3149 4412
rect -3150 4332 3149 4348
rect -3150 4268 3065 4332
rect 3129 4268 3149 4332
rect -3150 4252 3149 4268
rect -3150 4188 3065 4252
rect 3129 4188 3149 4252
rect -3150 4172 3149 4188
rect -3150 4108 3065 4172
rect 3129 4108 3149 4172
rect -3150 4092 3149 4108
rect -3150 4028 3065 4092
rect 3129 4028 3149 4092
rect -3150 4012 3149 4028
rect -3150 3948 3065 4012
rect 3129 3948 3149 4012
rect -3150 3932 3149 3948
rect -3150 3868 3065 3932
rect 3129 3868 3149 3932
rect -3150 3852 3149 3868
rect -3150 3788 3065 3852
rect 3129 3788 3149 3852
rect -3150 3772 3149 3788
rect -3150 3708 3065 3772
rect 3129 3708 3149 3772
rect -3150 3692 3149 3708
rect -3150 3628 3065 3692
rect 3129 3628 3149 3692
rect -3150 3612 3149 3628
rect -3150 3548 3065 3612
rect 3129 3548 3149 3612
rect -3150 3532 3149 3548
rect -3150 3468 3065 3532
rect 3129 3468 3149 3532
rect -3150 3452 3149 3468
rect -3150 3388 3065 3452
rect 3129 3388 3149 3452
rect -3150 3372 3149 3388
rect -3150 3308 3065 3372
rect 3129 3308 3149 3372
rect -3150 3292 3149 3308
rect -3150 3228 3065 3292
rect 3129 3228 3149 3292
rect -3150 3200 3149 3228
rect 3169 9372 9468 9400
rect 3169 9308 9384 9372
rect 9448 9308 9468 9372
rect 3169 9292 9468 9308
rect 3169 9228 9384 9292
rect 9448 9228 9468 9292
rect 3169 9212 9468 9228
rect 3169 9148 9384 9212
rect 9448 9148 9468 9212
rect 3169 9132 9468 9148
rect 3169 9068 9384 9132
rect 9448 9068 9468 9132
rect 3169 9052 9468 9068
rect 3169 8988 9384 9052
rect 9448 8988 9468 9052
rect 3169 8972 9468 8988
rect 3169 8908 9384 8972
rect 9448 8908 9468 8972
rect 3169 8892 9468 8908
rect 3169 8828 9384 8892
rect 9448 8828 9468 8892
rect 3169 8812 9468 8828
rect 3169 8748 9384 8812
rect 9448 8748 9468 8812
rect 3169 8732 9468 8748
rect 3169 8668 9384 8732
rect 9448 8668 9468 8732
rect 3169 8652 9468 8668
rect 3169 8588 9384 8652
rect 9448 8588 9468 8652
rect 3169 8572 9468 8588
rect 3169 8508 9384 8572
rect 9448 8508 9468 8572
rect 3169 8492 9468 8508
rect 3169 8428 9384 8492
rect 9448 8428 9468 8492
rect 3169 8412 9468 8428
rect 3169 8348 9384 8412
rect 9448 8348 9468 8412
rect 3169 8332 9468 8348
rect 3169 8268 9384 8332
rect 9448 8268 9468 8332
rect 3169 8252 9468 8268
rect 3169 8188 9384 8252
rect 9448 8188 9468 8252
rect 3169 8172 9468 8188
rect 3169 8108 9384 8172
rect 9448 8108 9468 8172
rect 3169 8092 9468 8108
rect 3169 8028 9384 8092
rect 9448 8028 9468 8092
rect 3169 8012 9468 8028
rect 3169 7948 9384 8012
rect 9448 7948 9468 8012
rect 3169 7932 9468 7948
rect 3169 7868 9384 7932
rect 9448 7868 9468 7932
rect 3169 7852 9468 7868
rect 3169 7788 9384 7852
rect 9448 7788 9468 7852
rect 3169 7772 9468 7788
rect 3169 7708 9384 7772
rect 9448 7708 9468 7772
rect 3169 7692 9468 7708
rect 3169 7628 9384 7692
rect 9448 7628 9468 7692
rect 3169 7612 9468 7628
rect 3169 7548 9384 7612
rect 9448 7548 9468 7612
rect 3169 7532 9468 7548
rect 3169 7468 9384 7532
rect 9448 7468 9468 7532
rect 3169 7452 9468 7468
rect 3169 7388 9384 7452
rect 9448 7388 9468 7452
rect 3169 7372 9468 7388
rect 3169 7308 9384 7372
rect 9448 7308 9468 7372
rect 3169 7292 9468 7308
rect 3169 7228 9384 7292
rect 9448 7228 9468 7292
rect 3169 7212 9468 7228
rect 3169 7148 9384 7212
rect 9448 7148 9468 7212
rect 3169 7132 9468 7148
rect 3169 7068 9384 7132
rect 9448 7068 9468 7132
rect 3169 7052 9468 7068
rect 3169 6988 9384 7052
rect 9448 6988 9468 7052
rect 3169 6972 9468 6988
rect 3169 6908 9384 6972
rect 9448 6908 9468 6972
rect 3169 6892 9468 6908
rect 3169 6828 9384 6892
rect 9448 6828 9468 6892
rect 3169 6812 9468 6828
rect 3169 6748 9384 6812
rect 9448 6748 9468 6812
rect 3169 6732 9468 6748
rect 3169 6668 9384 6732
rect 9448 6668 9468 6732
rect 3169 6652 9468 6668
rect 3169 6588 9384 6652
rect 9448 6588 9468 6652
rect 3169 6572 9468 6588
rect 3169 6508 9384 6572
rect 9448 6508 9468 6572
rect 3169 6492 9468 6508
rect 3169 6428 9384 6492
rect 9448 6428 9468 6492
rect 3169 6412 9468 6428
rect 3169 6348 9384 6412
rect 9448 6348 9468 6412
rect 3169 6332 9468 6348
rect 3169 6268 9384 6332
rect 9448 6268 9468 6332
rect 3169 6252 9468 6268
rect 3169 6188 9384 6252
rect 9448 6188 9468 6252
rect 3169 6172 9468 6188
rect 3169 6108 9384 6172
rect 9448 6108 9468 6172
rect 3169 6092 9468 6108
rect 3169 6028 9384 6092
rect 9448 6028 9468 6092
rect 3169 6012 9468 6028
rect 3169 5948 9384 6012
rect 9448 5948 9468 6012
rect 3169 5932 9468 5948
rect 3169 5868 9384 5932
rect 9448 5868 9468 5932
rect 3169 5852 9468 5868
rect 3169 5788 9384 5852
rect 9448 5788 9468 5852
rect 3169 5772 9468 5788
rect 3169 5708 9384 5772
rect 9448 5708 9468 5772
rect 3169 5692 9468 5708
rect 3169 5628 9384 5692
rect 9448 5628 9468 5692
rect 3169 5612 9468 5628
rect 3169 5548 9384 5612
rect 9448 5548 9468 5612
rect 3169 5532 9468 5548
rect 3169 5468 9384 5532
rect 9448 5468 9468 5532
rect 3169 5452 9468 5468
rect 3169 5388 9384 5452
rect 9448 5388 9468 5452
rect 3169 5372 9468 5388
rect 3169 5308 9384 5372
rect 9448 5308 9468 5372
rect 3169 5292 9468 5308
rect 3169 5228 9384 5292
rect 9448 5228 9468 5292
rect 3169 5212 9468 5228
rect 3169 5148 9384 5212
rect 9448 5148 9468 5212
rect 3169 5132 9468 5148
rect 3169 5068 9384 5132
rect 9448 5068 9468 5132
rect 3169 5052 9468 5068
rect 3169 4988 9384 5052
rect 9448 4988 9468 5052
rect 3169 4972 9468 4988
rect 3169 4908 9384 4972
rect 9448 4908 9468 4972
rect 3169 4892 9468 4908
rect 3169 4828 9384 4892
rect 9448 4828 9468 4892
rect 3169 4812 9468 4828
rect 3169 4748 9384 4812
rect 9448 4748 9468 4812
rect 3169 4732 9468 4748
rect 3169 4668 9384 4732
rect 9448 4668 9468 4732
rect 3169 4652 9468 4668
rect 3169 4588 9384 4652
rect 9448 4588 9468 4652
rect 3169 4572 9468 4588
rect 3169 4508 9384 4572
rect 9448 4508 9468 4572
rect 3169 4492 9468 4508
rect 3169 4428 9384 4492
rect 9448 4428 9468 4492
rect 3169 4412 9468 4428
rect 3169 4348 9384 4412
rect 9448 4348 9468 4412
rect 3169 4332 9468 4348
rect 3169 4268 9384 4332
rect 9448 4268 9468 4332
rect 3169 4252 9468 4268
rect 3169 4188 9384 4252
rect 9448 4188 9468 4252
rect 3169 4172 9468 4188
rect 3169 4108 9384 4172
rect 9448 4108 9468 4172
rect 3169 4092 9468 4108
rect 3169 4028 9384 4092
rect 9448 4028 9468 4092
rect 3169 4012 9468 4028
rect 3169 3948 9384 4012
rect 9448 3948 9468 4012
rect 3169 3932 9468 3948
rect 3169 3868 9384 3932
rect 9448 3868 9468 3932
rect 3169 3852 9468 3868
rect 3169 3788 9384 3852
rect 9448 3788 9468 3852
rect 3169 3772 9468 3788
rect 3169 3708 9384 3772
rect 9448 3708 9468 3772
rect 3169 3692 9468 3708
rect 3169 3628 9384 3692
rect 9448 3628 9468 3692
rect 3169 3612 9468 3628
rect 3169 3548 9384 3612
rect 9448 3548 9468 3612
rect 3169 3532 9468 3548
rect 3169 3468 9384 3532
rect 9448 3468 9468 3532
rect 3169 3452 9468 3468
rect 3169 3388 9384 3452
rect 9448 3388 9468 3452
rect 3169 3372 9468 3388
rect 3169 3308 9384 3372
rect 9448 3308 9468 3372
rect 3169 3292 9468 3308
rect 3169 3228 9384 3292
rect 9448 3228 9468 3292
rect 3169 3200 9468 3228
rect 9488 9372 15787 9400
rect 9488 9308 15703 9372
rect 15767 9308 15787 9372
rect 9488 9292 15787 9308
rect 9488 9228 15703 9292
rect 15767 9228 15787 9292
rect 9488 9212 15787 9228
rect 9488 9148 15703 9212
rect 15767 9148 15787 9212
rect 9488 9132 15787 9148
rect 9488 9068 15703 9132
rect 15767 9068 15787 9132
rect 9488 9052 15787 9068
rect 9488 8988 15703 9052
rect 15767 8988 15787 9052
rect 9488 8972 15787 8988
rect 9488 8908 15703 8972
rect 15767 8908 15787 8972
rect 9488 8892 15787 8908
rect 9488 8828 15703 8892
rect 15767 8828 15787 8892
rect 9488 8812 15787 8828
rect 9488 8748 15703 8812
rect 15767 8748 15787 8812
rect 9488 8732 15787 8748
rect 9488 8668 15703 8732
rect 15767 8668 15787 8732
rect 9488 8652 15787 8668
rect 9488 8588 15703 8652
rect 15767 8588 15787 8652
rect 9488 8572 15787 8588
rect 9488 8508 15703 8572
rect 15767 8508 15787 8572
rect 9488 8492 15787 8508
rect 9488 8428 15703 8492
rect 15767 8428 15787 8492
rect 9488 8412 15787 8428
rect 9488 8348 15703 8412
rect 15767 8348 15787 8412
rect 9488 8332 15787 8348
rect 9488 8268 15703 8332
rect 15767 8268 15787 8332
rect 9488 8252 15787 8268
rect 9488 8188 15703 8252
rect 15767 8188 15787 8252
rect 9488 8172 15787 8188
rect 9488 8108 15703 8172
rect 15767 8108 15787 8172
rect 9488 8092 15787 8108
rect 9488 8028 15703 8092
rect 15767 8028 15787 8092
rect 9488 8012 15787 8028
rect 9488 7948 15703 8012
rect 15767 7948 15787 8012
rect 9488 7932 15787 7948
rect 9488 7868 15703 7932
rect 15767 7868 15787 7932
rect 9488 7852 15787 7868
rect 9488 7788 15703 7852
rect 15767 7788 15787 7852
rect 9488 7772 15787 7788
rect 9488 7708 15703 7772
rect 15767 7708 15787 7772
rect 9488 7692 15787 7708
rect 9488 7628 15703 7692
rect 15767 7628 15787 7692
rect 9488 7612 15787 7628
rect 9488 7548 15703 7612
rect 15767 7548 15787 7612
rect 9488 7532 15787 7548
rect 9488 7468 15703 7532
rect 15767 7468 15787 7532
rect 9488 7452 15787 7468
rect 9488 7388 15703 7452
rect 15767 7388 15787 7452
rect 9488 7372 15787 7388
rect 9488 7308 15703 7372
rect 15767 7308 15787 7372
rect 9488 7292 15787 7308
rect 9488 7228 15703 7292
rect 15767 7228 15787 7292
rect 9488 7212 15787 7228
rect 9488 7148 15703 7212
rect 15767 7148 15787 7212
rect 9488 7132 15787 7148
rect 9488 7068 15703 7132
rect 15767 7068 15787 7132
rect 9488 7052 15787 7068
rect 9488 6988 15703 7052
rect 15767 6988 15787 7052
rect 9488 6972 15787 6988
rect 9488 6908 15703 6972
rect 15767 6908 15787 6972
rect 9488 6892 15787 6908
rect 9488 6828 15703 6892
rect 15767 6828 15787 6892
rect 9488 6812 15787 6828
rect 9488 6748 15703 6812
rect 15767 6748 15787 6812
rect 9488 6732 15787 6748
rect 9488 6668 15703 6732
rect 15767 6668 15787 6732
rect 9488 6652 15787 6668
rect 9488 6588 15703 6652
rect 15767 6588 15787 6652
rect 9488 6572 15787 6588
rect 9488 6508 15703 6572
rect 15767 6508 15787 6572
rect 9488 6492 15787 6508
rect 9488 6428 15703 6492
rect 15767 6428 15787 6492
rect 9488 6412 15787 6428
rect 9488 6348 15703 6412
rect 15767 6348 15787 6412
rect 9488 6332 15787 6348
rect 9488 6268 15703 6332
rect 15767 6268 15787 6332
rect 9488 6252 15787 6268
rect 9488 6188 15703 6252
rect 15767 6188 15787 6252
rect 9488 6172 15787 6188
rect 9488 6108 15703 6172
rect 15767 6108 15787 6172
rect 9488 6092 15787 6108
rect 9488 6028 15703 6092
rect 15767 6028 15787 6092
rect 9488 6012 15787 6028
rect 9488 5948 15703 6012
rect 15767 5948 15787 6012
rect 9488 5932 15787 5948
rect 9488 5868 15703 5932
rect 15767 5868 15787 5932
rect 9488 5852 15787 5868
rect 9488 5788 15703 5852
rect 15767 5788 15787 5852
rect 9488 5772 15787 5788
rect 9488 5708 15703 5772
rect 15767 5708 15787 5772
rect 9488 5692 15787 5708
rect 9488 5628 15703 5692
rect 15767 5628 15787 5692
rect 9488 5612 15787 5628
rect 9488 5548 15703 5612
rect 15767 5548 15787 5612
rect 9488 5532 15787 5548
rect 9488 5468 15703 5532
rect 15767 5468 15787 5532
rect 9488 5452 15787 5468
rect 9488 5388 15703 5452
rect 15767 5388 15787 5452
rect 9488 5372 15787 5388
rect 9488 5308 15703 5372
rect 15767 5308 15787 5372
rect 9488 5292 15787 5308
rect 9488 5228 15703 5292
rect 15767 5228 15787 5292
rect 9488 5212 15787 5228
rect 9488 5148 15703 5212
rect 15767 5148 15787 5212
rect 9488 5132 15787 5148
rect 9488 5068 15703 5132
rect 15767 5068 15787 5132
rect 9488 5052 15787 5068
rect 9488 4988 15703 5052
rect 15767 4988 15787 5052
rect 9488 4972 15787 4988
rect 9488 4908 15703 4972
rect 15767 4908 15787 4972
rect 9488 4892 15787 4908
rect 9488 4828 15703 4892
rect 15767 4828 15787 4892
rect 9488 4812 15787 4828
rect 9488 4748 15703 4812
rect 15767 4748 15787 4812
rect 9488 4732 15787 4748
rect 9488 4668 15703 4732
rect 15767 4668 15787 4732
rect 9488 4652 15787 4668
rect 9488 4588 15703 4652
rect 15767 4588 15787 4652
rect 9488 4572 15787 4588
rect 9488 4508 15703 4572
rect 15767 4508 15787 4572
rect 9488 4492 15787 4508
rect 9488 4428 15703 4492
rect 15767 4428 15787 4492
rect 9488 4412 15787 4428
rect 9488 4348 15703 4412
rect 15767 4348 15787 4412
rect 9488 4332 15787 4348
rect 9488 4268 15703 4332
rect 15767 4268 15787 4332
rect 9488 4252 15787 4268
rect 9488 4188 15703 4252
rect 15767 4188 15787 4252
rect 9488 4172 15787 4188
rect 9488 4108 15703 4172
rect 15767 4108 15787 4172
rect 9488 4092 15787 4108
rect 9488 4028 15703 4092
rect 15767 4028 15787 4092
rect 9488 4012 15787 4028
rect 9488 3948 15703 4012
rect 15767 3948 15787 4012
rect 9488 3932 15787 3948
rect 9488 3868 15703 3932
rect 15767 3868 15787 3932
rect 9488 3852 15787 3868
rect 9488 3788 15703 3852
rect 15767 3788 15787 3852
rect 9488 3772 15787 3788
rect 9488 3708 15703 3772
rect 15767 3708 15787 3772
rect 9488 3692 15787 3708
rect 9488 3628 15703 3692
rect 15767 3628 15787 3692
rect 9488 3612 15787 3628
rect 9488 3548 15703 3612
rect 15767 3548 15787 3612
rect 9488 3532 15787 3548
rect 9488 3468 15703 3532
rect 15767 3468 15787 3532
rect 9488 3452 15787 3468
rect 9488 3388 15703 3452
rect 15767 3388 15787 3452
rect 9488 3372 15787 3388
rect 9488 3308 15703 3372
rect 15767 3308 15787 3372
rect 9488 3292 15787 3308
rect 9488 3228 15703 3292
rect 15767 3228 15787 3292
rect 9488 3200 15787 3228
rect 15807 9372 22106 9400
rect 15807 9308 22022 9372
rect 22086 9308 22106 9372
rect 15807 9292 22106 9308
rect 15807 9228 22022 9292
rect 22086 9228 22106 9292
rect 15807 9212 22106 9228
rect 15807 9148 22022 9212
rect 22086 9148 22106 9212
rect 15807 9132 22106 9148
rect 15807 9068 22022 9132
rect 22086 9068 22106 9132
rect 15807 9052 22106 9068
rect 15807 8988 22022 9052
rect 22086 8988 22106 9052
rect 15807 8972 22106 8988
rect 15807 8908 22022 8972
rect 22086 8908 22106 8972
rect 15807 8892 22106 8908
rect 15807 8828 22022 8892
rect 22086 8828 22106 8892
rect 15807 8812 22106 8828
rect 15807 8748 22022 8812
rect 22086 8748 22106 8812
rect 15807 8732 22106 8748
rect 15807 8668 22022 8732
rect 22086 8668 22106 8732
rect 15807 8652 22106 8668
rect 15807 8588 22022 8652
rect 22086 8588 22106 8652
rect 15807 8572 22106 8588
rect 15807 8508 22022 8572
rect 22086 8508 22106 8572
rect 15807 8492 22106 8508
rect 15807 8428 22022 8492
rect 22086 8428 22106 8492
rect 15807 8412 22106 8428
rect 15807 8348 22022 8412
rect 22086 8348 22106 8412
rect 15807 8332 22106 8348
rect 15807 8268 22022 8332
rect 22086 8268 22106 8332
rect 15807 8252 22106 8268
rect 15807 8188 22022 8252
rect 22086 8188 22106 8252
rect 15807 8172 22106 8188
rect 15807 8108 22022 8172
rect 22086 8108 22106 8172
rect 15807 8092 22106 8108
rect 15807 8028 22022 8092
rect 22086 8028 22106 8092
rect 15807 8012 22106 8028
rect 15807 7948 22022 8012
rect 22086 7948 22106 8012
rect 15807 7932 22106 7948
rect 15807 7868 22022 7932
rect 22086 7868 22106 7932
rect 15807 7852 22106 7868
rect 15807 7788 22022 7852
rect 22086 7788 22106 7852
rect 15807 7772 22106 7788
rect 15807 7708 22022 7772
rect 22086 7708 22106 7772
rect 15807 7692 22106 7708
rect 15807 7628 22022 7692
rect 22086 7628 22106 7692
rect 15807 7612 22106 7628
rect 15807 7548 22022 7612
rect 22086 7548 22106 7612
rect 15807 7532 22106 7548
rect 15807 7468 22022 7532
rect 22086 7468 22106 7532
rect 15807 7452 22106 7468
rect 15807 7388 22022 7452
rect 22086 7388 22106 7452
rect 15807 7372 22106 7388
rect 15807 7308 22022 7372
rect 22086 7308 22106 7372
rect 15807 7292 22106 7308
rect 15807 7228 22022 7292
rect 22086 7228 22106 7292
rect 15807 7212 22106 7228
rect 15807 7148 22022 7212
rect 22086 7148 22106 7212
rect 15807 7132 22106 7148
rect 15807 7068 22022 7132
rect 22086 7068 22106 7132
rect 15807 7052 22106 7068
rect 15807 6988 22022 7052
rect 22086 6988 22106 7052
rect 15807 6972 22106 6988
rect 15807 6908 22022 6972
rect 22086 6908 22106 6972
rect 15807 6892 22106 6908
rect 15807 6828 22022 6892
rect 22086 6828 22106 6892
rect 15807 6812 22106 6828
rect 15807 6748 22022 6812
rect 22086 6748 22106 6812
rect 15807 6732 22106 6748
rect 15807 6668 22022 6732
rect 22086 6668 22106 6732
rect 15807 6652 22106 6668
rect 15807 6588 22022 6652
rect 22086 6588 22106 6652
rect 15807 6572 22106 6588
rect 15807 6508 22022 6572
rect 22086 6508 22106 6572
rect 15807 6492 22106 6508
rect 15807 6428 22022 6492
rect 22086 6428 22106 6492
rect 15807 6412 22106 6428
rect 15807 6348 22022 6412
rect 22086 6348 22106 6412
rect 15807 6332 22106 6348
rect 15807 6268 22022 6332
rect 22086 6268 22106 6332
rect 15807 6252 22106 6268
rect 15807 6188 22022 6252
rect 22086 6188 22106 6252
rect 15807 6172 22106 6188
rect 15807 6108 22022 6172
rect 22086 6108 22106 6172
rect 15807 6092 22106 6108
rect 15807 6028 22022 6092
rect 22086 6028 22106 6092
rect 15807 6012 22106 6028
rect 15807 5948 22022 6012
rect 22086 5948 22106 6012
rect 15807 5932 22106 5948
rect 15807 5868 22022 5932
rect 22086 5868 22106 5932
rect 15807 5852 22106 5868
rect 15807 5788 22022 5852
rect 22086 5788 22106 5852
rect 15807 5772 22106 5788
rect 15807 5708 22022 5772
rect 22086 5708 22106 5772
rect 15807 5692 22106 5708
rect 15807 5628 22022 5692
rect 22086 5628 22106 5692
rect 15807 5612 22106 5628
rect 15807 5548 22022 5612
rect 22086 5548 22106 5612
rect 15807 5532 22106 5548
rect 15807 5468 22022 5532
rect 22086 5468 22106 5532
rect 15807 5452 22106 5468
rect 15807 5388 22022 5452
rect 22086 5388 22106 5452
rect 15807 5372 22106 5388
rect 15807 5308 22022 5372
rect 22086 5308 22106 5372
rect 15807 5292 22106 5308
rect 15807 5228 22022 5292
rect 22086 5228 22106 5292
rect 15807 5212 22106 5228
rect 15807 5148 22022 5212
rect 22086 5148 22106 5212
rect 15807 5132 22106 5148
rect 15807 5068 22022 5132
rect 22086 5068 22106 5132
rect 15807 5052 22106 5068
rect 15807 4988 22022 5052
rect 22086 4988 22106 5052
rect 15807 4972 22106 4988
rect 15807 4908 22022 4972
rect 22086 4908 22106 4972
rect 15807 4892 22106 4908
rect 15807 4828 22022 4892
rect 22086 4828 22106 4892
rect 15807 4812 22106 4828
rect 15807 4748 22022 4812
rect 22086 4748 22106 4812
rect 15807 4732 22106 4748
rect 15807 4668 22022 4732
rect 22086 4668 22106 4732
rect 15807 4652 22106 4668
rect 15807 4588 22022 4652
rect 22086 4588 22106 4652
rect 15807 4572 22106 4588
rect 15807 4508 22022 4572
rect 22086 4508 22106 4572
rect 15807 4492 22106 4508
rect 15807 4428 22022 4492
rect 22086 4428 22106 4492
rect 15807 4412 22106 4428
rect 15807 4348 22022 4412
rect 22086 4348 22106 4412
rect 15807 4332 22106 4348
rect 15807 4268 22022 4332
rect 22086 4268 22106 4332
rect 15807 4252 22106 4268
rect 15807 4188 22022 4252
rect 22086 4188 22106 4252
rect 15807 4172 22106 4188
rect 15807 4108 22022 4172
rect 22086 4108 22106 4172
rect 15807 4092 22106 4108
rect 15807 4028 22022 4092
rect 22086 4028 22106 4092
rect 15807 4012 22106 4028
rect 15807 3948 22022 4012
rect 22086 3948 22106 4012
rect 15807 3932 22106 3948
rect 15807 3868 22022 3932
rect 22086 3868 22106 3932
rect 15807 3852 22106 3868
rect 15807 3788 22022 3852
rect 22086 3788 22106 3852
rect 15807 3772 22106 3788
rect 15807 3708 22022 3772
rect 22086 3708 22106 3772
rect 15807 3692 22106 3708
rect 15807 3628 22022 3692
rect 22086 3628 22106 3692
rect 15807 3612 22106 3628
rect 15807 3548 22022 3612
rect 22086 3548 22106 3612
rect 15807 3532 22106 3548
rect 15807 3468 22022 3532
rect 22086 3468 22106 3532
rect 15807 3452 22106 3468
rect 15807 3388 22022 3452
rect 22086 3388 22106 3452
rect 15807 3372 22106 3388
rect 15807 3308 22022 3372
rect 22086 3308 22106 3372
rect 15807 3292 22106 3308
rect 15807 3228 22022 3292
rect 22086 3228 22106 3292
rect 15807 3200 22106 3228
rect 22126 9372 28425 9400
rect 22126 9308 28341 9372
rect 28405 9308 28425 9372
rect 22126 9292 28425 9308
rect 22126 9228 28341 9292
rect 28405 9228 28425 9292
rect 22126 9212 28425 9228
rect 22126 9148 28341 9212
rect 28405 9148 28425 9212
rect 22126 9132 28425 9148
rect 22126 9068 28341 9132
rect 28405 9068 28425 9132
rect 22126 9052 28425 9068
rect 22126 8988 28341 9052
rect 28405 8988 28425 9052
rect 22126 8972 28425 8988
rect 22126 8908 28341 8972
rect 28405 8908 28425 8972
rect 22126 8892 28425 8908
rect 22126 8828 28341 8892
rect 28405 8828 28425 8892
rect 22126 8812 28425 8828
rect 22126 8748 28341 8812
rect 28405 8748 28425 8812
rect 22126 8732 28425 8748
rect 22126 8668 28341 8732
rect 28405 8668 28425 8732
rect 22126 8652 28425 8668
rect 22126 8588 28341 8652
rect 28405 8588 28425 8652
rect 22126 8572 28425 8588
rect 22126 8508 28341 8572
rect 28405 8508 28425 8572
rect 22126 8492 28425 8508
rect 22126 8428 28341 8492
rect 28405 8428 28425 8492
rect 22126 8412 28425 8428
rect 22126 8348 28341 8412
rect 28405 8348 28425 8412
rect 22126 8332 28425 8348
rect 22126 8268 28341 8332
rect 28405 8268 28425 8332
rect 22126 8252 28425 8268
rect 22126 8188 28341 8252
rect 28405 8188 28425 8252
rect 22126 8172 28425 8188
rect 22126 8108 28341 8172
rect 28405 8108 28425 8172
rect 22126 8092 28425 8108
rect 22126 8028 28341 8092
rect 28405 8028 28425 8092
rect 22126 8012 28425 8028
rect 22126 7948 28341 8012
rect 28405 7948 28425 8012
rect 22126 7932 28425 7948
rect 22126 7868 28341 7932
rect 28405 7868 28425 7932
rect 22126 7852 28425 7868
rect 22126 7788 28341 7852
rect 28405 7788 28425 7852
rect 22126 7772 28425 7788
rect 22126 7708 28341 7772
rect 28405 7708 28425 7772
rect 22126 7692 28425 7708
rect 22126 7628 28341 7692
rect 28405 7628 28425 7692
rect 22126 7612 28425 7628
rect 22126 7548 28341 7612
rect 28405 7548 28425 7612
rect 22126 7532 28425 7548
rect 22126 7468 28341 7532
rect 28405 7468 28425 7532
rect 22126 7452 28425 7468
rect 22126 7388 28341 7452
rect 28405 7388 28425 7452
rect 22126 7372 28425 7388
rect 22126 7308 28341 7372
rect 28405 7308 28425 7372
rect 22126 7292 28425 7308
rect 22126 7228 28341 7292
rect 28405 7228 28425 7292
rect 22126 7212 28425 7228
rect 22126 7148 28341 7212
rect 28405 7148 28425 7212
rect 22126 7132 28425 7148
rect 22126 7068 28341 7132
rect 28405 7068 28425 7132
rect 22126 7052 28425 7068
rect 22126 6988 28341 7052
rect 28405 6988 28425 7052
rect 22126 6972 28425 6988
rect 22126 6908 28341 6972
rect 28405 6908 28425 6972
rect 22126 6892 28425 6908
rect 22126 6828 28341 6892
rect 28405 6828 28425 6892
rect 22126 6812 28425 6828
rect 22126 6748 28341 6812
rect 28405 6748 28425 6812
rect 22126 6732 28425 6748
rect 22126 6668 28341 6732
rect 28405 6668 28425 6732
rect 22126 6652 28425 6668
rect 22126 6588 28341 6652
rect 28405 6588 28425 6652
rect 22126 6572 28425 6588
rect 22126 6508 28341 6572
rect 28405 6508 28425 6572
rect 22126 6492 28425 6508
rect 22126 6428 28341 6492
rect 28405 6428 28425 6492
rect 22126 6412 28425 6428
rect 22126 6348 28341 6412
rect 28405 6348 28425 6412
rect 22126 6332 28425 6348
rect 22126 6268 28341 6332
rect 28405 6268 28425 6332
rect 22126 6252 28425 6268
rect 22126 6188 28341 6252
rect 28405 6188 28425 6252
rect 22126 6172 28425 6188
rect 22126 6108 28341 6172
rect 28405 6108 28425 6172
rect 22126 6092 28425 6108
rect 22126 6028 28341 6092
rect 28405 6028 28425 6092
rect 22126 6012 28425 6028
rect 22126 5948 28341 6012
rect 28405 5948 28425 6012
rect 22126 5932 28425 5948
rect 22126 5868 28341 5932
rect 28405 5868 28425 5932
rect 22126 5852 28425 5868
rect 22126 5788 28341 5852
rect 28405 5788 28425 5852
rect 22126 5772 28425 5788
rect 22126 5708 28341 5772
rect 28405 5708 28425 5772
rect 22126 5692 28425 5708
rect 22126 5628 28341 5692
rect 28405 5628 28425 5692
rect 22126 5612 28425 5628
rect 22126 5548 28341 5612
rect 28405 5548 28425 5612
rect 22126 5532 28425 5548
rect 22126 5468 28341 5532
rect 28405 5468 28425 5532
rect 22126 5452 28425 5468
rect 22126 5388 28341 5452
rect 28405 5388 28425 5452
rect 22126 5372 28425 5388
rect 22126 5308 28341 5372
rect 28405 5308 28425 5372
rect 22126 5292 28425 5308
rect 22126 5228 28341 5292
rect 28405 5228 28425 5292
rect 22126 5212 28425 5228
rect 22126 5148 28341 5212
rect 28405 5148 28425 5212
rect 22126 5132 28425 5148
rect 22126 5068 28341 5132
rect 28405 5068 28425 5132
rect 22126 5052 28425 5068
rect 22126 4988 28341 5052
rect 28405 4988 28425 5052
rect 22126 4972 28425 4988
rect 22126 4908 28341 4972
rect 28405 4908 28425 4972
rect 22126 4892 28425 4908
rect 22126 4828 28341 4892
rect 28405 4828 28425 4892
rect 22126 4812 28425 4828
rect 22126 4748 28341 4812
rect 28405 4748 28425 4812
rect 22126 4732 28425 4748
rect 22126 4668 28341 4732
rect 28405 4668 28425 4732
rect 22126 4652 28425 4668
rect 22126 4588 28341 4652
rect 28405 4588 28425 4652
rect 22126 4572 28425 4588
rect 22126 4508 28341 4572
rect 28405 4508 28425 4572
rect 22126 4492 28425 4508
rect 22126 4428 28341 4492
rect 28405 4428 28425 4492
rect 22126 4412 28425 4428
rect 22126 4348 28341 4412
rect 28405 4348 28425 4412
rect 22126 4332 28425 4348
rect 22126 4268 28341 4332
rect 28405 4268 28425 4332
rect 22126 4252 28425 4268
rect 22126 4188 28341 4252
rect 28405 4188 28425 4252
rect 22126 4172 28425 4188
rect 22126 4108 28341 4172
rect 28405 4108 28425 4172
rect 22126 4092 28425 4108
rect 22126 4028 28341 4092
rect 28405 4028 28425 4092
rect 22126 4012 28425 4028
rect 22126 3948 28341 4012
rect 28405 3948 28425 4012
rect 22126 3932 28425 3948
rect 22126 3868 28341 3932
rect 28405 3868 28425 3932
rect 22126 3852 28425 3868
rect 22126 3788 28341 3852
rect 28405 3788 28425 3852
rect 22126 3772 28425 3788
rect 22126 3708 28341 3772
rect 28405 3708 28425 3772
rect 22126 3692 28425 3708
rect 22126 3628 28341 3692
rect 28405 3628 28425 3692
rect 22126 3612 28425 3628
rect 22126 3548 28341 3612
rect 28405 3548 28425 3612
rect 22126 3532 28425 3548
rect 22126 3468 28341 3532
rect 28405 3468 28425 3532
rect 22126 3452 28425 3468
rect 22126 3388 28341 3452
rect 28405 3388 28425 3452
rect 22126 3372 28425 3388
rect 22126 3308 28341 3372
rect 28405 3308 28425 3372
rect 22126 3292 28425 3308
rect 22126 3228 28341 3292
rect 28405 3228 28425 3292
rect 22126 3200 28425 3228
rect 28445 9372 34744 9400
rect 28445 9308 34660 9372
rect 34724 9308 34744 9372
rect 28445 9292 34744 9308
rect 28445 9228 34660 9292
rect 34724 9228 34744 9292
rect 28445 9212 34744 9228
rect 28445 9148 34660 9212
rect 34724 9148 34744 9212
rect 28445 9132 34744 9148
rect 28445 9068 34660 9132
rect 34724 9068 34744 9132
rect 28445 9052 34744 9068
rect 28445 8988 34660 9052
rect 34724 8988 34744 9052
rect 28445 8972 34744 8988
rect 28445 8908 34660 8972
rect 34724 8908 34744 8972
rect 28445 8892 34744 8908
rect 28445 8828 34660 8892
rect 34724 8828 34744 8892
rect 28445 8812 34744 8828
rect 28445 8748 34660 8812
rect 34724 8748 34744 8812
rect 28445 8732 34744 8748
rect 28445 8668 34660 8732
rect 34724 8668 34744 8732
rect 28445 8652 34744 8668
rect 28445 8588 34660 8652
rect 34724 8588 34744 8652
rect 28445 8572 34744 8588
rect 28445 8508 34660 8572
rect 34724 8508 34744 8572
rect 28445 8492 34744 8508
rect 28445 8428 34660 8492
rect 34724 8428 34744 8492
rect 28445 8412 34744 8428
rect 28445 8348 34660 8412
rect 34724 8348 34744 8412
rect 28445 8332 34744 8348
rect 28445 8268 34660 8332
rect 34724 8268 34744 8332
rect 28445 8252 34744 8268
rect 28445 8188 34660 8252
rect 34724 8188 34744 8252
rect 28445 8172 34744 8188
rect 28445 8108 34660 8172
rect 34724 8108 34744 8172
rect 28445 8092 34744 8108
rect 28445 8028 34660 8092
rect 34724 8028 34744 8092
rect 28445 8012 34744 8028
rect 28445 7948 34660 8012
rect 34724 7948 34744 8012
rect 28445 7932 34744 7948
rect 28445 7868 34660 7932
rect 34724 7868 34744 7932
rect 28445 7852 34744 7868
rect 28445 7788 34660 7852
rect 34724 7788 34744 7852
rect 28445 7772 34744 7788
rect 28445 7708 34660 7772
rect 34724 7708 34744 7772
rect 28445 7692 34744 7708
rect 28445 7628 34660 7692
rect 34724 7628 34744 7692
rect 28445 7612 34744 7628
rect 28445 7548 34660 7612
rect 34724 7548 34744 7612
rect 28445 7532 34744 7548
rect 28445 7468 34660 7532
rect 34724 7468 34744 7532
rect 28445 7452 34744 7468
rect 28445 7388 34660 7452
rect 34724 7388 34744 7452
rect 28445 7372 34744 7388
rect 28445 7308 34660 7372
rect 34724 7308 34744 7372
rect 28445 7292 34744 7308
rect 28445 7228 34660 7292
rect 34724 7228 34744 7292
rect 28445 7212 34744 7228
rect 28445 7148 34660 7212
rect 34724 7148 34744 7212
rect 28445 7132 34744 7148
rect 28445 7068 34660 7132
rect 34724 7068 34744 7132
rect 28445 7052 34744 7068
rect 28445 6988 34660 7052
rect 34724 6988 34744 7052
rect 28445 6972 34744 6988
rect 28445 6908 34660 6972
rect 34724 6908 34744 6972
rect 28445 6892 34744 6908
rect 28445 6828 34660 6892
rect 34724 6828 34744 6892
rect 28445 6812 34744 6828
rect 28445 6748 34660 6812
rect 34724 6748 34744 6812
rect 28445 6732 34744 6748
rect 28445 6668 34660 6732
rect 34724 6668 34744 6732
rect 28445 6652 34744 6668
rect 28445 6588 34660 6652
rect 34724 6588 34744 6652
rect 28445 6572 34744 6588
rect 28445 6508 34660 6572
rect 34724 6508 34744 6572
rect 28445 6492 34744 6508
rect 28445 6428 34660 6492
rect 34724 6428 34744 6492
rect 28445 6412 34744 6428
rect 28445 6348 34660 6412
rect 34724 6348 34744 6412
rect 28445 6332 34744 6348
rect 28445 6268 34660 6332
rect 34724 6268 34744 6332
rect 28445 6252 34744 6268
rect 28445 6188 34660 6252
rect 34724 6188 34744 6252
rect 28445 6172 34744 6188
rect 28445 6108 34660 6172
rect 34724 6108 34744 6172
rect 28445 6092 34744 6108
rect 28445 6028 34660 6092
rect 34724 6028 34744 6092
rect 28445 6012 34744 6028
rect 28445 5948 34660 6012
rect 34724 5948 34744 6012
rect 28445 5932 34744 5948
rect 28445 5868 34660 5932
rect 34724 5868 34744 5932
rect 28445 5852 34744 5868
rect 28445 5788 34660 5852
rect 34724 5788 34744 5852
rect 28445 5772 34744 5788
rect 28445 5708 34660 5772
rect 34724 5708 34744 5772
rect 28445 5692 34744 5708
rect 28445 5628 34660 5692
rect 34724 5628 34744 5692
rect 28445 5612 34744 5628
rect 28445 5548 34660 5612
rect 34724 5548 34744 5612
rect 28445 5532 34744 5548
rect 28445 5468 34660 5532
rect 34724 5468 34744 5532
rect 28445 5452 34744 5468
rect 28445 5388 34660 5452
rect 34724 5388 34744 5452
rect 28445 5372 34744 5388
rect 28445 5308 34660 5372
rect 34724 5308 34744 5372
rect 28445 5292 34744 5308
rect 28445 5228 34660 5292
rect 34724 5228 34744 5292
rect 28445 5212 34744 5228
rect 28445 5148 34660 5212
rect 34724 5148 34744 5212
rect 28445 5132 34744 5148
rect 28445 5068 34660 5132
rect 34724 5068 34744 5132
rect 28445 5052 34744 5068
rect 28445 4988 34660 5052
rect 34724 4988 34744 5052
rect 28445 4972 34744 4988
rect 28445 4908 34660 4972
rect 34724 4908 34744 4972
rect 28445 4892 34744 4908
rect 28445 4828 34660 4892
rect 34724 4828 34744 4892
rect 28445 4812 34744 4828
rect 28445 4748 34660 4812
rect 34724 4748 34744 4812
rect 28445 4732 34744 4748
rect 28445 4668 34660 4732
rect 34724 4668 34744 4732
rect 28445 4652 34744 4668
rect 28445 4588 34660 4652
rect 34724 4588 34744 4652
rect 28445 4572 34744 4588
rect 28445 4508 34660 4572
rect 34724 4508 34744 4572
rect 28445 4492 34744 4508
rect 28445 4428 34660 4492
rect 34724 4428 34744 4492
rect 28445 4412 34744 4428
rect 28445 4348 34660 4412
rect 34724 4348 34744 4412
rect 28445 4332 34744 4348
rect 28445 4268 34660 4332
rect 34724 4268 34744 4332
rect 28445 4252 34744 4268
rect 28445 4188 34660 4252
rect 34724 4188 34744 4252
rect 28445 4172 34744 4188
rect 28445 4108 34660 4172
rect 34724 4108 34744 4172
rect 28445 4092 34744 4108
rect 28445 4028 34660 4092
rect 34724 4028 34744 4092
rect 28445 4012 34744 4028
rect 28445 3948 34660 4012
rect 34724 3948 34744 4012
rect 28445 3932 34744 3948
rect 28445 3868 34660 3932
rect 34724 3868 34744 3932
rect 28445 3852 34744 3868
rect 28445 3788 34660 3852
rect 34724 3788 34744 3852
rect 28445 3772 34744 3788
rect 28445 3708 34660 3772
rect 34724 3708 34744 3772
rect 28445 3692 34744 3708
rect 28445 3628 34660 3692
rect 34724 3628 34744 3692
rect 28445 3612 34744 3628
rect 28445 3548 34660 3612
rect 34724 3548 34744 3612
rect 28445 3532 34744 3548
rect 28445 3468 34660 3532
rect 34724 3468 34744 3532
rect 28445 3452 34744 3468
rect 28445 3388 34660 3452
rect 34724 3388 34744 3452
rect 28445 3372 34744 3388
rect 28445 3308 34660 3372
rect 34724 3308 34744 3372
rect 28445 3292 34744 3308
rect 28445 3228 34660 3292
rect 34724 3228 34744 3292
rect 28445 3200 34744 3228
rect 34764 9372 41063 9400
rect 34764 9308 40979 9372
rect 41043 9308 41063 9372
rect 34764 9292 41063 9308
rect 34764 9228 40979 9292
rect 41043 9228 41063 9292
rect 34764 9212 41063 9228
rect 34764 9148 40979 9212
rect 41043 9148 41063 9212
rect 34764 9132 41063 9148
rect 34764 9068 40979 9132
rect 41043 9068 41063 9132
rect 34764 9052 41063 9068
rect 34764 8988 40979 9052
rect 41043 8988 41063 9052
rect 34764 8972 41063 8988
rect 34764 8908 40979 8972
rect 41043 8908 41063 8972
rect 34764 8892 41063 8908
rect 34764 8828 40979 8892
rect 41043 8828 41063 8892
rect 34764 8812 41063 8828
rect 34764 8748 40979 8812
rect 41043 8748 41063 8812
rect 34764 8732 41063 8748
rect 34764 8668 40979 8732
rect 41043 8668 41063 8732
rect 34764 8652 41063 8668
rect 34764 8588 40979 8652
rect 41043 8588 41063 8652
rect 34764 8572 41063 8588
rect 34764 8508 40979 8572
rect 41043 8508 41063 8572
rect 34764 8492 41063 8508
rect 34764 8428 40979 8492
rect 41043 8428 41063 8492
rect 34764 8412 41063 8428
rect 34764 8348 40979 8412
rect 41043 8348 41063 8412
rect 34764 8332 41063 8348
rect 34764 8268 40979 8332
rect 41043 8268 41063 8332
rect 34764 8252 41063 8268
rect 34764 8188 40979 8252
rect 41043 8188 41063 8252
rect 34764 8172 41063 8188
rect 34764 8108 40979 8172
rect 41043 8108 41063 8172
rect 34764 8092 41063 8108
rect 34764 8028 40979 8092
rect 41043 8028 41063 8092
rect 34764 8012 41063 8028
rect 34764 7948 40979 8012
rect 41043 7948 41063 8012
rect 34764 7932 41063 7948
rect 34764 7868 40979 7932
rect 41043 7868 41063 7932
rect 34764 7852 41063 7868
rect 34764 7788 40979 7852
rect 41043 7788 41063 7852
rect 34764 7772 41063 7788
rect 34764 7708 40979 7772
rect 41043 7708 41063 7772
rect 34764 7692 41063 7708
rect 34764 7628 40979 7692
rect 41043 7628 41063 7692
rect 34764 7612 41063 7628
rect 34764 7548 40979 7612
rect 41043 7548 41063 7612
rect 34764 7532 41063 7548
rect 34764 7468 40979 7532
rect 41043 7468 41063 7532
rect 34764 7452 41063 7468
rect 34764 7388 40979 7452
rect 41043 7388 41063 7452
rect 34764 7372 41063 7388
rect 34764 7308 40979 7372
rect 41043 7308 41063 7372
rect 34764 7292 41063 7308
rect 34764 7228 40979 7292
rect 41043 7228 41063 7292
rect 34764 7212 41063 7228
rect 34764 7148 40979 7212
rect 41043 7148 41063 7212
rect 34764 7132 41063 7148
rect 34764 7068 40979 7132
rect 41043 7068 41063 7132
rect 34764 7052 41063 7068
rect 34764 6988 40979 7052
rect 41043 6988 41063 7052
rect 34764 6972 41063 6988
rect 34764 6908 40979 6972
rect 41043 6908 41063 6972
rect 34764 6892 41063 6908
rect 34764 6828 40979 6892
rect 41043 6828 41063 6892
rect 34764 6812 41063 6828
rect 34764 6748 40979 6812
rect 41043 6748 41063 6812
rect 34764 6732 41063 6748
rect 34764 6668 40979 6732
rect 41043 6668 41063 6732
rect 34764 6652 41063 6668
rect 34764 6588 40979 6652
rect 41043 6588 41063 6652
rect 34764 6572 41063 6588
rect 34764 6508 40979 6572
rect 41043 6508 41063 6572
rect 34764 6492 41063 6508
rect 34764 6428 40979 6492
rect 41043 6428 41063 6492
rect 34764 6412 41063 6428
rect 34764 6348 40979 6412
rect 41043 6348 41063 6412
rect 34764 6332 41063 6348
rect 34764 6268 40979 6332
rect 41043 6268 41063 6332
rect 34764 6252 41063 6268
rect 34764 6188 40979 6252
rect 41043 6188 41063 6252
rect 34764 6172 41063 6188
rect 34764 6108 40979 6172
rect 41043 6108 41063 6172
rect 34764 6092 41063 6108
rect 34764 6028 40979 6092
rect 41043 6028 41063 6092
rect 34764 6012 41063 6028
rect 34764 5948 40979 6012
rect 41043 5948 41063 6012
rect 34764 5932 41063 5948
rect 34764 5868 40979 5932
rect 41043 5868 41063 5932
rect 34764 5852 41063 5868
rect 34764 5788 40979 5852
rect 41043 5788 41063 5852
rect 34764 5772 41063 5788
rect 34764 5708 40979 5772
rect 41043 5708 41063 5772
rect 34764 5692 41063 5708
rect 34764 5628 40979 5692
rect 41043 5628 41063 5692
rect 34764 5612 41063 5628
rect 34764 5548 40979 5612
rect 41043 5548 41063 5612
rect 34764 5532 41063 5548
rect 34764 5468 40979 5532
rect 41043 5468 41063 5532
rect 34764 5452 41063 5468
rect 34764 5388 40979 5452
rect 41043 5388 41063 5452
rect 34764 5372 41063 5388
rect 34764 5308 40979 5372
rect 41043 5308 41063 5372
rect 34764 5292 41063 5308
rect 34764 5228 40979 5292
rect 41043 5228 41063 5292
rect 34764 5212 41063 5228
rect 34764 5148 40979 5212
rect 41043 5148 41063 5212
rect 34764 5132 41063 5148
rect 34764 5068 40979 5132
rect 41043 5068 41063 5132
rect 34764 5052 41063 5068
rect 34764 4988 40979 5052
rect 41043 4988 41063 5052
rect 34764 4972 41063 4988
rect 34764 4908 40979 4972
rect 41043 4908 41063 4972
rect 34764 4892 41063 4908
rect 34764 4828 40979 4892
rect 41043 4828 41063 4892
rect 34764 4812 41063 4828
rect 34764 4748 40979 4812
rect 41043 4748 41063 4812
rect 34764 4732 41063 4748
rect 34764 4668 40979 4732
rect 41043 4668 41063 4732
rect 34764 4652 41063 4668
rect 34764 4588 40979 4652
rect 41043 4588 41063 4652
rect 34764 4572 41063 4588
rect 34764 4508 40979 4572
rect 41043 4508 41063 4572
rect 34764 4492 41063 4508
rect 34764 4428 40979 4492
rect 41043 4428 41063 4492
rect 34764 4412 41063 4428
rect 34764 4348 40979 4412
rect 41043 4348 41063 4412
rect 34764 4332 41063 4348
rect 34764 4268 40979 4332
rect 41043 4268 41063 4332
rect 34764 4252 41063 4268
rect 34764 4188 40979 4252
rect 41043 4188 41063 4252
rect 34764 4172 41063 4188
rect 34764 4108 40979 4172
rect 41043 4108 41063 4172
rect 34764 4092 41063 4108
rect 34764 4028 40979 4092
rect 41043 4028 41063 4092
rect 34764 4012 41063 4028
rect 34764 3948 40979 4012
rect 41043 3948 41063 4012
rect 34764 3932 41063 3948
rect 34764 3868 40979 3932
rect 41043 3868 41063 3932
rect 34764 3852 41063 3868
rect 34764 3788 40979 3852
rect 41043 3788 41063 3852
rect 34764 3772 41063 3788
rect 34764 3708 40979 3772
rect 41043 3708 41063 3772
rect 34764 3692 41063 3708
rect 34764 3628 40979 3692
rect 41043 3628 41063 3692
rect 34764 3612 41063 3628
rect 34764 3548 40979 3612
rect 41043 3548 41063 3612
rect 34764 3532 41063 3548
rect 34764 3468 40979 3532
rect 41043 3468 41063 3532
rect 34764 3452 41063 3468
rect 34764 3388 40979 3452
rect 41043 3388 41063 3452
rect 34764 3372 41063 3388
rect 34764 3308 40979 3372
rect 41043 3308 41063 3372
rect 34764 3292 41063 3308
rect 34764 3228 40979 3292
rect 41043 3228 41063 3292
rect 34764 3200 41063 3228
rect 41083 9372 47382 9400
rect 41083 9308 47298 9372
rect 47362 9308 47382 9372
rect 41083 9292 47382 9308
rect 41083 9228 47298 9292
rect 47362 9228 47382 9292
rect 41083 9212 47382 9228
rect 41083 9148 47298 9212
rect 47362 9148 47382 9212
rect 41083 9132 47382 9148
rect 41083 9068 47298 9132
rect 47362 9068 47382 9132
rect 41083 9052 47382 9068
rect 41083 8988 47298 9052
rect 47362 8988 47382 9052
rect 41083 8972 47382 8988
rect 41083 8908 47298 8972
rect 47362 8908 47382 8972
rect 41083 8892 47382 8908
rect 41083 8828 47298 8892
rect 47362 8828 47382 8892
rect 41083 8812 47382 8828
rect 41083 8748 47298 8812
rect 47362 8748 47382 8812
rect 41083 8732 47382 8748
rect 41083 8668 47298 8732
rect 47362 8668 47382 8732
rect 41083 8652 47382 8668
rect 41083 8588 47298 8652
rect 47362 8588 47382 8652
rect 41083 8572 47382 8588
rect 41083 8508 47298 8572
rect 47362 8508 47382 8572
rect 41083 8492 47382 8508
rect 41083 8428 47298 8492
rect 47362 8428 47382 8492
rect 41083 8412 47382 8428
rect 41083 8348 47298 8412
rect 47362 8348 47382 8412
rect 41083 8332 47382 8348
rect 41083 8268 47298 8332
rect 47362 8268 47382 8332
rect 41083 8252 47382 8268
rect 41083 8188 47298 8252
rect 47362 8188 47382 8252
rect 41083 8172 47382 8188
rect 41083 8108 47298 8172
rect 47362 8108 47382 8172
rect 41083 8092 47382 8108
rect 41083 8028 47298 8092
rect 47362 8028 47382 8092
rect 41083 8012 47382 8028
rect 41083 7948 47298 8012
rect 47362 7948 47382 8012
rect 41083 7932 47382 7948
rect 41083 7868 47298 7932
rect 47362 7868 47382 7932
rect 41083 7852 47382 7868
rect 41083 7788 47298 7852
rect 47362 7788 47382 7852
rect 41083 7772 47382 7788
rect 41083 7708 47298 7772
rect 47362 7708 47382 7772
rect 41083 7692 47382 7708
rect 41083 7628 47298 7692
rect 47362 7628 47382 7692
rect 41083 7612 47382 7628
rect 41083 7548 47298 7612
rect 47362 7548 47382 7612
rect 41083 7532 47382 7548
rect 41083 7468 47298 7532
rect 47362 7468 47382 7532
rect 41083 7452 47382 7468
rect 41083 7388 47298 7452
rect 47362 7388 47382 7452
rect 41083 7372 47382 7388
rect 41083 7308 47298 7372
rect 47362 7308 47382 7372
rect 41083 7292 47382 7308
rect 41083 7228 47298 7292
rect 47362 7228 47382 7292
rect 41083 7212 47382 7228
rect 41083 7148 47298 7212
rect 47362 7148 47382 7212
rect 41083 7132 47382 7148
rect 41083 7068 47298 7132
rect 47362 7068 47382 7132
rect 41083 7052 47382 7068
rect 41083 6988 47298 7052
rect 47362 6988 47382 7052
rect 41083 6972 47382 6988
rect 41083 6908 47298 6972
rect 47362 6908 47382 6972
rect 41083 6892 47382 6908
rect 41083 6828 47298 6892
rect 47362 6828 47382 6892
rect 41083 6812 47382 6828
rect 41083 6748 47298 6812
rect 47362 6748 47382 6812
rect 41083 6732 47382 6748
rect 41083 6668 47298 6732
rect 47362 6668 47382 6732
rect 41083 6652 47382 6668
rect 41083 6588 47298 6652
rect 47362 6588 47382 6652
rect 41083 6572 47382 6588
rect 41083 6508 47298 6572
rect 47362 6508 47382 6572
rect 41083 6492 47382 6508
rect 41083 6428 47298 6492
rect 47362 6428 47382 6492
rect 41083 6412 47382 6428
rect 41083 6348 47298 6412
rect 47362 6348 47382 6412
rect 41083 6332 47382 6348
rect 41083 6268 47298 6332
rect 47362 6268 47382 6332
rect 41083 6252 47382 6268
rect 41083 6188 47298 6252
rect 47362 6188 47382 6252
rect 41083 6172 47382 6188
rect 41083 6108 47298 6172
rect 47362 6108 47382 6172
rect 41083 6092 47382 6108
rect 41083 6028 47298 6092
rect 47362 6028 47382 6092
rect 41083 6012 47382 6028
rect 41083 5948 47298 6012
rect 47362 5948 47382 6012
rect 41083 5932 47382 5948
rect 41083 5868 47298 5932
rect 47362 5868 47382 5932
rect 41083 5852 47382 5868
rect 41083 5788 47298 5852
rect 47362 5788 47382 5852
rect 41083 5772 47382 5788
rect 41083 5708 47298 5772
rect 47362 5708 47382 5772
rect 41083 5692 47382 5708
rect 41083 5628 47298 5692
rect 47362 5628 47382 5692
rect 41083 5612 47382 5628
rect 41083 5548 47298 5612
rect 47362 5548 47382 5612
rect 41083 5532 47382 5548
rect 41083 5468 47298 5532
rect 47362 5468 47382 5532
rect 41083 5452 47382 5468
rect 41083 5388 47298 5452
rect 47362 5388 47382 5452
rect 41083 5372 47382 5388
rect 41083 5308 47298 5372
rect 47362 5308 47382 5372
rect 41083 5292 47382 5308
rect 41083 5228 47298 5292
rect 47362 5228 47382 5292
rect 41083 5212 47382 5228
rect 41083 5148 47298 5212
rect 47362 5148 47382 5212
rect 41083 5132 47382 5148
rect 41083 5068 47298 5132
rect 47362 5068 47382 5132
rect 41083 5052 47382 5068
rect 41083 4988 47298 5052
rect 47362 4988 47382 5052
rect 41083 4972 47382 4988
rect 41083 4908 47298 4972
rect 47362 4908 47382 4972
rect 41083 4892 47382 4908
rect 41083 4828 47298 4892
rect 47362 4828 47382 4892
rect 41083 4812 47382 4828
rect 41083 4748 47298 4812
rect 47362 4748 47382 4812
rect 41083 4732 47382 4748
rect 41083 4668 47298 4732
rect 47362 4668 47382 4732
rect 41083 4652 47382 4668
rect 41083 4588 47298 4652
rect 47362 4588 47382 4652
rect 41083 4572 47382 4588
rect 41083 4508 47298 4572
rect 47362 4508 47382 4572
rect 41083 4492 47382 4508
rect 41083 4428 47298 4492
rect 47362 4428 47382 4492
rect 41083 4412 47382 4428
rect 41083 4348 47298 4412
rect 47362 4348 47382 4412
rect 41083 4332 47382 4348
rect 41083 4268 47298 4332
rect 47362 4268 47382 4332
rect 41083 4252 47382 4268
rect 41083 4188 47298 4252
rect 47362 4188 47382 4252
rect 41083 4172 47382 4188
rect 41083 4108 47298 4172
rect 47362 4108 47382 4172
rect 41083 4092 47382 4108
rect 41083 4028 47298 4092
rect 47362 4028 47382 4092
rect 41083 4012 47382 4028
rect 41083 3948 47298 4012
rect 47362 3948 47382 4012
rect 41083 3932 47382 3948
rect 41083 3868 47298 3932
rect 47362 3868 47382 3932
rect 41083 3852 47382 3868
rect 41083 3788 47298 3852
rect 47362 3788 47382 3852
rect 41083 3772 47382 3788
rect 41083 3708 47298 3772
rect 47362 3708 47382 3772
rect 41083 3692 47382 3708
rect 41083 3628 47298 3692
rect 47362 3628 47382 3692
rect 41083 3612 47382 3628
rect 41083 3548 47298 3612
rect 47362 3548 47382 3612
rect 41083 3532 47382 3548
rect 41083 3468 47298 3532
rect 47362 3468 47382 3532
rect 41083 3452 47382 3468
rect 41083 3388 47298 3452
rect 47362 3388 47382 3452
rect 41083 3372 47382 3388
rect 41083 3308 47298 3372
rect 47362 3308 47382 3372
rect 41083 3292 47382 3308
rect 41083 3228 47298 3292
rect 47362 3228 47382 3292
rect 41083 3200 47382 3228
rect -47383 3072 -41084 3100
rect -47383 3008 -41168 3072
rect -41104 3008 -41084 3072
rect -47383 2992 -41084 3008
rect -47383 2928 -41168 2992
rect -41104 2928 -41084 2992
rect -47383 2912 -41084 2928
rect -47383 2848 -41168 2912
rect -41104 2848 -41084 2912
rect -47383 2832 -41084 2848
rect -47383 2768 -41168 2832
rect -41104 2768 -41084 2832
rect -47383 2752 -41084 2768
rect -47383 2688 -41168 2752
rect -41104 2688 -41084 2752
rect -47383 2672 -41084 2688
rect -47383 2608 -41168 2672
rect -41104 2608 -41084 2672
rect -47383 2592 -41084 2608
rect -47383 2528 -41168 2592
rect -41104 2528 -41084 2592
rect -47383 2512 -41084 2528
rect -47383 2448 -41168 2512
rect -41104 2448 -41084 2512
rect -47383 2432 -41084 2448
rect -47383 2368 -41168 2432
rect -41104 2368 -41084 2432
rect -47383 2352 -41084 2368
rect -47383 2288 -41168 2352
rect -41104 2288 -41084 2352
rect -47383 2272 -41084 2288
rect -47383 2208 -41168 2272
rect -41104 2208 -41084 2272
rect -47383 2192 -41084 2208
rect -47383 2128 -41168 2192
rect -41104 2128 -41084 2192
rect -47383 2112 -41084 2128
rect -47383 2048 -41168 2112
rect -41104 2048 -41084 2112
rect -47383 2032 -41084 2048
rect -47383 1968 -41168 2032
rect -41104 1968 -41084 2032
rect -47383 1952 -41084 1968
rect -47383 1888 -41168 1952
rect -41104 1888 -41084 1952
rect -47383 1872 -41084 1888
rect -47383 1808 -41168 1872
rect -41104 1808 -41084 1872
rect -47383 1792 -41084 1808
rect -47383 1728 -41168 1792
rect -41104 1728 -41084 1792
rect -47383 1712 -41084 1728
rect -47383 1648 -41168 1712
rect -41104 1648 -41084 1712
rect -47383 1632 -41084 1648
rect -47383 1568 -41168 1632
rect -41104 1568 -41084 1632
rect -47383 1552 -41084 1568
rect -47383 1488 -41168 1552
rect -41104 1488 -41084 1552
rect -47383 1472 -41084 1488
rect -47383 1408 -41168 1472
rect -41104 1408 -41084 1472
rect -47383 1392 -41084 1408
rect -47383 1328 -41168 1392
rect -41104 1328 -41084 1392
rect -47383 1312 -41084 1328
rect -47383 1248 -41168 1312
rect -41104 1248 -41084 1312
rect -47383 1232 -41084 1248
rect -47383 1168 -41168 1232
rect -41104 1168 -41084 1232
rect -47383 1152 -41084 1168
rect -47383 1088 -41168 1152
rect -41104 1088 -41084 1152
rect -47383 1072 -41084 1088
rect -47383 1008 -41168 1072
rect -41104 1008 -41084 1072
rect -47383 992 -41084 1008
rect -47383 928 -41168 992
rect -41104 928 -41084 992
rect -47383 912 -41084 928
rect -47383 848 -41168 912
rect -41104 848 -41084 912
rect -47383 832 -41084 848
rect -47383 768 -41168 832
rect -41104 768 -41084 832
rect -47383 752 -41084 768
rect -47383 688 -41168 752
rect -41104 688 -41084 752
rect -47383 672 -41084 688
rect -47383 608 -41168 672
rect -41104 608 -41084 672
rect -47383 592 -41084 608
rect -47383 528 -41168 592
rect -41104 528 -41084 592
rect -47383 512 -41084 528
rect -47383 448 -41168 512
rect -41104 448 -41084 512
rect -47383 432 -41084 448
rect -47383 368 -41168 432
rect -41104 368 -41084 432
rect -47383 352 -41084 368
rect -47383 288 -41168 352
rect -41104 288 -41084 352
rect -47383 272 -41084 288
rect -47383 208 -41168 272
rect -41104 208 -41084 272
rect -47383 192 -41084 208
rect -47383 128 -41168 192
rect -41104 128 -41084 192
rect -47383 112 -41084 128
rect -47383 48 -41168 112
rect -41104 48 -41084 112
rect -47383 32 -41084 48
rect -47383 -32 -41168 32
rect -41104 -32 -41084 32
rect -47383 -48 -41084 -32
rect -47383 -112 -41168 -48
rect -41104 -112 -41084 -48
rect -47383 -128 -41084 -112
rect -47383 -192 -41168 -128
rect -41104 -192 -41084 -128
rect -47383 -208 -41084 -192
rect -47383 -272 -41168 -208
rect -41104 -272 -41084 -208
rect -47383 -288 -41084 -272
rect -47383 -352 -41168 -288
rect -41104 -352 -41084 -288
rect -47383 -368 -41084 -352
rect -47383 -432 -41168 -368
rect -41104 -432 -41084 -368
rect -47383 -448 -41084 -432
rect -47383 -512 -41168 -448
rect -41104 -512 -41084 -448
rect -47383 -528 -41084 -512
rect -47383 -592 -41168 -528
rect -41104 -592 -41084 -528
rect -47383 -608 -41084 -592
rect -47383 -672 -41168 -608
rect -41104 -672 -41084 -608
rect -47383 -688 -41084 -672
rect -47383 -752 -41168 -688
rect -41104 -752 -41084 -688
rect -47383 -768 -41084 -752
rect -47383 -832 -41168 -768
rect -41104 -832 -41084 -768
rect -47383 -848 -41084 -832
rect -47383 -912 -41168 -848
rect -41104 -912 -41084 -848
rect -47383 -928 -41084 -912
rect -47383 -992 -41168 -928
rect -41104 -992 -41084 -928
rect -47383 -1008 -41084 -992
rect -47383 -1072 -41168 -1008
rect -41104 -1072 -41084 -1008
rect -47383 -1088 -41084 -1072
rect -47383 -1152 -41168 -1088
rect -41104 -1152 -41084 -1088
rect -47383 -1168 -41084 -1152
rect -47383 -1232 -41168 -1168
rect -41104 -1232 -41084 -1168
rect -47383 -1248 -41084 -1232
rect -47383 -1312 -41168 -1248
rect -41104 -1312 -41084 -1248
rect -47383 -1328 -41084 -1312
rect -47383 -1392 -41168 -1328
rect -41104 -1392 -41084 -1328
rect -47383 -1408 -41084 -1392
rect -47383 -1472 -41168 -1408
rect -41104 -1472 -41084 -1408
rect -47383 -1488 -41084 -1472
rect -47383 -1552 -41168 -1488
rect -41104 -1552 -41084 -1488
rect -47383 -1568 -41084 -1552
rect -47383 -1632 -41168 -1568
rect -41104 -1632 -41084 -1568
rect -47383 -1648 -41084 -1632
rect -47383 -1712 -41168 -1648
rect -41104 -1712 -41084 -1648
rect -47383 -1728 -41084 -1712
rect -47383 -1792 -41168 -1728
rect -41104 -1792 -41084 -1728
rect -47383 -1808 -41084 -1792
rect -47383 -1872 -41168 -1808
rect -41104 -1872 -41084 -1808
rect -47383 -1888 -41084 -1872
rect -47383 -1952 -41168 -1888
rect -41104 -1952 -41084 -1888
rect -47383 -1968 -41084 -1952
rect -47383 -2032 -41168 -1968
rect -41104 -2032 -41084 -1968
rect -47383 -2048 -41084 -2032
rect -47383 -2112 -41168 -2048
rect -41104 -2112 -41084 -2048
rect -47383 -2128 -41084 -2112
rect -47383 -2192 -41168 -2128
rect -41104 -2192 -41084 -2128
rect -47383 -2208 -41084 -2192
rect -47383 -2272 -41168 -2208
rect -41104 -2272 -41084 -2208
rect -47383 -2288 -41084 -2272
rect -47383 -2352 -41168 -2288
rect -41104 -2352 -41084 -2288
rect -47383 -2368 -41084 -2352
rect -47383 -2432 -41168 -2368
rect -41104 -2432 -41084 -2368
rect -47383 -2448 -41084 -2432
rect -47383 -2512 -41168 -2448
rect -41104 -2512 -41084 -2448
rect -47383 -2528 -41084 -2512
rect -47383 -2592 -41168 -2528
rect -41104 -2592 -41084 -2528
rect -47383 -2608 -41084 -2592
rect -47383 -2672 -41168 -2608
rect -41104 -2672 -41084 -2608
rect -47383 -2688 -41084 -2672
rect -47383 -2752 -41168 -2688
rect -41104 -2752 -41084 -2688
rect -47383 -2768 -41084 -2752
rect -47383 -2832 -41168 -2768
rect -41104 -2832 -41084 -2768
rect -47383 -2848 -41084 -2832
rect -47383 -2912 -41168 -2848
rect -41104 -2912 -41084 -2848
rect -47383 -2928 -41084 -2912
rect -47383 -2992 -41168 -2928
rect -41104 -2992 -41084 -2928
rect -47383 -3008 -41084 -2992
rect -47383 -3072 -41168 -3008
rect -41104 -3072 -41084 -3008
rect -47383 -3100 -41084 -3072
rect -41064 3072 -34765 3100
rect -41064 3008 -34849 3072
rect -34785 3008 -34765 3072
rect -41064 2992 -34765 3008
rect -41064 2928 -34849 2992
rect -34785 2928 -34765 2992
rect -41064 2912 -34765 2928
rect -41064 2848 -34849 2912
rect -34785 2848 -34765 2912
rect -41064 2832 -34765 2848
rect -41064 2768 -34849 2832
rect -34785 2768 -34765 2832
rect -41064 2752 -34765 2768
rect -41064 2688 -34849 2752
rect -34785 2688 -34765 2752
rect -41064 2672 -34765 2688
rect -41064 2608 -34849 2672
rect -34785 2608 -34765 2672
rect -41064 2592 -34765 2608
rect -41064 2528 -34849 2592
rect -34785 2528 -34765 2592
rect -41064 2512 -34765 2528
rect -41064 2448 -34849 2512
rect -34785 2448 -34765 2512
rect -41064 2432 -34765 2448
rect -41064 2368 -34849 2432
rect -34785 2368 -34765 2432
rect -41064 2352 -34765 2368
rect -41064 2288 -34849 2352
rect -34785 2288 -34765 2352
rect -41064 2272 -34765 2288
rect -41064 2208 -34849 2272
rect -34785 2208 -34765 2272
rect -41064 2192 -34765 2208
rect -41064 2128 -34849 2192
rect -34785 2128 -34765 2192
rect -41064 2112 -34765 2128
rect -41064 2048 -34849 2112
rect -34785 2048 -34765 2112
rect -41064 2032 -34765 2048
rect -41064 1968 -34849 2032
rect -34785 1968 -34765 2032
rect -41064 1952 -34765 1968
rect -41064 1888 -34849 1952
rect -34785 1888 -34765 1952
rect -41064 1872 -34765 1888
rect -41064 1808 -34849 1872
rect -34785 1808 -34765 1872
rect -41064 1792 -34765 1808
rect -41064 1728 -34849 1792
rect -34785 1728 -34765 1792
rect -41064 1712 -34765 1728
rect -41064 1648 -34849 1712
rect -34785 1648 -34765 1712
rect -41064 1632 -34765 1648
rect -41064 1568 -34849 1632
rect -34785 1568 -34765 1632
rect -41064 1552 -34765 1568
rect -41064 1488 -34849 1552
rect -34785 1488 -34765 1552
rect -41064 1472 -34765 1488
rect -41064 1408 -34849 1472
rect -34785 1408 -34765 1472
rect -41064 1392 -34765 1408
rect -41064 1328 -34849 1392
rect -34785 1328 -34765 1392
rect -41064 1312 -34765 1328
rect -41064 1248 -34849 1312
rect -34785 1248 -34765 1312
rect -41064 1232 -34765 1248
rect -41064 1168 -34849 1232
rect -34785 1168 -34765 1232
rect -41064 1152 -34765 1168
rect -41064 1088 -34849 1152
rect -34785 1088 -34765 1152
rect -41064 1072 -34765 1088
rect -41064 1008 -34849 1072
rect -34785 1008 -34765 1072
rect -41064 992 -34765 1008
rect -41064 928 -34849 992
rect -34785 928 -34765 992
rect -41064 912 -34765 928
rect -41064 848 -34849 912
rect -34785 848 -34765 912
rect -41064 832 -34765 848
rect -41064 768 -34849 832
rect -34785 768 -34765 832
rect -41064 752 -34765 768
rect -41064 688 -34849 752
rect -34785 688 -34765 752
rect -41064 672 -34765 688
rect -41064 608 -34849 672
rect -34785 608 -34765 672
rect -41064 592 -34765 608
rect -41064 528 -34849 592
rect -34785 528 -34765 592
rect -41064 512 -34765 528
rect -41064 448 -34849 512
rect -34785 448 -34765 512
rect -41064 432 -34765 448
rect -41064 368 -34849 432
rect -34785 368 -34765 432
rect -41064 352 -34765 368
rect -41064 288 -34849 352
rect -34785 288 -34765 352
rect -41064 272 -34765 288
rect -41064 208 -34849 272
rect -34785 208 -34765 272
rect -41064 192 -34765 208
rect -41064 128 -34849 192
rect -34785 128 -34765 192
rect -41064 112 -34765 128
rect -41064 48 -34849 112
rect -34785 48 -34765 112
rect -41064 32 -34765 48
rect -41064 -32 -34849 32
rect -34785 -32 -34765 32
rect -41064 -48 -34765 -32
rect -41064 -112 -34849 -48
rect -34785 -112 -34765 -48
rect -41064 -128 -34765 -112
rect -41064 -192 -34849 -128
rect -34785 -192 -34765 -128
rect -41064 -208 -34765 -192
rect -41064 -272 -34849 -208
rect -34785 -272 -34765 -208
rect -41064 -288 -34765 -272
rect -41064 -352 -34849 -288
rect -34785 -352 -34765 -288
rect -41064 -368 -34765 -352
rect -41064 -432 -34849 -368
rect -34785 -432 -34765 -368
rect -41064 -448 -34765 -432
rect -41064 -512 -34849 -448
rect -34785 -512 -34765 -448
rect -41064 -528 -34765 -512
rect -41064 -592 -34849 -528
rect -34785 -592 -34765 -528
rect -41064 -608 -34765 -592
rect -41064 -672 -34849 -608
rect -34785 -672 -34765 -608
rect -41064 -688 -34765 -672
rect -41064 -752 -34849 -688
rect -34785 -752 -34765 -688
rect -41064 -768 -34765 -752
rect -41064 -832 -34849 -768
rect -34785 -832 -34765 -768
rect -41064 -848 -34765 -832
rect -41064 -912 -34849 -848
rect -34785 -912 -34765 -848
rect -41064 -928 -34765 -912
rect -41064 -992 -34849 -928
rect -34785 -992 -34765 -928
rect -41064 -1008 -34765 -992
rect -41064 -1072 -34849 -1008
rect -34785 -1072 -34765 -1008
rect -41064 -1088 -34765 -1072
rect -41064 -1152 -34849 -1088
rect -34785 -1152 -34765 -1088
rect -41064 -1168 -34765 -1152
rect -41064 -1232 -34849 -1168
rect -34785 -1232 -34765 -1168
rect -41064 -1248 -34765 -1232
rect -41064 -1312 -34849 -1248
rect -34785 -1312 -34765 -1248
rect -41064 -1328 -34765 -1312
rect -41064 -1392 -34849 -1328
rect -34785 -1392 -34765 -1328
rect -41064 -1408 -34765 -1392
rect -41064 -1472 -34849 -1408
rect -34785 -1472 -34765 -1408
rect -41064 -1488 -34765 -1472
rect -41064 -1552 -34849 -1488
rect -34785 -1552 -34765 -1488
rect -41064 -1568 -34765 -1552
rect -41064 -1632 -34849 -1568
rect -34785 -1632 -34765 -1568
rect -41064 -1648 -34765 -1632
rect -41064 -1712 -34849 -1648
rect -34785 -1712 -34765 -1648
rect -41064 -1728 -34765 -1712
rect -41064 -1792 -34849 -1728
rect -34785 -1792 -34765 -1728
rect -41064 -1808 -34765 -1792
rect -41064 -1872 -34849 -1808
rect -34785 -1872 -34765 -1808
rect -41064 -1888 -34765 -1872
rect -41064 -1952 -34849 -1888
rect -34785 -1952 -34765 -1888
rect -41064 -1968 -34765 -1952
rect -41064 -2032 -34849 -1968
rect -34785 -2032 -34765 -1968
rect -41064 -2048 -34765 -2032
rect -41064 -2112 -34849 -2048
rect -34785 -2112 -34765 -2048
rect -41064 -2128 -34765 -2112
rect -41064 -2192 -34849 -2128
rect -34785 -2192 -34765 -2128
rect -41064 -2208 -34765 -2192
rect -41064 -2272 -34849 -2208
rect -34785 -2272 -34765 -2208
rect -41064 -2288 -34765 -2272
rect -41064 -2352 -34849 -2288
rect -34785 -2352 -34765 -2288
rect -41064 -2368 -34765 -2352
rect -41064 -2432 -34849 -2368
rect -34785 -2432 -34765 -2368
rect -41064 -2448 -34765 -2432
rect -41064 -2512 -34849 -2448
rect -34785 -2512 -34765 -2448
rect -41064 -2528 -34765 -2512
rect -41064 -2592 -34849 -2528
rect -34785 -2592 -34765 -2528
rect -41064 -2608 -34765 -2592
rect -41064 -2672 -34849 -2608
rect -34785 -2672 -34765 -2608
rect -41064 -2688 -34765 -2672
rect -41064 -2752 -34849 -2688
rect -34785 -2752 -34765 -2688
rect -41064 -2768 -34765 -2752
rect -41064 -2832 -34849 -2768
rect -34785 -2832 -34765 -2768
rect -41064 -2848 -34765 -2832
rect -41064 -2912 -34849 -2848
rect -34785 -2912 -34765 -2848
rect -41064 -2928 -34765 -2912
rect -41064 -2992 -34849 -2928
rect -34785 -2992 -34765 -2928
rect -41064 -3008 -34765 -2992
rect -41064 -3072 -34849 -3008
rect -34785 -3072 -34765 -3008
rect -41064 -3100 -34765 -3072
rect -34745 3072 -28446 3100
rect -34745 3008 -28530 3072
rect -28466 3008 -28446 3072
rect -34745 2992 -28446 3008
rect -34745 2928 -28530 2992
rect -28466 2928 -28446 2992
rect -34745 2912 -28446 2928
rect -34745 2848 -28530 2912
rect -28466 2848 -28446 2912
rect -34745 2832 -28446 2848
rect -34745 2768 -28530 2832
rect -28466 2768 -28446 2832
rect -34745 2752 -28446 2768
rect -34745 2688 -28530 2752
rect -28466 2688 -28446 2752
rect -34745 2672 -28446 2688
rect -34745 2608 -28530 2672
rect -28466 2608 -28446 2672
rect -34745 2592 -28446 2608
rect -34745 2528 -28530 2592
rect -28466 2528 -28446 2592
rect -34745 2512 -28446 2528
rect -34745 2448 -28530 2512
rect -28466 2448 -28446 2512
rect -34745 2432 -28446 2448
rect -34745 2368 -28530 2432
rect -28466 2368 -28446 2432
rect -34745 2352 -28446 2368
rect -34745 2288 -28530 2352
rect -28466 2288 -28446 2352
rect -34745 2272 -28446 2288
rect -34745 2208 -28530 2272
rect -28466 2208 -28446 2272
rect -34745 2192 -28446 2208
rect -34745 2128 -28530 2192
rect -28466 2128 -28446 2192
rect -34745 2112 -28446 2128
rect -34745 2048 -28530 2112
rect -28466 2048 -28446 2112
rect -34745 2032 -28446 2048
rect -34745 1968 -28530 2032
rect -28466 1968 -28446 2032
rect -34745 1952 -28446 1968
rect -34745 1888 -28530 1952
rect -28466 1888 -28446 1952
rect -34745 1872 -28446 1888
rect -34745 1808 -28530 1872
rect -28466 1808 -28446 1872
rect -34745 1792 -28446 1808
rect -34745 1728 -28530 1792
rect -28466 1728 -28446 1792
rect -34745 1712 -28446 1728
rect -34745 1648 -28530 1712
rect -28466 1648 -28446 1712
rect -34745 1632 -28446 1648
rect -34745 1568 -28530 1632
rect -28466 1568 -28446 1632
rect -34745 1552 -28446 1568
rect -34745 1488 -28530 1552
rect -28466 1488 -28446 1552
rect -34745 1472 -28446 1488
rect -34745 1408 -28530 1472
rect -28466 1408 -28446 1472
rect -34745 1392 -28446 1408
rect -34745 1328 -28530 1392
rect -28466 1328 -28446 1392
rect -34745 1312 -28446 1328
rect -34745 1248 -28530 1312
rect -28466 1248 -28446 1312
rect -34745 1232 -28446 1248
rect -34745 1168 -28530 1232
rect -28466 1168 -28446 1232
rect -34745 1152 -28446 1168
rect -34745 1088 -28530 1152
rect -28466 1088 -28446 1152
rect -34745 1072 -28446 1088
rect -34745 1008 -28530 1072
rect -28466 1008 -28446 1072
rect -34745 992 -28446 1008
rect -34745 928 -28530 992
rect -28466 928 -28446 992
rect -34745 912 -28446 928
rect -34745 848 -28530 912
rect -28466 848 -28446 912
rect -34745 832 -28446 848
rect -34745 768 -28530 832
rect -28466 768 -28446 832
rect -34745 752 -28446 768
rect -34745 688 -28530 752
rect -28466 688 -28446 752
rect -34745 672 -28446 688
rect -34745 608 -28530 672
rect -28466 608 -28446 672
rect -34745 592 -28446 608
rect -34745 528 -28530 592
rect -28466 528 -28446 592
rect -34745 512 -28446 528
rect -34745 448 -28530 512
rect -28466 448 -28446 512
rect -34745 432 -28446 448
rect -34745 368 -28530 432
rect -28466 368 -28446 432
rect -34745 352 -28446 368
rect -34745 288 -28530 352
rect -28466 288 -28446 352
rect -34745 272 -28446 288
rect -34745 208 -28530 272
rect -28466 208 -28446 272
rect -34745 192 -28446 208
rect -34745 128 -28530 192
rect -28466 128 -28446 192
rect -34745 112 -28446 128
rect -34745 48 -28530 112
rect -28466 48 -28446 112
rect -34745 32 -28446 48
rect -34745 -32 -28530 32
rect -28466 -32 -28446 32
rect -34745 -48 -28446 -32
rect -34745 -112 -28530 -48
rect -28466 -112 -28446 -48
rect -34745 -128 -28446 -112
rect -34745 -192 -28530 -128
rect -28466 -192 -28446 -128
rect -34745 -208 -28446 -192
rect -34745 -272 -28530 -208
rect -28466 -272 -28446 -208
rect -34745 -288 -28446 -272
rect -34745 -352 -28530 -288
rect -28466 -352 -28446 -288
rect -34745 -368 -28446 -352
rect -34745 -432 -28530 -368
rect -28466 -432 -28446 -368
rect -34745 -448 -28446 -432
rect -34745 -512 -28530 -448
rect -28466 -512 -28446 -448
rect -34745 -528 -28446 -512
rect -34745 -592 -28530 -528
rect -28466 -592 -28446 -528
rect -34745 -608 -28446 -592
rect -34745 -672 -28530 -608
rect -28466 -672 -28446 -608
rect -34745 -688 -28446 -672
rect -34745 -752 -28530 -688
rect -28466 -752 -28446 -688
rect -34745 -768 -28446 -752
rect -34745 -832 -28530 -768
rect -28466 -832 -28446 -768
rect -34745 -848 -28446 -832
rect -34745 -912 -28530 -848
rect -28466 -912 -28446 -848
rect -34745 -928 -28446 -912
rect -34745 -992 -28530 -928
rect -28466 -992 -28446 -928
rect -34745 -1008 -28446 -992
rect -34745 -1072 -28530 -1008
rect -28466 -1072 -28446 -1008
rect -34745 -1088 -28446 -1072
rect -34745 -1152 -28530 -1088
rect -28466 -1152 -28446 -1088
rect -34745 -1168 -28446 -1152
rect -34745 -1232 -28530 -1168
rect -28466 -1232 -28446 -1168
rect -34745 -1248 -28446 -1232
rect -34745 -1312 -28530 -1248
rect -28466 -1312 -28446 -1248
rect -34745 -1328 -28446 -1312
rect -34745 -1392 -28530 -1328
rect -28466 -1392 -28446 -1328
rect -34745 -1408 -28446 -1392
rect -34745 -1472 -28530 -1408
rect -28466 -1472 -28446 -1408
rect -34745 -1488 -28446 -1472
rect -34745 -1552 -28530 -1488
rect -28466 -1552 -28446 -1488
rect -34745 -1568 -28446 -1552
rect -34745 -1632 -28530 -1568
rect -28466 -1632 -28446 -1568
rect -34745 -1648 -28446 -1632
rect -34745 -1712 -28530 -1648
rect -28466 -1712 -28446 -1648
rect -34745 -1728 -28446 -1712
rect -34745 -1792 -28530 -1728
rect -28466 -1792 -28446 -1728
rect -34745 -1808 -28446 -1792
rect -34745 -1872 -28530 -1808
rect -28466 -1872 -28446 -1808
rect -34745 -1888 -28446 -1872
rect -34745 -1952 -28530 -1888
rect -28466 -1952 -28446 -1888
rect -34745 -1968 -28446 -1952
rect -34745 -2032 -28530 -1968
rect -28466 -2032 -28446 -1968
rect -34745 -2048 -28446 -2032
rect -34745 -2112 -28530 -2048
rect -28466 -2112 -28446 -2048
rect -34745 -2128 -28446 -2112
rect -34745 -2192 -28530 -2128
rect -28466 -2192 -28446 -2128
rect -34745 -2208 -28446 -2192
rect -34745 -2272 -28530 -2208
rect -28466 -2272 -28446 -2208
rect -34745 -2288 -28446 -2272
rect -34745 -2352 -28530 -2288
rect -28466 -2352 -28446 -2288
rect -34745 -2368 -28446 -2352
rect -34745 -2432 -28530 -2368
rect -28466 -2432 -28446 -2368
rect -34745 -2448 -28446 -2432
rect -34745 -2512 -28530 -2448
rect -28466 -2512 -28446 -2448
rect -34745 -2528 -28446 -2512
rect -34745 -2592 -28530 -2528
rect -28466 -2592 -28446 -2528
rect -34745 -2608 -28446 -2592
rect -34745 -2672 -28530 -2608
rect -28466 -2672 -28446 -2608
rect -34745 -2688 -28446 -2672
rect -34745 -2752 -28530 -2688
rect -28466 -2752 -28446 -2688
rect -34745 -2768 -28446 -2752
rect -34745 -2832 -28530 -2768
rect -28466 -2832 -28446 -2768
rect -34745 -2848 -28446 -2832
rect -34745 -2912 -28530 -2848
rect -28466 -2912 -28446 -2848
rect -34745 -2928 -28446 -2912
rect -34745 -2992 -28530 -2928
rect -28466 -2992 -28446 -2928
rect -34745 -3008 -28446 -2992
rect -34745 -3072 -28530 -3008
rect -28466 -3072 -28446 -3008
rect -34745 -3100 -28446 -3072
rect -28426 3072 -22127 3100
rect -28426 3008 -22211 3072
rect -22147 3008 -22127 3072
rect -28426 2992 -22127 3008
rect -28426 2928 -22211 2992
rect -22147 2928 -22127 2992
rect -28426 2912 -22127 2928
rect -28426 2848 -22211 2912
rect -22147 2848 -22127 2912
rect -28426 2832 -22127 2848
rect -28426 2768 -22211 2832
rect -22147 2768 -22127 2832
rect -28426 2752 -22127 2768
rect -28426 2688 -22211 2752
rect -22147 2688 -22127 2752
rect -28426 2672 -22127 2688
rect -28426 2608 -22211 2672
rect -22147 2608 -22127 2672
rect -28426 2592 -22127 2608
rect -28426 2528 -22211 2592
rect -22147 2528 -22127 2592
rect -28426 2512 -22127 2528
rect -28426 2448 -22211 2512
rect -22147 2448 -22127 2512
rect -28426 2432 -22127 2448
rect -28426 2368 -22211 2432
rect -22147 2368 -22127 2432
rect -28426 2352 -22127 2368
rect -28426 2288 -22211 2352
rect -22147 2288 -22127 2352
rect -28426 2272 -22127 2288
rect -28426 2208 -22211 2272
rect -22147 2208 -22127 2272
rect -28426 2192 -22127 2208
rect -28426 2128 -22211 2192
rect -22147 2128 -22127 2192
rect -28426 2112 -22127 2128
rect -28426 2048 -22211 2112
rect -22147 2048 -22127 2112
rect -28426 2032 -22127 2048
rect -28426 1968 -22211 2032
rect -22147 1968 -22127 2032
rect -28426 1952 -22127 1968
rect -28426 1888 -22211 1952
rect -22147 1888 -22127 1952
rect -28426 1872 -22127 1888
rect -28426 1808 -22211 1872
rect -22147 1808 -22127 1872
rect -28426 1792 -22127 1808
rect -28426 1728 -22211 1792
rect -22147 1728 -22127 1792
rect -28426 1712 -22127 1728
rect -28426 1648 -22211 1712
rect -22147 1648 -22127 1712
rect -28426 1632 -22127 1648
rect -28426 1568 -22211 1632
rect -22147 1568 -22127 1632
rect -28426 1552 -22127 1568
rect -28426 1488 -22211 1552
rect -22147 1488 -22127 1552
rect -28426 1472 -22127 1488
rect -28426 1408 -22211 1472
rect -22147 1408 -22127 1472
rect -28426 1392 -22127 1408
rect -28426 1328 -22211 1392
rect -22147 1328 -22127 1392
rect -28426 1312 -22127 1328
rect -28426 1248 -22211 1312
rect -22147 1248 -22127 1312
rect -28426 1232 -22127 1248
rect -28426 1168 -22211 1232
rect -22147 1168 -22127 1232
rect -28426 1152 -22127 1168
rect -28426 1088 -22211 1152
rect -22147 1088 -22127 1152
rect -28426 1072 -22127 1088
rect -28426 1008 -22211 1072
rect -22147 1008 -22127 1072
rect -28426 992 -22127 1008
rect -28426 928 -22211 992
rect -22147 928 -22127 992
rect -28426 912 -22127 928
rect -28426 848 -22211 912
rect -22147 848 -22127 912
rect -28426 832 -22127 848
rect -28426 768 -22211 832
rect -22147 768 -22127 832
rect -28426 752 -22127 768
rect -28426 688 -22211 752
rect -22147 688 -22127 752
rect -28426 672 -22127 688
rect -28426 608 -22211 672
rect -22147 608 -22127 672
rect -28426 592 -22127 608
rect -28426 528 -22211 592
rect -22147 528 -22127 592
rect -28426 512 -22127 528
rect -28426 448 -22211 512
rect -22147 448 -22127 512
rect -28426 432 -22127 448
rect -28426 368 -22211 432
rect -22147 368 -22127 432
rect -28426 352 -22127 368
rect -28426 288 -22211 352
rect -22147 288 -22127 352
rect -28426 272 -22127 288
rect -28426 208 -22211 272
rect -22147 208 -22127 272
rect -28426 192 -22127 208
rect -28426 128 -22211 192
rect -22147 128 -22127 192
rect -28426 112 -22127 128
rect -28426 48 -22211 112
rect -22147 48 -22127 112
rect -28426 32 -22127 48
rect -28426 -32 -22211 32
rect -22147 -32 -22127 32
rect -28426 -48 -22127 -32
rect -28426 -112 -22211 -48
rect -22147 -112 -22127 -48
rect -28426 -128 -22127 -112
rect -28426 -192 -22211 -128
rect -22147 -192 -22127 -128
rect -28426 -208 -22127 -192
rect -28426 -272 -22211 -208
rect -22147 -272 -22127 -208
rect -28426 -288 -22127 -272
rect -28426 -352 -22211 -288
rect -22147 -352 -22127 -288
rect -28426 -368 -22127 -352
rect -28426 -432 -22211 -368
rect -22147 -432 -22127 -368
rect -28426 -448 -22127 -432
rect -28426 -512 -22211 -448
rect -22147 -512 -22127 -448
rect -28426 -528 -22127 -512
rect -28426 -592 -22211 -528
rect -22147 -592 -22127 -528
rect -28426 -608 -22127 -592
rect -28426 -672 -22211 -608
rect -22147 -672 -22127 -608
rect -28426 -688 -22127 -672
rect -28426 -752 -22211 -688
rect -22147 -752 -22127 -688
rect -28426 -768 -22127 -752
rect -28426 -832 -22211 -768
rect -22147 -832 -22127 -768
rect -28426 -848 -22127 -832
rect -28426 -912 -22211 -848
rect -22147 -912 -22127 -848
rect -28426 -928 -22127 -912
rect -28426 -992 -22211 -928
rect -22147 -992 -22127 -928
rect -28426 -1008 -22127 -992
rect -28426 -1072 -22211 -1008
rect -22147 -1072 -22127 -1008
rect -28426 -1088 -22127 -1072
rect -28426 -1152 -22211 -1088
rect -22147 -1152 -22127 -1088
rect -28426 -1168 -22127 -1152
rect -28426 -1232 -22211 -1168
rect -22147 -1232 -22127 -1168
rect -28426 -1248 -22127 -1232
rect -28426 -1312 -22211 -1248
rect -22147 -1312 -22127 -1248
rect -28426 -1328 -22127 -1312
rect -28426 -1392 -22211 -1328
rect -22147 -1392 -22127 -1328
rect -28426 -1408 -22127 -1392
rect -28426 -1472 -22211 -1408
rect -22147 -1472 -22127 -1408
rect -28426 -1488 -22127 -1472
rect -28426 -1552 -22211 -1488
rect -22147 -1552 -22127 -1488
rect -28426 -1568 -22127 -1552
rect -28426 -1632 -22211 -1568
rect -22147 -1632 -22127 -1568
rect -28426 -1648 -22127 -1632
rect -28426 -1712 -22211 -1648
rect -22147 -1712 -22127 -1648
rect -28426 -1728 -22127 -1712
rect -28426 -1792 -22211 -1728
rect -22147 -1792 -22127 -1728
rect -28426 -1808 -22127 -1792
rect -28426 -1872 -22211 -1808
rect -22147 -1872 -22127 -1808
rect -28426 -1888 -22127 -1872
rect -28426 -1952 -22211 -1888
rect -22147 -1952 -22127 -1888
rect -28426 -1968 -22127 -1952
rect -28426 -2032 -22211 -1968
rect -22147 -2032 -22127 -1968
rect -28426 -2048 -22127 -2032
rect -28426 -2112 -22211 -2048
rect -22147 -2112 -22127 -2048
rect -28426 -2128 -22127 -2112
rect -28426 -2192 -22211 -2128
rect -22147 -2192 -22127 -2128
rect -28426 -2208 -22127 -2192
rect -28426 -2272 -22211 -2208
rect -22147 -2272 -22127 -2208
rect -28426 -2288 -22127 -2272
rect -28426 -2352 -22211 -2288
rect -22147 -2352 -22127 -2288
rect -28426 -2368 -22127 -2352
rect -28426 -2432 -22211 -2368
rect -22147 -2432 -22127 -2368
rect -28426 -2448 -22127 -2432
rect -28426 -2512 -22211 -2448
rect -22147 -2512 -22127 -2448
rect -28426 -2528 -22127 -2512
rect -28426 -2592 -22211 -2528
rect -22147 -2592 -22127 -2528
rect -28426 -2608 -22127 -2592
rect -28426 -2672 -22211 -2608
rect -22147 -2672 -22127 -2608
rect -28426 -2688 -22127 -2672
rect -28426 -2752 -22211 -2688
rect -22147 -2752 -22127 -2688
rect -28426 -2768 -22127 -2752
rect -28426 -2832 -22211 -2768
rect -22147 -2832 -22127 -2768
rect -28426 -2848 -22127 -2832
rect -28426 -2912 -22211 -2848
rect -22147 -2912 -22127 -2848
rect -28426 -2928 -22127 -2912
rect -28426 -2992 -22211 -2928
rect -22147 -2992 -22127 -2928
rect -28426 -3008 -22127 -2992
rect -28426 -3072 -22211 -3008
rect -22147 -3072 -22127 -3008
rect -28426 -3100 -22127 -3072
rect -22107 3072 -15808 3100
rect -22107 3008 -15892 3072
rect -15828 3008 -15808 3072
rect -22107 2992 -15808 3008
rect -22107 2928 -15892 2992
rect -15828 2928 -15808 2992
rect -22107 2912 -15808 2928
rect -22107 2848 -15892 2912
rect -15828 2848 -15808 2912
rect -22107 2832 -15808 2848
rect -22107 2768 -15892 2832
rect -15828 2768 -15808 2832
rect -22107 2752 -15808 2768
rect -22107 2688 -15892 2752
rect -15828 2688 -15808 2752
rect -22107 2672 -15808 2688
rect -22107 2608 -15892 2672
rect -15828 2608 -15808 2672
rect -22107 2592 -15808 2608
rect -22107 2528 -15892 2592
rect -15828 2528 -15808 2592
rect -22107 2512 -15808 2528
rect -22107 2448 -15892 2512
rect -15828 2448 -15808 2512
rect -22107 2432 -15808 2448
rect -22107 2368 -15892 2432
rect -15828 2368 -15808 2432
rect -22107 2352 -15808 2368
rect -22107 2288 -15892 2352
rect -15828 2288 -15808 2352
rect -22107 2272 -15808 2288
rect -22107 2208 -15892 2272
rect -15828 2208 -15808 2272
rect -22107 2192 -15808 2208
rect -22107 2128 -15892 2192
rect -15828 2128 -15808 2192
rect -22107 2112 -15808 2128
rect -22107 2048 -15892 2112
rect -15828 2048 -15808 2112
rect -22107 2032 -15808 2048
rect -22107 1968 -15892 2032
rect -15828 1968 -15808 2032
rect -22107 1952 -15808 1968
rect -22107 1888 -15892 1952
rect -15828 1888 -15808 1952
rect -22107 1872 -15808 1888
rect -22107 1808 -15892 1872
rect -15828 1808 -15808 1872
rect -22107 1792 -15808 1808
rect -22107 1728 -15892 1792
rect -15828 1728 -15808 1792
rect -22107 1712 -15808 1728
rect -22107 1648 -15892 1712
rect -15828 1648 -15808 1712
rect -22107 1632 -15808 1648
rect -22107 1568 -15892 1632
rect -15828 1568 -15808 1632
rect -22107 1552 -15808 1568
rect -22107 1488 -15892 1552
rect -15828 1488 -15808 1552
rect -22107 1472 -15808 1488
rect -22107 1408 -15892 1472
rect -15828 1408 -15808 1472
rect -22107 1392 -15808 1408
rect -22107 1328 -15892 1392
rect -15828 1328 -15808 1392
rect -22107 1312 -15808 1328
rect -22107 1248 -15892 1312
rect -15828 1248 -15808 1312
rect -22107 1232 -15808 1248
rect -22107 1168 -15892 1232
rect -15828 1168 -15808 1232
rect -22107 1152 -15808 1168
rect -22107 1088 -15892 1152
rect -15828 1088 -15808 1152
rect -22107 1072 -15808 1088
rect -22107 1008 -15892 1072
rect -15828 1008 -15808 1072
rect -22107 992 -15808 1008
rect -22107 928 -15892 992
rect -15828 928 -15808 992
rect -22107 912 -15808 928
rect -22107 848 -15892 912
rect -15828 848 -15808 912
rect -22107 832 -15808 848
rect -22107 768 -15892 832
rect -15828 768 -15808 832
rect -22107 752 -15808 768
rect -22107 688 -15892 752
rect -15828 688 -15808 752
rect -22107 672 -15808 688
rect -22107 608 -15892 672
rect -15828 608 -15808 672
rect -22107 592 -15808 608
rect -22107 528 -15892 592
rect -15828 528 -15808 592
rect -22107 512 -15808 528
rect -22107 448 -15892 512
rect -15828 448 -15808 512
rect -22107 432 -15808 448
rect -22107 368 -15892 432
rect -15828 368 -15808 432
rect -22107 352 -15808 368
rect -22107 288 -15892 352
rect -15828 288 -15808 352
rect -22107 272 -15808 288
rect -22107 208 -15892 272
rect -15828 208 -15808 272
rect -22107 192 -15808 208
rect -22107 128 -15892 192
rect -15828 128 -15808 192
rect -22107 112 -15808 128
rect -22107 48 -15892 112
rect -15828 48 -15808 112
rect -22107 32 -15808 48
rect -22107 -32 -15892 32
rect -15828 -32 -15808 32
rect -22107 -48 -15808 -32
rect -22107 -112 -15892 -48
rect -15828 -112 -15808 -48
rect -22107 -128 -15808 -112
rect -22107 -192 -15892 -128
rect -15828 -192 -15808 -128
rect -22107 -208 -15808 -192
rect -22107 -272 -15892 -208
rect -15828 -272 -15808 -208
rect -22107 -288 -15808 -272
rect -22107 -352 -15892 -288
rect -15828 -352 -15808 -288
rect -22107 -368 -15808 -352
rect -22107 -432 -15892 -368
rect -15828 -432 -15808 -368
rect -22107 -448 -15808 -432
rect -22107 -512 -15892 -448
rect -15828 -512 -15808 -448
rect -22107 -528 -15808 -512
rect -22107 -592 -15892 -528
rect -15828 -592 -15808 -528
rect -22107 -608 -15808 -592
rect -22107 -672 -15892 -608
rect -15828 -672 -15808 -608
rect -22107 -688 -15808 -672
rect -22107 -752 -15892 -688
rect -15828 -752 -15808 -688
rect -22107 -768 -15808 -752
rect -22107 -832 -15892 -768
rect -15828 -832 -15808 -768
rect -22107 -848 -15808 -832
rect -22107 -912 -15892 -848
rect -15828 -912 -15808 -848
rect -22107 -928 -15808 -912
rect -22107 -992 -15892 -928
rect -15828 -992 -15808 -928
rect -22107 -1008 -15808 -992
rect -22107 -1072 -15892 -1008
rect -15828 -1072 -15808 -1008
rect -22107 -1088 -15808 -1072
rect -22107 -1152 -15892 -1088
rect -15828 -1152 -15808 -1088
rect -22107 -1168 -15808 -1152
rect -22107 -1232 -15892 -1168
rect -15828 -1232 -15808 -1168
rect -22107 -1248 -15808 -1232
rect -22107 -1312 -15892 -1248
rect -15828 -1312 -15808 -1248
rect -22107 -1328 -15808 -1312
rect -22107 -1392 -15892 -1328
rect -15828 -1392 -15808 -1328
rect -22107 -1408 -15808 -1392
rect -22107 -1472 -15892 -1408
rect -15828 -1472 -15808 -1408
rect -22107 -1488 -15808 -1472
rect -22107 -1552 -15892 -1488
rect -15828 -1552 -15808 -1488
rect -22107 -1568 -15808 -1552
rect -22107 -1632 -15892 -1568
rect -15828 -1632 -15808 -1568
rect -22107 -1648 -15808 -1632
rect -22107 -1712 -15892 -1648
rect -15828 -1712 -15808 -1648
rect -22107 -1728 -15808 -1712
rect -22107 -1792 -15892 -1728
rect -15828 -1792 -15808 -1728
rect -22107 -1808 -15808 -1792
rect -22107 -1872 -15892 -1808
rect -15828 -1872 -15808 -1808
rect -22107 -1888 -15808 -1872
rect -22107 -1952 -15892 -1888
rect -15828 -1952 -15808 -1888
rect -22107 -1968 -15808 -1952
rect -22107 -2032 -15892 -1968
rect -15828 -2032 -15808 -1968
rect -22107 -2048 -15808 -2032
rect -22107 -2112 -15892 -2048
rect -15828 -2112 -15808 -2048
rect -22107 -2128 -15808 -2112
rect -22107 -2192 -15892 -2128
rect -15828 -2192 -15808 -2128
rect -22107 -2208 -15808 -2192
rect -22107 -2272 -15892 -2208
rect -15828 -2272 -15808 -2208
rect -22107 -2288 -15808 -2272
rect -22107 -2352 -15892 -2288
rect -15828 -2352 -15808 -2288
rect -22107 -2368 -15808 -2352
rect -22107 -2432 -15892 -2368
rect -15828 -2432 -15808 -2368
rect -22107 -2448 -15808 -2432
rect -22107 -2512 -15892 -2448
rect -15828 -2512 -15808 -2448
rect -22107 -2528 -15808 -2512
rect -22107 -2592 -15892 -2528
rect -15828 -2592 -15808 -2528
rect -22107 -2608 -15808 -2592
rect -22107 -2672 -15892 -2608
rect -15828 -2672 -15808 -2608
rect -22107 -2688 -15808 -2672
rect -22107 -2752 -15892 -2688
rect -15828 -2752 -15808 -2688
rect -22107 -2768 -15808 -2752
rect -22107 -2832 -15892 -2768
rect -15828 -2832 -15808 -2768
rect -22107 -2848 -15808 -2832
rect -22107 -2912 -15892 -2848
rect -15828 -2912 -15808 -2848
rect -22107 -2928 -15808 -2912
rect -22107 -2992 -15892 -2928
rect -15828 -2992 -15808 -2928
rect -22107 -3008 -15808 -2992
rect -22107 -3072 -15892 -3008
rect -15828 -3072 -15808 -3008
rect -22107 -3100 -15808 -3072
rect -15788 3072 -9489 3100
rect -15788 3008 -9573 3072
rect -9509 3008 -9489 3072
rect -15788 2992 -9489 3008
rect -15788 2928 -9573 2992
rect -9509 2928 -9489 2992
rect -15788 2912 -9489 2928
rect -15788 2848 -9573 2912
rect -9509 2848 -9489 2912
rect -15788 2832 -9489 2848
rect -15788 2768 -9573 2832
rect -9509 2768 -9489 2832
rect -15788 2752 -9489 2768
rect -15788 2688 -9573 2752
rect -9509 2688 -9489 2752
rect -15788 2672 -9489 2688
rect -15788 2608 -9573 2672
rect -9509 2608 -9489 2672
rect -15788 2592 -9489 2608
rect -15788 2528 -9573 2592
rect -9509 2528 -9489 2592
rect -15788 2512 -9489 2528
rect -15788 2448 -9573 2512
rect -9509 2448 -9489 2512
rect -15788 2432 -9489 2448
rect -15788 2368 -9573 2432
rect -9509 2368 -9489 2432
rect -15788 2352 -9489 2368
rect -15788 2288 -9573 2352
rect -9509 2288 -9489 2352
rect -15788 2272 -9489 2288
rect -15788 2208 -9573 2272
rect -9509 2208 -9489 2272
rect -15788 2192 -9489 2208
rect -15788 2128 -9573 2192
rect -9509 2128 -9489 2192
rect -15788 2112 -9489 2128
rect -15788 2048 -9573 2112
rect -9509 2048 -9489 2112
rect -15788 2032 -9489 2048
rect -15788 1968 -9573 2032
rect -9509 1968 -9489 2032
rect -15788 1952 -9489 1968
rect -15788 1888 -9573 1952
rect -9509 1888 -9489 1952
rect -15788 1872 -9489 1888
rect -15788 1808 -9573 1872
rect -9509 1808 -9489 1872
rect -15788 1792 -9489 1808
rect -15788 1728 -9573 1792
rect -9509 1728 -9489 1792
rect -15788 1712 -9489 1728
rect -15788 1648 -9573 1712
rect -9509 1648 -9489 1712
rect -15788 1632 -9489 1648
rect -15788 1568 -9573 1632
rect -9509 1568 -9489 1632
rect -15788 1552 -9489 1568
rect -15788 1488 -9573 1552
rect -9509 1488 -9489 1552
rect -15788 1472 -9489 1488
rect -15788 1408 -9573 1472
rect -9509 1408 -9489 1472
rect -15788 1392 -9489 1408
rect -15788 1328 -9573 1392
rect -9509 1328 -9489 1392
rect -15788 1312 -9489 1328
rect -15788 1248 -9573 1312
rect -9509 1248 -9489 1312
rect -15788 1232 -9489 1248
rect -15788 1168 -9573 1232
rect -9509 1168 -9489 1232
rect -15788 1152 -9489 1168
rect -15788 1088 -9573 1152
rect -9509 1088 -9489 1152
rect -15788 1072 -9489 1088
rect -15788 1008 -9573 1072
rect -9509 1008 -9489 1072
rect -15788 992 -9489 1008
rect -15788 928 -9573 992
rect -9509 928 -9489 992
rect -15788 912 -9489 928
rect -15788 848 -9573 912
rect -9509 848 -9489 912
rect -15788 832 -9489 848
rect -15788 768 -9573 832
rect -9509 768 -9489 832
rect -15788 752 -9489 768
rect -15788 688 -9573 752
rect -9509 688 -9489 752
rect -15788 672 -9489 688
rect -15788 608 -9573 672
rect -9509 608 -9489 672
rect -15788 592 -9489 608
rect -15788 528 -9573 592
rect -9509 528 -9489 592
rect -15788 512 -9489 528
rect -15788 448 -9573 512
rect -9509 448 -9489 512
rect -15788 432 -9489 448
rect -15788 368 -9573 432
rect -9509 368 -9489 432
rect -15788 352 -9489 368
rect -15788 288 -9573 352
rect -9509 288 -9489 352
rect -15788 272 -9489 288
rect -15788 208 -9573 272
rect -9509 208 -9489 272
rect -15788 192 -9489 208
rect -15788 128 -9573 192
rect -9509 128 -9489 192
rect -15788 112 -9489 128
rect -15788 48 -9573 112
rect -9509 48 -9489 112
rect -15788 32 -9489 48
rect -15788 -32 -9573 32
rect -9509 -32 -9489 32
rect -15788 -48 -9489 -32
rect -15788 -112 -9573 -48
rect -9509 -112 -9489 -48
rect -15788 -128 -9489 -112
rect -15788 -192 -9573 -128
rect -9509 -192 -9489 -128
rect -15788 -208 -9489 -192
rect -15788 -272 -9573 -208
rect -9509 -272 -9489 -208
rect -15788 -288 -9489 -272
rect -15788 -352 -9573 -288
rect -9509 -352 -9489 -288
rect -15788 -368 -9489 -352
rect -15788 -432 -9573 -368
rect -9509 -432 -9489 -368
rect -15788 -448 -9489 -432
rect -15788 -512 -9573 -448
rect -9509 -512 -9489 -448
rect -15788 -528 -9489 -512
rect -15788 -592 -9573 -528
rect -9509 -592 -9489 -528
rect -15788 -608 -9489 -592
rect -15788 -672 -9573 -608
rect -9509 -672 -9489 -608
rect -15788 -688 -9489 -672
rect -15788 -752 -9573 -688
rect -9509 -752 -9489 -688
rect -15788 -768 -9489 -752
rect -15788 -832 -9573 -768
rect -9509 -832 -9489 -768
rect -15788 -848 -9489 -832
rect -15788 -912 -9573 -848
rect -9509 -912 -9489 -848
rect -15788 -928 -9489 -912
rect -15788 -992 -9573 -928
rect -9509 -992 -9489 -928
rect -15788 -1008 -9489 -992
rect -15788 -1072 -9573 -1008
rect -9509 -1072 -9489 -1008
rect -15788 -1088 -9489 -1072
rect -15788 -1152 -9573 -1088
rect -9509 -1152 -9489 -1088
rect -15788 -1168 -9489 -1152
rect -15788 -1232 -9573 -1168
rect -9509 -1232 -9489 -1168
rect -15788 -1248 -9489 -1232
rect -15788 -1312 -9573 -1248
rect -9509 -1312 -9489 -1248
rect -15788 -1328 -9489 -1312
rect -15788 -1392 -9573 -1328
rect -9509 -1392 -9489 -1328
rect -15788 -1408 -9489 -1392
rect -15788 -1472 -9573 -1408
rect -9509 -1472 -9489 -1408
rect -15788 -1488 -9489 -1472
rect -15788 -1552 -9573 -1488
rect -9509 -1552 -9489 -1488
rect -15788 -1568 -9489 -1552
rect -15788 -1632 -9573 -1568
rect -9509 -1632 -9489 -1568
rect -15788 -1648 -9489 -1632
rect -15788 -1712 -9573 -1648
rect -9509 -1712 -9489 -1648
rect -15788 -1728 -9489 -1712
rect -15788 -1792 -9573 -1728
rect -9509 -1792 -9489 -1728
rect -15788 -1808 -9489 -1792
rect -15788 -1872 -9573 -1808
rect -9509 -1872 -9489 -1808
rect -15788 -1888 -9489 -1872
rect -15788 -1952 -9573 -1888
rect -9509 -1952 -9489 -1888
rect -15788 -1968 -9489 -1952
rect -15788 -2032 -9573 -1968
rect -9509 -2032 -9489 -1968
rect -15788 -2048 -9489 -2032
rect -15788 -2112 -9573 -2048
rect -9509 -2112 -9489 -2048
rect -15788 -2128 -9489 -2112
rect -15788 -2192 -9573 -2128
rect -9509 -2192 -9489 -2128
rect -15788 -2208 -9489 -2192
rect -15788 -2272 -9573 -2208
rect -9509 -2272 -9489 -2208
rect -15788 -2288 -9489 -2272
rect -15788 -2352 -9573 -2288
rect -9509 -2352 -9489 -2288
rect -15788 -2368 -9489 -2352
rect -15788 -2432 -9573 -2368
rect -9509 -2432 -9489 -2368
rect -15788 -2448 -9489 -2432
rect -15788 -2512 -9573 -2448
rect -9509 -2512 -9489 -2448
rect -15788 -2528 -9489 -2512
rect -15788 -2592 -9573 -2528
rect -9509 -2592 -9489 -2528
rect -15788 -2608 -9489 -2592
rect -15788 -2672 -9573 -2608
rect -9509 -2672 -9489 -2608
rect -15788 -2688 -9489 -2672
rect -15788 -2752 -9573 -2688
rect -9509 -2752 -9489 -2688
rect -15788 -2768 -9489 -2752
rect -15788 -2832 -9573 -2768
rect -9509 -2832 -9489 -2768
rect -15788 -2848 -9489 -2832
rect -15788 -2912 -9573 -2848
rect -9509 -2912 -9489 -2848
rect -15788 -2928 -9489 -2912
rect -15788 -2992 -9573 -2928
rect -9509 -2992 -9489 -2928
rect -15788 -3008 -9489 -2992
rect -15788 -3072 -9573 -3008
rect -9509 -3072 -9489 -3008
rect -15788 -3100 -9489 -3072
rect -9469 3072 -3170 3100
rect -9469 3008 -3254 3072
rect -3190 3008 -3170 3072
rect -9469 2992 -3170 3008
rect -9469 2928 -3254 2992
rect -3190 2928 -3170 2992
rect -9469 2912 -3170 2928
rect -9469 2848 -3254 2912
rect -3190 2848 -3170 2912
rect -9469 2832 -3170 2848
rect -9469 2768 -3254 2832
rect -3190 2768 -3170 2832
rect -9469 2752 -3170 2768
rect -9469 2688 -3254 2752
rect -3190 2688 -3170 2752
rect -9469 2672 -3170 2688
rect -9469 2608 -3254 2672
rect -3190 2608 -3170 2672
rect -9469 2592 -3170 2608
rect -9469 2528 -3254 2592
rect -3190 2528 -3170 2592
rect -9469 2512 -3170 2528
rect -9469 2448 -3254 2512
rect -3190 2448 -3170 2512
rect -9469 2432 -3170 2448
rect -9469 2368 -3254 2432
rect -3190 2368 -3170 2432
rect -9469 2352 -3170 2368
rect -9469 2288 -3254 2352
rect -3190 2288 -3170 2352
rect -9469 2272 -3170 2288
rect -9469 2208 -3254 2272
rect -3190 2208 -3170 2272
rect -9469 2192 -3170 2208
rect -9469 2128 -3254 2192
rect -3190 2128 -3170 2192
rect -9469 2112 -3170 2128
rect -9469 2048 -3254 2112
rect -3190 2048 -3170 2112
rect -9469 2032 -3170 2048
rect -9469 1968 -3254 2032
rect -3190 1968 -3170 2032
rect -9469 1952 -3170 1968
rect -9469 1888 -3254 1952
rect -3190 1888 -3170 1952
rect -9469 1872 -3170 1888
rect -9469 1808 -3254 1872
rect -3190 1808 -3170 1872
rect -9469 1792 -3170 1808
rect -9469 1728 -3254 1792
rect -3190 1728 -3170 1792
rect -9469 1712 -3170 1728
rect -9469 1648 -3254 1712
rect -3190 1648 -3170 1712
rect -9469 1632 -3170 1648
rect -9469 1568 -3254 1632
rect -3190 1568 -3170 1632
rect -9469 1552 -3170 1568
rect -9469 1488 -3254 1552
rect -3190 1488 -3170 1552
rect -9469 1472 -3170 1488
rect -9469 1408 -3254 1472
rect -3190 1408 -3170 1472
rect -9469 1392 -3170 1408
rect -9469 1328 -3254 1392
rect -3190 1328 -3170 1392
rect -9469 1312 -3170 1328
rect -9469 1248 -3254 1312
rect -3190 1248 -3170 1312
rect -9469 1232 -3170 1248
rect -9469 1168 -3254 1232
rect -3190 1168 -3170 1232
rect -9469 1152 -3170 1168
rect -9469 1088 -3254 1152
rect -3190 1088 -3170 1152
rect -9469 1072 -3170 1088
rect -9469 1008 -3254 1072
rect -3190 1008 -3170 1072
rect -9469 992 -3170 1008
rect -9469 928 -3254 992
rect -3190 928 -3170 992
rect -9469 912 -3170 928
rect -9469 848 -3254 912
rect -3190 848 -3170 912
rect -9469 832 -3170 848
rect -9469 768 -3254 832
rect -3190 768 -3170 832
rect -9469 752 -3170 768
rect -9469 688 -3254 752
rect -3190 688 -3170 752
rect -9469 672 -3170 688
rect -9469 608 -3254 672
rect -3190 608 -3170 672
rect -9469 592 -3170 608
rect -9469 528 -3254 592
rect -3190 528 -3170 592
rect -9469 512 -3170 528
rect -9469 448 -3254 512
rect -3190 448 -3170 512
rect -9469 432 -3170 448
rect -9469 368 -3254 432
rect -3190 368 -3170 432
rect -9469 352 -3170 368
rect -9469 288 -3254 352
rect -3190 288 -3170 352
rect -9469 272 -3170 288
rect -9469 208 -3254 272
rect -3190 208 -3170 272
rect -9469 192 -3170 208
rect -9469 128 -3254 192
rect -3190 128 -3170 192
rect -9469 112 -3170 128
rect -9469 48 -3254 112
rect -3190 48 -3170 112
rect -9469 32 -3170 48
rect -9469 -32 -3254 32
rect -3190 -32 -3170 32
rect -9469 -48 -3170 -32
rect -9469 -112 -3254 -48
rect -3190 -112 -3170 -48
rect -9469 -128 -3170 -112
rect -9469 -192 -3254 -128
rect -3190 -192 -3170 -128
rect -9469 -208 -3170 -192
rect -9469 -272 -3254 -208
rect -3190 -272 -3170 -208
rect -9469 -288 -3170 -272
rect -9469 -352 -3254 -288
rect -3190 -352 -3170 -288
rect -9469 -368 -3170 -352
rect -9469 -432 -3254 -368
rect -3190 -432 -3170 -368
rect -9469 -448 -3170 -432
rect -9469 -512 -3254 -448
rect -3190 -512 -3170 -448
rect -9469 -528 -3170 -512
rect -9469 -592 -3254 -528
rect -3190 -592 -3170 -528
rect -9469 -608 -3170 -592
rect -9469 -672 -3254 -608
rect -3190 -672 -3170 -608
rect -9469 -688 -3170 -672
rect -9469 -752 -3254 -688
rect -3190 -752 -3170 -688
rect -9469 -768 -3170 -752
rect -9469 -832 -3254 -768
rect -3190 -832 -3170 -768
rect -9469 -848 -3170 -832
rect -9469 -912 -3254 -848
rect -3190 -912 -3170 -848
rect -9469 -928 -3170 -912
rect -9469 -992 -3254 -928
rect -3190 -992 -3170 -928
rect -9469 -1008 -3170 -992
rect -9469 -1072 -3254 -1008
rect -3190 -1072 -3170 -1008
rect -9469 -1088 -3170 -1072
rect -9469 -1152 -3254 -1088
rect -3190 -1152 -3170 -1088
rect -9469 -1168 -3170 -1152
rect -9469 -1232 -3254 -1168
rect -3190 -1232 -3170 -1168
rect -9469 -1248 -3170 -1232
rect -9469 -1312 -3254 -1248
rect -3190 -1312 -3170 -1248
rect -9469 -1328 -3170 -1312
rect -9469 -1392 -3254 -1328
rect -3190 -1392 -3170 -1328
rect -9469 -1408 -3170 -1392
rect -9469 -1472 -3254 -1408
rect -3190 -1472 -3170 -1408
rect -9469 -1488 -3170 -1472
rect -9469 -1552 -3254 -1488
rect -3190 -1552 -3170 -1488
rect -9469 -1568 -3170 -1552
rect -9469 -1632 -3254 -1568
rect -3190 -1632 -3170 -1568
rect -9469 -1648 -3170 -1632
rect -9469 -1712 -3254 -1648
rect -3190 -1712 -3170 -1648
rect -9469 -1728 -3170 -1712
rect -9469 -1792 -3254 -1728
rect -3190 -1792 -3170 -1728
rect -9469 -1808 -3170 -1792
rect -9469 -1872 -3254 -1808
rect -3190 -1872 -3170 -1808
rect -9469 -1888 -3170 -1872
rect -9469 -1952 -3254 -1888
rect -3190 -1952 -3170 -1888
rect -9469 -1968 -3170 -1952
rect -9469 -2032 -3254 -1968
rect -3190 -2032 -3170 -1968
rect -9469 -2048 -3170 -2032
rect -9469 -2112 -3254 -2048
rect -3190 -2112 -3170 -2048
rect -9469 -2128 -3170 -2112
rect -9469 -2192 -3254 -2128
rect -3190 -2192 -3170 -2128
rect -9469 -2208 -3170 -2192
rect -9469 -2272 -3254 -2208
rect -3190 -2272 -3170 -2208
rect -9469 -2288 -3170 -2272
rect -9469 -2352 -3254 -2288
rect -3190 -2352 -3170 -2288
rect -9469 -2368 -3170 -2352
rect -9469 -2432 -3254 -2368
rect -3190 -2432 -3170 -2368
rect -9469 -2448 -3170 -2432
rect -9469 -2512 -3254 -2448
rect -3190 -2512 -3170 -2448
rect -9469 -2528 -3170 -2512
rect -9469 -2592 -3254 -2528
rect -3190 -2592 -3170 -2528
rect -9469 -2608 -3170 -2592
rect -9469 -2672 -3254 -2608
rect -3190 -2672 -3170 -2608
rect -9469 -2688 -3170 -2672
rect -9469 -2752 -3254 -2688
rect -3190 -2752 -3170 -2688
rect -9469 -2768 -3170 -2752
rect -9469 -2832 -3254 -2768
rect -3190 -2832 -3170 -2768
rect -9469 -2848 -3170 -2832
rect -9469 -2912 -3254 -2848
rect -3190 -2912 -3170 -2848
rect -9469 -2928 -3170 -2912
rect -9469 -2992 -3254 -2928
rect -3190 -2992 -3170 -2928
rect -9469 -3008 -3170 -2992
rect -9469 -3072 -3254 -3008
rect -3190 -3072 -3170 -3008
rect -9469 -3100 -3170 -3072
rect -3150 3072 3149 3100
rect -3150 3008 3065 3072
rect 3129 3008 3149 3072
rect -3150 2992 3149 3008
rect -3150 2928 3065 2992
rect 3129 2928 3149 2992
rect -3150 2912 3149 2928
rect -3150 2848 3065 2912
rect 3129 2848 3149 2912
rect -3150 2832 3149 2848
rect -3150 2768 3065 2832
rect 3129 2768 3149 2832
rect -3150 2752 3149 2768
rect -3150 2688 3065 2752
rect 3129 2688 3149 2752
rect -3150 2672 3149 2688
rect -3150 2608 3065 2672
rect 3129 2608 3149 2672
rect -3150 2592 3149 2608
rect -3150 2528 3065 2592
rect 3129 2528 3149 2592
rect -3150 2512 3149 2528
rect -3150 2448 3065 2512
rect 3129 2448 3149 2512
rect -3150 2432 3149 2448
rect -3150 2368 3065 2432
rect 3129 2368 3149 2432
rect -3150 2352 3149 2368
rect -3150 2288 3065 2352
rect 3129 2288 3149 2352
rect -3150 2272 3149 2288
rect -3150 2208 3065 2272
rect 3129 2208 3149 2272
rect -3150 2192 3149 2208
rect -3150 2128 3065 2192
rect 3129 2128 3149 2192
rect -3150 2112 3149 2128
rect -3150 2048 3065 2112
rect 3129 2048 3149 2112
rect -3150 2032 3149 2048
rect -3150 1968 3065 2032
rect 3129 1968 3149 2032
rect -3150 1952 3149 1968
rect -3150 1888 3065 1952
rect 3129 1888 3149 1952
rect -3150 1872 3149 1888
rect -3150 1808 3065 1872
rect 3129 1808 3149 1872
rect -3150 1792 3149 1808
rect -3150 1728 3065 1792
rect 3129 1728 3149 1792
rect -3150 1712 3149 1728
rect -3150 1648 3065 1712
rect 3129 1648 3149 1712
rect -3150 1632 3149 1648
rect -3150 1568 3065 1632
rect 3129 1568 3149 1632
rect -3150 1552 3149 1568
rect -3150 1488 3065 1552
rect 3129 1488 3149 1552
rect -3150 1472 3149 1488
rect -3150 1408 3065 1472
rect 3129 1408 3149 1472
rect -3150 1392 3149 1408
rect -3150 1328 3065 1392
rect 3129 1328 3149 1392
rect -3150 1312 3149 1328
rect -3150 1248 3065 1312
rect 3129 1248 3149 1312
rect -3150 1232 3149 1248
rect -3150 1168 3065 1232
rect 3129 1168 3149 1232
rect -3150 1152 3149 1168
rect -3150 1088 3065 1152
rect 3129 1088 3149 1152
rect -3150 1072 3149 1088
rect -3150 1008 3065 1072
rect 3129 1008 3149 1072
rect -3150 992 3149 1008
rect -3150 928 3065 992
rect 3129 928 3149 992
rect -3150 912 3149 928
rect -3150 848 3065 912
rect 3129 848 3149 912
rect -3150 832 3149 848
rect -3150 768 3065 832
rect 3129 768 3149 832
rect -3150 752 3149 768
rect -3150 688 3065 752
rect 3129 688 3149 752
rect -3150 672 3149 688
rect -3150 608 3065 672
rect 3129 608 3149 672
rect -3150 592 3149 608
rect -3150 528 3065 592
rect 3129 528 3149 592
rect -3150 512 3149 528
rect -3150 448 3065 512
rect 3129 448 3149 512
rect -3150 432 3149 448
rect -3150 368 3065 432
rect 3129 368 3149 432
rect -3150 352 3149 368
rect -3150 288 3065 352
rect 3129 288 3149 352
rect -3150 272 3149 288
rect -3150 208 3065 272
rect 3129 208 3149 272
rect -3150 192 3149 208
rect -3150 128 3065 192
rect 3129 128 3149 192
rect -3150 112 3149 128
rect -3150 48 3065 112
rect 3129 48 3149 112
rect -3150 32 3149 48
rect -3150 -32 3065 32
rect 3129 -32 3149 32
rect -3150 -48 3149 -32
rect -3150 -112 3065 -48
rect 3129 -112 3149 -48
rect -3150 -128 3149 -112
rect -3150 -192 3065 -128
rect 3129 -192 3149 -128
rect -3150 -208 3149 -192
rect -3150 -272 3065 -208
rect 3129 -272 3149 -208
rect -3150 -288 3149 -272
rect -3150 -352 3065 -288
rect 3129 -352 3149 -288
rect -3150 -368 3149 -352
rect -3150 -432 3065 -368
rect 3129 -432 3149 -368
rect -3150 -448 3149 -432
rect -3150 -512 3065 -448
rect 3129 -512 3149 -448
rect -3150 -528 3149 -512
rect -3150 -592 3065 -528
rect 3129 -592 3149 -528
rect -3150 -608 3149 -592
rect -3150 -672 3065 -608
rect 3129 -672 3149 -608
rect -3150 -688 3149 -672
rect -3150 -752 3065 -688
rect 3129 -752 3149 -688
rect -3150 -768 3149 -752
rect -3150 -832 3065 -768
rect 3129 -832 3149 -768
rect -3150 -848 3149 -832
rect -3150 -912 3065 -848
rect 3129 -912 3149 -848
rect -3150 -928 3149 -912
rect -3150 -992 3065 -928
rect 3129 -992 3149 -928
rect -3150 -1008 3149 -992
rect -3150 -1072 3065 -1008
rect 3129 -1072 3149 -1008
rect -3150 -1088 3149 -1072
rect -3150 -1152 3065 -1088
rect 3129 -1152 3149 -1088
rect -3150 -1168 3149 -1152
rect -3150 -1232 3065 -1168
rect 3129 -1232 3149 -1168
rect -3150 -1248 3149 -1232
rect -3150 -1312 3065 -1248
rect 3129 -1312 3149 -1248
rect -3150 -1328 3149 -1312
rect -3150 -1392 3065 -1328
rect 3129 -1392 3149 -1328
rect -3150 -1408 3149 -1392
rect -3150 -1472 3065 -1408
rect 3129 -1472 3149 -1408
rect -3150 -1488 3149 -1472
rect -3150 -1552 3065 -1488
rect 3129 -1552 3149 -1488
rect -3150 -1568 3149 -1552
rect -3150 -1632 3065 -1568
rect 3129 -1632 3149 -1568
rect -3150 -1648 3149 -1632
rect -3150 -1712 3065 -1648
rect 3129 -1712 3149 -1648
rect -3150 -1728 3149 -1712
rect -3150 -1792 3065 -1728
rect 3129 -1792 3149 -1728
rect -3150 -1808 3149 -1792
rect -3150 -1872 3065 -1808
rect 3129 -1872 3149 -1808
rect -3150 -1888 3149 -1872
rect -3150 -1952 3065 -1888
rect 3129 -1952 3149 -1888
rect -3150 -1968 3149 -1952
rect -3150 -2032 3065 -1968
rect 3129 -2032 3149 -1968
rect -3150 -2048 3149 -2032
rect -3150 -2112 3065 -2048
rect 3129 -2112 3149 -2048
rect -3150 -2128 3149 -2112
rect -3150 -2192 3065 -2128
rect 3129 -2192 3149 -2128
rect -3150 -2208 3149 -2192
rect -3150 -2272 3065 -2208
rect 3129 -2272 3149 -2208
rect -3150 -2288 3149 -2272
rect -3150 -2352 3065 -2288
rect 3129 -2352 3149 -2288
rect -3150 -2368 3149 -2352
rect -3150 -2432 3065 -2368
rect 3129 -2432 3149 -2368
rect -3150 -2448 3149 -2432
rect -3150 -2512 3065 -2448
rect 3129 -2512 3149 -2448
rect -3150 -2528 3149 -2512
rect -3150 -2592 3065 -2528
rect 3129 -2592 3149 -2528
rect -3150 -2608 3149 -2592
rect -3150 -2672 3065 -2608
rect 3129 -2672 3149 -2608
rect -3150 -2688 3149 -2672
rect -3150 -2752 3065 -2688
rect 3129 -2752 3149 -2688
rect -3150 -2768 3149 -2752
rect -3150 -2832 3065 -2768
rect 3129 -2832 3149 -2768
rect -3150 -2848 3149 -2832
rect -3150 -2912 3065 -2848
rect 3129 -2912 3149 -2848
rect -3150 -2928 3149 -2912
rect -3150 -2992 3065 -2928
rect 3129 -2992 3149 -2928
rect -3150 -3008 3149 -2992
rect -3150 -3072 3065 -3008
rect 3129 -3072 3149 -3008
rect -3150 -3100 3149 -3072
rect 3169 3072 9468 3100
rect 3169 3008 9384 3072
rect 9448 3008 9468 3072
rect 3169 2992 9468 3008
rect 3169 2928 9384 2992
rect 9448 2928 9468 2992
rect 3169 2912 9468 2928
rect 3169 2848 9384 2912
rect 9448 2848 9468 2912
rect 3169 2832 9468 2848
rect 3169 2768 9384 2832
rect 9448 2768 9468 2832
rect 3169 2752 9468 2768
rect 3169 2688 9384 2752
rect 9448 2688 9468 2752
rect 3169 2672 9468 2688
rect 3169 2608 9384 2672
rect 9448 2608 9468 2672
rect 3169 2592 9468 2608
rect 3169 2528 9384 2592
rect 9448 2528 9468 2592
rect 3169 2512 9468 2528
rect 3169 2448 9384 2512
rect 9448 2448 9468 2512
rect 3169 2432 9468 2448
rect 3169 2368 9384 2432
rect 9448 2368 9468 2432
rect 3169 2352 9468 2368
rect 3169 2288 9384 2352
rect 9448 2288 9468 2352
rect 3169 2272 9468 2288
rect 3169 2208 9384 2272
rect 9448 2208 9468 2272
rect 3169 2192 9468 2208
rect 3169 2128 9384 2192
rect 9448 2128 9468 2192
rect 3169 2112 9468 2128
rect 3169 2048 9384 2112
rect 9448 2048 9468 2112
rect 3169 2032 9468 2048
rect 3169 1968 9384 2032
rect 9448 1968 9468 2032
rect 3169 1952 9468 1968
rect 3169 1888 9384 1952
rect 9448 1888 9468 1952
rect 3169 1872 9468 1888
rect 3169 1808 9384 1872
rect 9448 1808 9468 1872
rect 3169 1792 9468 1808
rect 3169 1728 9384 1792
rect 9448 1728 9468 1792
rect 3169 1712 9468 1728
rect 3169 1648 9384 1712
rect 9448 1648 9468 1712
rect 3169 1632 9468 1648
rect 3169 1568 9384 1632
rect 9448 1568 9468 1632
rect 3169 1552 9468 1568
rect 3169 1488 9384 1552
rect 9448 1488 9468 1552
rect 3169 1472 9468 1488
rect 3169 1408 9384 1472
rect 9448 1408 9468 1472
rect 3169 1392 9468 1408
rect 3169 1328 9384 1392
rect 9448 1328 9468 1392
rect 3169 1312 9468 1328
rect 3169 1248 9384 1312
rect 9448 1248 9468 1312
rect 3169 1232 9468 1248
rect 3169 1168 9384 1232
rect 9448 1168 9468 1232
rect 3169 1152 9468 1168
rect 3169 1088 9384 1152
rect 9448 1088 9468 1152
rect 3169 1072 9468 1088
rect 3169 1008 9384 1072
rect 9448 1008 9468 1072
rect 3169 992 9468 1008
rect 3169 928 9384 992
rect 9448 928 9468 992
rect 3169 912 9468 928
rect 3169 848 9384 912
rect 9448 848 9468 912
rect 3169 832 9468 848
rect 3169 768 9384 832
rect 9448 768 9468 832
rect 3169 752 9468 768
rect 3169 688 9384 752
rect 9448 688 9468 752
rect 3169 672 9468 688
rect 3169 608 9384 672
rect 9448 608 9468 672
rect 3169 592 9468 608
rect 3169 528 9384 592
rect 9448 528 9468 592
rect 3169 512 9468 528
rect 3169 448 9384 512
rect 9448 448 9468 512
rect 3169 432 9468 448
rect 3169 368 9384 432
rect 9448 368 9468 432
rect 3169 352 9468 368
rect 3169 288 9384 352
rect 9448 288 9468 352
rect 3169 272 9468 288
rect 3169 208 9384 272
rect 9448 208 9468 272
rect 3169 192 9468 208
rect 3169 128 9384 192
rect 9448 128 9468 192
rect 3169 112 9468 128
rect 3169 48 9384 112
rect 9448 48 9468 112
rect 3169 32 9468 48
rect 3169 -32 9384 32
rect 9448 -32 9468 32
rect 3169 -48 9468 -32
rect 3169 -112 9384 -48
rect 9448 -112 9468 -48
rect 3169 -128 9468 -112
rect 3169 -192 9384 -128
rect 9448 -192 9468 -128
rect 3169 -208 9468 -192
rect 3169 -272 9384 -208
rect 9448 -272 9468 -208
rect 3169 -288 9468 -272
rect 3169 -352 9384 -288
rect 9448 -352 9468 -288
rect 3169 -368 9468 -352
rect 3169 -432 9384 -368
rect 9448 -432 9468 -368
rect 3169 -448 9468 -432
rect 3169 -512 9384 -448
rect 9448 -512 9468 -448
rect 3169 -528 9468 -512
rect 3169 -592 9384 -528
rect 9448 -592 9468 -528
rect 3169 -608 9468 -592
rect 3169 -672 9384 -608
rect 9448 -672 9468 -608
rect 3169 -688 9468 -672
rect 3169 -752 9384 -688
rect 9448 -752 9468 -688
rect 3169 -768 9468 -752
rect 3169 -832 9384 -768
rect 9448 -832 9468 -768
rect 3169 -848 9468 -832
rect 3169 -912 9384 -848
rect 9448 -912 9468 -848
rect 3169 -928 9468 -912
rect 3169 -992 9384 -928
rect 9448 -992 9468 -928
rect 3169 -1008 9468 -992
rect 3169 -1072 9384 -1008
rect 9448 -1072 9468 -1008
rect 3169 -1088 9468 -1072
rect 3169 -1152 9384 -1088
rect 9448 -1152 9468 -1088
rect 3169 -1168 9468 -1152
rect 3169 -1232 9384 -1168
rect 9448 -1232 9468 -1168
rect 3169 -1248 9468 -1232
rect 3169 -1312 9384 -1248
rect 9448 -1312 9468 -1248
rect 3169 -1328 9468 -1312
rect 3169 -1392 9384 -1328
rect 9448 -1392 9468 -1328
rect 3169 -1408 9468 -1392
rect 3169 -1472 9384 -1408
rect 9448 -1472 9468 -1408
rect 3169 -1488 9468 -1472
rect 3169 -1552 9384 -1488
rect 9448 -1552 9468 -1488
rect 3169 -1568 9468 -1552
rect 3169 -1632 9384 -1568
rect 9448 -1632 9468 -1568
rect 3169 -1648 9468 -1632
rect 3169 -1712 9384 -1648
rect 9448 -1712 9468 -1648
rect 3169 -1728 9468 -1712
rect 3169 -1792 9384 -1728
rect 9448 -1792 9468 -1728
rect 3169 -1808 9468 -1792
rect 3169 -1872 9384 -1808
rect 9448 -1872 9468 -1808
rect 3169 -1888 9468 -1872
rect 3169 -1952 9384 -1888
rect 9448 -1952 9468 -1888
rect 3169 -1968 9468 -1952
rect 3169 -2032 9384 -1968
rect 9448 -2032 9468 -1968
rect 3169 -2048 9468 -2032
rect 3169 -2112 9384 -2048
rect 9448 -2112 9468 -2048
rect 3169 -2128 9468 -2112
rect 3169 -2192 9384 -2128
rect 9448 -2192 9468 -2128
rect 3169 -2208 9468 -2192
rect 3169 -2272 9384 -2208
rect 9448 -2272 9468 -2208
rect 3169 -2288 9468 -2272
rect 3169 -2352 9384 -2288
rect 9448 -2352 9468 -2288
rect 3169 -2368 9468 -2352
rect 3169 -2432 9384 -2368
rect 9448 -2432 9468 -2368
rect 3169 -2448 9468 -2432
rect 3169 -2512 9384 -2448
rect 9448 -2512 9468 -2448
rect 3169 -2528 9468 -2512
rect 3169 -2592 9384 -2528
rect 9448 -2592 9468 -2528
rect 3169 -2608 9468 -2592
rect 3169 -2672 9384 -2608
rect 9448 -2672 9468 -2608
rect 3169 -2688 9468 -2672
rect 3169 -2752 9384 -2688
rect 9448 -2752 9468 -2688
rect 3169 -2768 9468 -2752
rect 3169 -2832 9384 -2768
rect 9448 -2832 9468 -2768
rect 3169 -2848 9468 -2832
rect 3169 -2912 9384 -2848
rect 9448 -2912 9468 -2848
rect 3169 -2928 9468 -2912
rect 3169 -2992 9384 -2928
rect 9448 -2992 9468 -2928
rect 3169 -3008 9468 -2992
rect 3169 -3072 9384 -3008
rect 9448 -3072 9468 -3008
rect 3169 -3100 9468 -3072
rect 9488 3072 15787 3100
rect 9488 3008 15703 3072
rect 15767 3008 15787 3072
rect 9488 2992 15787 3008
rect 9488 2928 15703 2992
rect 15767 2928 15787 2992
rect 9488 2912 15787 2928
rect 9488 2848 15703 2912
rect 15767 2848 15787 2912
rect 9488 2832 15787 2848
rect 9488 2768 15703 2832
rect 15767 2768 15787 2832
rect 9488 2752 15787 2768
rect 9488 2688 15703 2752
rect 15767 2688 15787 2752
rect 9488 2672 15787 2688
rect 9488 2608 15703 2672
rect 15767 2608 15787 2672
rect 9488 2592 15787 2608
rect 9488 2528 15703 2592
rect 15767 2528 15787 2592
rect 9488 2512 15787 2528
rect 9488 2448 15703 2512
rect 15767 2448 15787 2512
rect 9488 2432 15787 2448
rect 9488 2368 15703 2432
rect 15767 2368 15787 2432
rect 9488 2352 15787 2368
rect 9488 2288 15703 2352
rect 15767 2288 15787 2352
rect 9488 2272 15787 2288
rect 9488 2208 15703 2272
rect 15767 2208 15787 2272
rect 9488 2192 15787 2208
rect 9488 2128 15703 2192
rect 15767 2128 15787 2192
rect 9488 2112 15787 2128
rect 9488 2048 15703 2112
rect 15767 2048 15787 2112
rect 9488 2032 15787 2048
rect 9488 1968 15703 2032
rect 15767 1968 15787 2032
rect 9488 1952 15787 1968
rect 9488 1888 15703 1952
rect 15767 1888 15787 1952
rect 9488 1872 15787 1888
rect 9488 1808 15703 1872
rect 15767 1808 15787 1872
rect 9488 1792 15787 1808
rect 9488 1728 15703 1792
rect 15767 1728 15787 1792
rect 9488 1712 15787 1728
rect 9488 1648 15703 1712
rect 15767 1648 15787 1712
rect 9488 1632 15787 1648
rect 9488 1568 15703 1632
rect 15767 1568 15787 1632
rect 9488 1552 15787 1568
rect 9488 1488 15703 1552
rect 15767 1488 15787 1552
rect 9488 1472 15787 1488
rect 9488 1408 15703 1472
rect 15767 1408 15787 1472
rect 9488 1392 15787 1408
rect 9488 1328 15703 1392
rect 15767 1328 15787 1392
rect 9488 1312 15787 1328
rect 9488 1248 15703 1312
rect 15767 1248 15787 1312
rect 9488 1232 15787 1248
rect 9488 1168 15703 1232
rect 15767 1168 15787 1232
rect 9488 1152 15787 1168
rect 9488 1088 15703 1152
rect 15767 1088 15787 1152
rect 9488 1072 15787 1088
rect 9488 1008 15703 1072
rect 15767 1008 15787 1072
rect 9488 992 15787 1008
rect 9488 928 15703 992
rect 15767 928 15787 992
rect 9488 912 15787 928
rect 9488 848 15703 912
rect 15767 848 15787 912
rect 9488 832 15787 848
rect 9488 768 15703 832
rect 15767 768 15787 832
rect 9488 752 15787 768
rect 9488 688 15703 752
rect 15767 688 15787 752
rect 9488 672 15787 688
rect 9488 608 15703 672
rect 15767 608 15787 672
rect 9488 592 15787 608
rect 9488 528 15703 592
rect 15767 528 15787 592
rect 9488 512 15787 528
rect 9488 448 15703 512
rect 15767 448 15787 512
rect 9488 432 15787 448
rect 9488 368 15703 432
rect 15767 368 15787 432
rect 9488 352 15787 368
rect 9488 288 15703 352
rect 15767 288 15787 352
rect 9488 272 15787 288
rect 9488 208 15703 272
rect 15767 208 15787 272
rect 9488 192 15787 208
rect 9488 128 15703 192
rect 15767 128 15787 192
rect 9488 112 15787 128
rect 9488 48 15703 112
rect 15767 48 15787 112
rect 9488 32 15787 48
rect 9488 -32 15703 32
rect 15767 -32 15787 32
rect 9488 -48 15787 -32
rect 9488 -112 15703 -48
rect 15767 -112 15787 -48
rect 9488 -128 15787 -112
rect 9488 -192 15703 -128
rect 15767 -192 15787 -128
rect 9488 -208 15787 -192
rect 9488 -272 15703 -208
rect 15767 -272 15787 -208
rect 9488 -288 15787 -272
rect 9488 -352 15703 -288
rect 15767 -352 15787 -288
rect 9488 -368 15787 -352
rect 9488 -432 15703 -368
rect 15767 -432 15787 -368
rect 9488 -448 15787 -432
rect 9488 -512 15703 -448
rect 15767 -512 15787 -448
rect 9488 -528 15787 -512
rect 9488 -592 15703 -528
rect 15767 -592 15787 -528
rect 9488 -608 15787 -592
rect 9488 -672 15703 -608
rect 15767 -672 15787 -608
rect 9488 -688 15787 -672
rect 9488 -752 15703 -688
rect 15767 -752 15787 -688
rect 9488 -768 15787 -752
rect 9488 -832 15703 -768
rect 15767 -832 15787 -768
rect 9488 -848 15787 -832
rect 9488 -912 15703 -848
rect 15767 -912 15787 -848
rect 9488 -928 15787 -912
rect 9488 -992 15703 -928
rect 15767 -992 15787 -928
rect 9488 -1008 15787 -992
rect 9488 -1072 15703 -1008
rect 15767 -1072 15787 -1008
rect 9488 -1088 15787 -1072
rect 9488 -1152 15703 -1088
rect 15767 -1152 15787 -1088
rect 9488 -1168 15787 -1152
rect 9488 -1232 15703 -1168
rect 15767 -1232 15787 -1168
rect 9488 -1248 15787 -1232
rect 9488 -1312 15703 -1248
rect 15767 -1312 15787 -1248
rect 9488 -1328 15787 -1312
rect 9488 -1392 15703 -1328
rect 15767 -1392 15787 -1328
rect 9488 -1408 15787 -1392
rect 9488 -1472 15703 -1408
rect 15767 -1472 15787 -1408
rect 9488 -1488 15787 -1472
rect 9488 -1552 15703 -1488
rect 15767 -1552 15787 -1488
rect 9488 -1568 15787 -1552
rect 9488 -1632 15703 -1568
rect 15767 -1632 15787 -1568
rect 9488 -1648 15787 -1632
rect 9488 -1712 15703 -1648
rect 15767 -1712 15787 -1648
rect 9488 -1728 15787 -1712
rect 9488 -1792 15703 -1728
rect 15767 -1792 15787 -1728
rect 9488 -1808 15787 -1792
rect 9488 -1872 15703 -1808
rect 15767 -1872 15787 -1808
rect 9488 -1888 15787 -1872
rect 9488 -1952 15703 -1888
rect 15767 -1952 15787 -1888
rect 9488 -1968 15787 -1952
rect 9488 -2032 15703 -1968
rect 15767 -2032 15787 -1968
rect 9488 -2048 15787 -2032
rect 9488 -2112 15703 -2048
rect 15767 -2112 15787 -2048
rect 9488 -2128 15787 -2112
rect 9488 -2192 15703 -2128
rect 15767 -2192 15787 -2128
rect 9488 -2208 15787 -2192
rect 9488 -2272 15703 -2208
rect 15767 -2272 15787 -2208
rect 9488 -2288 15787 -2272
rect 9488 -2352 15703 -2288
rect 15767 -2352 15787 -2288
rect 9488 -2368 15787 -2352
rect 9488 -2432 15703 -2368
rect 15767 -2432 15787 -2368
rect 9488 -2448 15787 -2432
rect 9488 -2512 15703 -2448
rect 15767 -2512 15787 -2448
rect 9488 -2528 15787 -2512
rect 9488 -2592 15703 -2528
rect 15767 -2592 15787 -2528
rect 9488 -2608 15787 -2592
rect 9488 -2672 15703 -2608
rect 15767 -2672 15787 -2608
rect 9488 -2688 15787 -2672
rect 9488 -2752 15703 -2688
rect 15767 -2752 15787 -2688
rect 9488 -2768 15787 -2752
rect 9488 -2832 15703 -2768
rect 15767 -2832 15787 -2768
rect 9488 -2848 15787 -2832
rect 9488 -2912 15703 -2848
rect 15767 -2912 15787 -2848
rect 9488 -2928 15787 -2912
rect 9488 -2992 15703 -2928
rect 15767 -2992 15787 -2928
rect 9488 -3008 15787 -2992
rect 9488 -3072 15703 -3008
rect 15767 -3072 15787 -3008
rect 9488 -3100 15787 -3072
rect 15807 3072 22106 3100
rect 15807 3008 22022 3072
rect 22086 3008 22106 3072
rect 15807 2992 22106 3008
rect 15807 2928 22022 2992
rect 22086 2928 22106 2992
rect 15807 2912 22106 2928
rect 15807 2848 22022 2912
rect 22086 2848 22106 2912
rect 15807 2832 22106 2848
rect 15807 2768 22022 2832
rect 22086 2768 22106 2832
rect 15807 2752 22106 2768
rect 15807 2688 22022 2752
rect 22086 2688 22106 2752
rect 15807 2672 22106 2688
rect 15807 2608 22022 2672
rect 22086 2608 22106 2672
rect 15807 2592 22106 2608
rect 15807 2528 22022 2592
rect 22086 2528 22106 2592
rect 15807 2512 22106 2528
rect 15807 2448 22022 2512
rect 22086 2448 22106 2512
rect 15807 2432 22106 2448
rect 15807 2368 22022 2432
rect 22086 2368 22106 2432
rect 15807 2352 22106 2368
rect 15807 2288 22022 2352
rect 22086 2288 22106 2352
rect 15807 2272 22106 2288
rect 15807 2208 22022 2272
rect 22086 2208 22106 2272
rect 15807 2192 22106 2208
rect 15807 2128 22022 2192
rect 22086 2128 22106 2192
rect 15807 2112 22106 2128
rect 15807 2048 22022 2112
rect 22086 2048 22106 2112
rect 15807 2032 22106 2048
rect 15807 1968 22022 2032
rect 22086 1968 22106 2032
rect 15807 1952 22106 1968
rect 15807 1888 22022 1952
rect 22086 1888 22106 1952
rect 15807 1872 22106 1888
rect 15807 1808 22022 1872
rect 22086 1808 22106 1872
rect 15807 1792 22106 1808
rect 15807 1728 22022 1792
rect 22086 1728 22106 1792
rect 15807 1712 22106 1728
rect 15807 1648 22022 1712
rect 22086 1648 22106 1712
rect 15807 1632 22106 1648
rect 15807 1568 22022 1632
rect 22086 1568 22106 1632
rect 15807 1552 22106 1568
rect 15807 1488 22022 1552
rect 22086 1488 22106 1552
rect 15807 1472 22106 1488
rect 15807 1408 22022 1472
rect 22086 1408 22106 1472
rect 15807 1392 22106 1408
rect 15807 1328 22022 1392
rect 22086 1328 22106 1392
rect 15807 1312 22106 1328
rect 15807 1248 22022 1312
rect 22086 1248 22106 1312
rect 15807 1232 22106 1248
rect 15807 1168 22022 1232
rect 22086 1168 22106 1232
rect 15807 1152 22106 1168
rect 15807 1088 22022 1152
rect 22086 1088 22106 1152
rect 15807 1072 22106 1088
rect 15807 1008 22022 1072
rect 22086 1008 22106 1072
rect 15807 992 22106 1008
rect 15807 928 22022 992
rect 22086 928 22106 992
rect 15807 912 22106 928
rect 15807 848 22022 912
rect 22086 848 22106 912
rect 15807 832 22106 848
rect 15807 768 22022 832
rect 22086 768 22106 832
rect 15807 752 22106 768
rect 15807 688 22022 752
rect 22086 688 22106 752
rect 15807 672 22106 688
rect 15807 608 22022 672
rect 22086 608 22106 672
rect 15807 592 22106 608
rect 15807 528 22022 592
rect 22086 528 22106 592
rect 15807 512 22106 528
rect 15807 448 22022 512
rect 22086 448 22106 512
rect 15807 432 22106 448
rect 15807 368 22022 432
rect 22086 368 22106 432
rect 15807 352 22106 368
rect 15807 288 22022 352
rect 22086 288 22106 352
rect 15807 272 22106 288
rect 15807 208 22022 272
rect 22086 208 22106 272
rect 15807 192 22106 208
rect 15807 128 22022 192
rect 22086 128 22106 192
rect 15807 112 22106 128
rect 15807 48 22022 112
rect 22086 48 22106 112
rect 15807 32 22106 48
rect 15807 -32 22022 32
rect 22086 -32 22106 32
rect 15807 -48 22106 -32
rect 15807 -112 22022 -48
rect 22086 -112 22106 -48
rect 15807 -128 22106 -112
rect 15807 -192 22022 -128
rect 22086 -192 22106 -128
rect 15807 -208 22106 -192
rect 15807 -272 22022 -208
rect 22086 -272 22106 -208
rect 15807 -288 22106 -272
rect 15807 -352 22022 -288
rect 22086 -352 22106 -288
rect 15807 -368 22106 -352
rect 15807 -432 22022 -368
rect 22086 -432 22106 -368
rect 15807 -448 22106 -432
rect 15807 -512 22022 -448
rect 22086 -512 22106 -448
rect 15807 -528 22106 -512
rect 15807 -592 22022 -528
rect 22086 -592 22106 -528
rect 15807 -608 22106 -592
rect 15807 -672 22022 -608
rect 22086 -672 22106 -608
rect 15807 -688 22106 -672
rect 15807 -752 22022 -688
rect 22086 -752 22106 -688
rect 15807 -768 22106 -752
rect 15807 -832 22022 -768
rect 22086 -832 22106 -768
rect 15807 -848 22106 -832
rect 15807 -912 22022 -848
rect 22086 -912 22106 -848
rect 15807 -928 22106 -912
rect 15807 -992 22022 -928
rect 22086 -992 22106 -928
rect 15807 -1008 22106 -992
rect 15807 -1072 22022 -1008
rect 22086 -1072 22106 -1008
rect 15807 -1088 22106 -1072
rect 15807 -1152 22022 -1088
rect 22086 -1152 22106 -1088
rect 15807 -1168 22106 -1152
rect 15807 -1232 22022 -1168
rect 22086 -1232 22106 -1168
rect 15807 -1248 22106 -1232
rect 15807 -1312 22022 -1248
rect 22086 -1312 22106 -1248
rect 15807 -1328 22106 -1312
rect 15807 -1392 22022 -1328
rect 22086 -1392 22106 -1328
rect 15807 -1408 22106 -1392
rect 15807 -1472 22022 -1408
rect 22086 -1472 22106 -1408
rect 15807 -1488 22106 -1472
rect 15807 -1552 22022 -1488
rect 22086 -1552 22106 -1488
rect 15807 -1568 22106 -1552
rect 15807 -1632 22022 -1568
rect 22086 -1632 22106 -1568
rect 15807 -1648 22106 -1632
rect 15807 -1712 22022 -1648
rect 22086 -1712 22106 -1648
rect 15807 -1728 22106 -1712
rect 15807 -1792 22022 -1728
rect 22086 -1792 22106 -1728
rect 15807 -1808 22106 -1792
rect 15807 -1872 22022 -1808
rect 22086 -1872 22106 -1808
rect 15807 -1888 22106 -1872
rect 15807 -1952 22022 -1888
rect 22086 -1952 22106 -1888
rect 15807 -1968 22106 -1952
rect 15807 -2032 22022 -1968
rect 22086 -2032 22106 -1968
rect 15807 -2048 22106 -2032
rect 15807 -2112 22022 -2048
rect 22086 -2112 22106 -2048
rect 15807 -2128 22106 -2112
rect 15807 -2192 22022 -2128
rect 22086 -2192 22106 -2128
rect 15807 -2208 22106 -2192
rect 15807 -2272 22022 -2208
rect 22086 -2272 22106 -2208
rect 15807 -2288 22106 -2272
rect 15807 -2352 22022 -2288
rect 22086 -2352 22106 -2288
rect 15807 -2368 22106 -2352
rect 15807 -2432 22022 -2368
rect 22086 -2432 22106 -2368
rect 15807 -2448 22106 -2432
rect 15807 -2512 22022 -2448
rect 22086 -2512 22106 -2448
rect 15807 -2528 22106 -2512
rect 15807 -2592 22022 -2528
rect 22086 -2592 22106 -2528
rect 15807 -2608 22106 -2592
rect 15807 -2672 22022 -2608
rect 22086 -2672 22106 -2608
rect 15807 -2688 22106 -2672
rect 15807 -2752 22022 -2688
rect 22086 -2752 22106 -2688
rect 15807 -2768 22106 -2752
rect 15807 -2832 22022 -2768
rect 22086 -2832 22106 -2768
rect 15807 -2848 22106 -2832
rect 15807 -2912 22022 -2848
rect 22086 -2912 22106 -2848
rect 15807 -2928 22106 -2912
rect 15807 -2992 22022 -2928
rect 22086 -2992 22106 -2928
rect 15807 -3008 22106 -2992
rect 15807 -3072 22022 -3008
rect 22086 -3072 22106 -3008
rect 15807 -3100 22106 -3072
rect 22126 3072 28425 3100
rect 22126 3008 28341 3072
rect 28405 3008 28425 3072
rect 22126 2992 28425 3008
rect 22126 2928 28341 2992
rect 28405 2928 28425 2992
rect 22126 2912 28425 2928
rect 22126 2848 28341 2912
rect 28405 2848 28425 2912
rect 22126 2832 28425 2848
rect 22126 2768 28341 2832
rect 28405 2768 28425 2832
rect 22126 2752 28425 2768
rect 22126 2688 28341 2752
rect 28405 2688 28425 2752
rect 22126 2672 28425 2688
rect 22126 2608 28341 2672
rect 28405 2608 28425 2672
rect 22126 2592 28425 2608
rect 22126 2528 28341 2592
rect 28405 2528 28425 2592
rect 22126 2512 28425 2528
rect 22126 2448 28341 2512
rect 28405 2448 28425 2512
rect 22126 2432 28425 2448
rect 22126 2368 28341 2432
rect 28405 2368 28425 2432
rect 22126 2352 28425 2368
rect 22126 2288 28341 2352
rect 28405 2288 28425 2352
rect 22126 2272 28425 2288
rect 22126 2208 28341 2272
rect 28405 2208 28425 2272
rect 22126 2192 28425 2208
rect 22126 2128 28341 2192
rect 28405 2128 28425 2192
rect 22126 2112 28425 2128
rect 22126 2048 28341 2112
rect 28405 2048 28425 2112
rect 22126 2032 28425 2048
rect 22126 1968 28341 2032
rect 28405 1968 28425 2032
rect 22126 1952 28425 1968
rect 22126 1888 28341 1952
rect 28405 1888 28425 1952
rect 22126 1872 28425 1888
rect 22126 1808 28341 1872
rect 28405 1808 28425 1872
rect 22126 1792 28425 1808
rect 22126 1728 28341 1792
rect 28405 1728 28425 1792
rect 22126 1712 28425 1728
rect 22126 1648 28341 1712
rect 28405 1648 28425 1712
rect 22126 1632 28425 1648
rect 22126 1568 28341 1632
rect 28405 1568 28425 1632
rect 22126 1552 28425 1568
rect 22126 1488 28341 1552
rect 28405 1488 28425 1552
rect 22126 1472 28425 1488
rect 22126 1408 28341 1472
rect 28405 1408 28425 1472
rect 22126 1392 28425 1408
rect 22126 1328 28341 1392
rect 28405 1328 28425 1392
rect 22126 1312 28425 1328
rect 22126 1248 28341 1312
rect 28405 1248 28425 1312
rect 22126 1232 28425 1248
rect 22126 1168 28341 1232
rect 28405 1168 28425 1232
rect 22126 1152 28425 1168
rect 22126 1088 28341 1152
rect 28405 1088 28425 1152
rect 22126 1072 28425 1088
rect 22126 1008 28341 1072
rect 28405 1008 28425 1072
rect 22126 992 28425 1008
rect 22126 928 28341 992
rect 28405 928 28425 992
rect 22126 912 28425 928
rect 22126 848 28341 912
rect 28405 848 28425 912
rect 22126 832 28425 848
rect 22126 768 28341 832
rect 28405 768 28425 832
rect 22126 752 28425 768
rect 22126 688 28341 752
rect 28405 688 28425 752
rect 22126 672 28425 688
rect 22126 608 28341 672
rect 28405 608 28425 672
rect 22126 592 28425 608
rect 22126 528 28341 592
rect 28405 528 28425 592
rect 22126 512 28425 528
rect 22126 448 28341 512
rect 28405 448 28425 512
rect 22126 432 28425 448
rect 22126 368 28341 432
rect 28405 368 28425 432
rect 22126 352 28425 368
rect 22126 288 28341 352
rect 28405 288 28425 352
rect 22126 272 28425 288
rect 22126 208 28341 272
rect 28405 208 28425 272
rect 22126 192 28425 208
rect 22126 128 28341 192
rect 28405 128 28425 192
rect 22126 112 28425 128
rect 22126 48 28341 112
rect 28405 48 28425 112
rect 22126 32 28425 48
rect 22126 -32 28341 32
rect 28405 -32 28425 32
rect 22126 -48 28425 -32
rect 22126 -112 28341 -48
rect 28405 -112 28425 -48
rect 22126 -128 28425 -112
rect 22126 -192 28341 -128
rect 28405 -192 28425 -128
rect 22126 -208 28425 -192
rect 22126 -272 28341 -208
rect 28405 -272 28425 -208
rect 22126 -288 28425 -272
rect 22126 -352 28341 -288
rect 28405 -352 28425 -288
rect 22126 -368 28425 -352
rect 22126 -432 28341 -368
rect 28405 -432 28425 -368
rect 22126 -448 28425 -432
rect 22126 -512 28341 -448
rect 28405 -512 28425 -448
rect 22126 -528 28425 -512
rect 22126 -592 28341 -528
rect 28405 -592 28425 -528
rect 22126 -608 28425 -592
rect 22126 -672 28341 -608
rect 28405 -672 28425 -608
rect 22126 -688 28425 -672
rect 22126 -752 28341 -688
rect 28405 -752 28425 -688
rect 22126 -768 28425 -752
rect 22126 -832 28341 -768
rect 28405 -832 28425 -768
rect 22126 -848 28425 -832
rect 22126 -912 28341 -848
rect 28405 -912 28425 -848
rect 22126 -928 28425 -912
rect 22126 -992 28341 -928
rect 28405 -992 28425 -928
rect 22126 -1008 28425 -992
rect 22126 -1072 28341 -1008
rect 28405 -1072 28425 -1008
rect 22126 -1088 28425 -1072
rect 22126 -1152 28341 -1088
rect 28405 -1152 28425 -1088
rect 22126 -1168 28425 -1152
rect 22126 -1232 28341 -1168
rect 28405 -1232 28425 -1168
rect 22126 -1248 28425 -1232
rect 22126 -1312 28341 -1248
rect 28405 -1312 28425 -1248
rect 22126 -1328 28425 -1312
rect 22126 -1392 28341 -1328
rect 28405 -1392 28425 -1328
rect 22126 -1408 28425 -1392
rect 22126 -1472 28341 -1408
rect 28405 -1472 28425 -1408
rect 22126 -1488 28425 -1472
rect 22126 -1552 28341 -1488
rect 28405 -1552 28425 -1488
rect 22126 -1568 28425 -1552
rect 22126 -1632 28341 -1568
rect 28405 -1632 28425 -1568
rect 22126 -1648 28425 -1632
rect 22126 -1712 28341 -1648
rect 28405 -1712 28425 -1648
rect 22126 -1728 28425 -1712
rect 22126 -1792 28341 -1728
rect 28405 -1792 28425 -1728
rect 22126 -1808 28425 -1792
rect 22126 -1872 28341 -1808
rect 28405 -1872 28425 -1808
rect 22126 -1888 28425 -1872
rect 22126 -1952 28341 -1888
rect 28405 -1952 28425 -1888
rect 22126 -1968 28425 -1952
rect 22126 -2032 28341 -1968
rect 28405 -2032 28425 -1968
rect 22126 -2048 28425 -2032
rect 22126 -2112 28341 -2048
rect 28405 -2112 28425 -2048
rect 22126 -2128 28425 -2112
rect 22126 -2192 28341 -2128
rect 28405 -2192 28425 -2128
rect 22126 -2208 28425 -2192
rect 22126 -2272 28341 -2208
rect 28405 -2272 28425 -2208
rect 22126 -2288 28425 -2272
rect 22126 -2352 28341 -2288
rect 28405 -2352 28425 -2288
rect 22126 -2368 28425 -2352
rect 22126 -2432 28341 -2368
rect 28405 -2432 28425 -2368
rect 22126 -2448 28425 -2432
rect 22126 -2512 28341 -2448
rect 28405 -2512 28425 -2448
rect 22126 -2528 28425 -2512
rect 22126 -2592 28341 -2528
rect 28405 -2592 28425 -2528
rect 22126 -2608 28425 -2592
rect 22126 -2672 28341 -2608
rect 28405 -2672 28425 -2608
rect 22126 -2688 28425 -2672
rect 22126 -2752 28341 -2688
rect 28405 -2752 28425 -2688
rect 22126 -2768 28425 -2752
rect 22126 -2832 28341 -2768
rect 28405 -2832 28425 -2768
rect 22126 -2848 28425 -2832
rect 22126 -2912 28341 -2848
rect 28405 -2912 28425 -2848
rect 22126 -2928 28425 -2912
rect 22126 -2992 28341 -2928
rect 28405 -2992 28425 -2928
rect 22126 -3008 28425 -2992
rect 22126 -3072 28341 -3008
rect 28405 -3072 28425 -3008
rect 22126 -3100 28425 -3072
rect 28445 3072 34744 3100
rect 28445 3008 34660 3072
rect 34724 3008 34744 3072
rect 28445 2992 34744 3008
rect 28445 2928 34660 2992
rect 34724 2928 34744 2992
rect 28445 2912 34744 2928
rect 28445 2848 34660 2912
rect 34724 2848 34744 2912
rect 28445 2832 34744 2848
rect 28445 2768 34660 2832
rect 34724 2768 34744 2832
rect 28445 2752 34744 2768
rect 28445 2688 34660 2752
rect 34724 2688 34744 2752
rect 28445 2672 34744 2688
rect 28445 2608 34660 2672
rect 34724 2608 34744 2672
rect 28445 2592 34744 2608
rect 28445 2528 34660 2592
rect 34724 2528 34744 2592
rect 28445 2512 34744 2528
rect 28445 2448 34660 2512
rect 34724 2448 34744 2512
rect 28445 2432 34744 2448
rect 28445 2368 34660 2432
rect 34724 2368 34744 2432
rect 28445 2352 34744 2368
rect 28445 2288 34660 2352
rect 34724 2288 34744 2352
rect 28445 2272 34744 2288
rect 28445 2208 34660 2272
rect 34724 2208 34744 2272
rect 28445 2192 34744 2208
rect 28445 2128 34660 2192
rect 34724 2128 34744 2192
rect 28445 2112 34744 2128
rect 28445 2048 34660 2112
rect 34724 2048 34744 2112
rect 28445 2032 34744 2048
rect 28445 1968 34660 2032
rect 34724 1968 34744 2032
rect 28445 1952 34744 1968
rect 28445 1888 34660 1952
rect 34724 1888 34744 1952
rect 28445 1872 34744 1888
rect 28445 1808 34660 1872
rect 34724 1808 34744 1872
rect 28445 1792 34744 1808
rect 28445 1728 34660 1792
rect 34724 1728 34744 1792
rect 28445 1712 34744 1728
rect 28445 1648 34660 1712
rect 34724 1648 34744 1712
rect 28445 1632 34744 1648
rect 28445 1568 34660 1632
rect 34724 1568 34744 1632
rect 28445 1552 34744 1568
rect 28445 1488 34660 1552
rect 34724 1488 34744 1552
rect 28445 1472 34744 1488
rect 28445 1408 34660 1472
rect 34724 1408 34744 1472
rect 28445 1392 34744 1408
rect 28445 1328 34660 1392
rect 34724 1328 34744 1392
rect 28445 1312 34744 1328
rect 28445 1248 34660 1312
rect 34724 1248 34744 1312
rect 28445 1232 34744 1248
rect 28445 1168 34660 1232
rect 34724 1168 34744 1232
rect 28445 1152 34744 1168
rect 28445 1088 34660 1152
rect 34724 1088 34744 1152
rect 28445 1072 34744 1088
rect 28445 1008 34660 1072
rect 34724 1008 34744 1072
rect 28445 992 34744 1008
rect 28445 928 34660 992
rect 34724 928 34744 992
rect 28445 912 34744 928
rect 28445 848 34660 912
rect 34724 848 34744 912
rect 28445 832 34744 848
rect 28445 768 34660 832
rect 34724 768 34744 832
rect 28445 752 34744 768
rect 28445 688 34660 752
rect 34724 688 34744 752
rect 28445 672 34744 688
rect 28445 608 34660 672
rect 34724 608 34744 672
rect 28445 592 34744 608
rect 28445 528 34660 592
rect 34724 528 34744 592
rect 28445 512 34744 528
rect 28445 448 34660 512
rect 34724 448 34744 512
rect 28445 432 34744 448
rect 28445 368 34660 432
rect 34724 368 34744 432
rect 28445 352 34744 368
rect 28445 288 34660 352
rect 34724 288 34744 352
rect 28445 272 34744 288
rect 28445 208 34660 272
rect 34724 208 34744 272
rect 28445 192 34744 208
rect 28445 128 34660 192
rect 34724 128 34744 192
rect 28445 112 34744 128
rect 28445 48 34660 112
rect 34724 48 34744 112
rect 28445 32 34744 48
rect 28445 -32 34660 32
rect 34724 -32 34744 32
rect 28445 -48 34744 -32
rect 28445 -112 34660 -48
rect 34724 -112 34744 -48
rect 28445 -128 34744 -112
rect 28445 -192 34660 -128
rect 34724 -192 34744 -128
rect 28445 -208 34744 -192
rect 28445 -272 34660 -208
rect 34724 -272 34744 -208
rect 28445 -288 34744 -272
rect 28445 -352 34660 -288
rect 34724 -352 34744 -288
rect 28445 -368 34744 -352
rect 28445 -432 34660 -368
rect 34724 -432 34744 -368
rect 28445 -448 34744 -432
rect 28445 -512 34660 -448
rect 34724 -512 34744 -448
rect 28445 -528 34744 -512
rect 28445 -592 34660 -528
rect 34724 -592 34744 -528
rect 28445 -608 34744 -592
rect 28445 -672 34660 -608
rect 34724 -672 34744 -608
rect 28445 -688 34744 -672
rect 28445 -752 34660 -688
rect 34724 -752 34744 -688
rect 28445 -768 34744 -752
rect 28445 -832 34660 -768
rect 34724 -832 34744 -768
rect 28445 -848 34744 -832
rect 28445 -912 34660 -848
rect 34724 -912 34744 -848
rect 28445 -928 34744 -912
rect 28445 -992 34660 -928
rect 34724 -992 34744 -928
rect 28445 -1008 34744 -992
rect 28445 -1072 34660 -1008
rect 34724 -1072 34744 -1008
rect 28445 -1088 34744 -1072
rect 28445 -1152 34660 -1088
rect 34724 -1152 34744 -1088
rect 28445 -1168 34744 -1152
rect 28445 -1232 34660 -1168
rect 34724 -1232 34744 -1168
rect 28445 -1248 34744 -1232
rect 28445 -1312 34660 -1248
rect 34724 -1312 34744 -1248
rect 28445 -1328 34744 -1312
rect 28445 -1392 34660 -1328
rect 34724 -1392 34744 -1328
rect 28445 -1408 34744 -1392
rect 28445 -1472 34660 -1408
rect 34724 -1472 34744 -1408
rect 28445 -1488 34744 -1472
rect 28445 -1552 34660 -1488
rect 34724 -1552 34744 -1488
rect 28445 -1568 34744 -1552
rect 28445 -1632 34660 -1568
rect 34724 -1632 34744 -1568
rect 28445 -1648 34744 -1632
rect 28445 -1712 34660 -1648
rect 34724 -1712 34744 -1648
rect 28445 -1728 34744 -1712
rect 28445 -1792 34660 -1728
rect 34724 -1792 34744 -1728
rect 28445 -1808 34744 -1792
rect 28445 -1872 34660 -1808
rect 34724 -1872 34744 -1808
rect 28445 -1888 34744 -1872
rect 28445 -1952 34660 -1888
rect 34724 -1952 34744 -1888
rect 28445 -1968 34744 -1952
rect 28445 -2032 34660 -1968
rect 34724 -2032 34744 -1968
rect 28445 -2048 34744 -2032
rect 28445 -2112 34660 -2048
rect 34724 -2112 34744 -2048
rect 28445 -2128 34744 -2112
rect 28445 -2192 34660 -2128
rect 34724 -2192 34744 -2128
rect 28445 -2208 34744 -2192
rect 28445 -2272 34660 -2208
rect 34724 -2272 34744 -2208
rect 28445 -2288 34744 -2272
rect 28445 -2352 34660 -2288
rect 34724 -2352 34744 -2288
rect 28445 -2368 34744 -2352
rect 28445 -2432 34660 -2368
rect 34724 -2432 34744 -2368
rect 28445 -2448 34744 -2432
rect 28445 -2512 34660 -2448
rect 34724 -2512 34744 -2448
rect 28445 -2528 34744 -2512
rect 28445 -2592 34660 -2528
rect 34724 -2592 34744 -2528
rect 28445 -2608 34744 -2592
rect 28445 -2672 34660 -2608
rect 34724 -2672 34744 -2608
rect 28445 -2688 34744 -2672
rect 28445 -2752 34660 -2688
rect 34724 -2752 34744 -2688
rect 28445 -2768 34744 -2752
rect 28445 -2832 34660 -2768
rect 34724 -2832 34744 -2768
rect 28445 -2848 34744 -2832
rect 28445 -2912 34660 -2848
rect 34724 -2912 34744 -2848
rect 28445 -2928 34744 -2912
rect 28445 -2992 34660 -2928
rect 34724 -2992 34744 -2928
rect 28445 -3008 34744 -2992
rect 28445 -3072 34660 -3008
rect 34724 -3072 34744 -3008
rect 28445 -3100 34744 -3072
rect 34764 3072 41063 3100
rect 34764 3008 40979 3072
rect 41043 3008 41063 3072
rect 34764 2992 41063 3008
rect 34764 2928 40979 2992
rect 41043 2928 41063 2992
rect 34764 2912 41063 2928
rect 34764 2848 40979 2912
rect 41043 2848 41063 2912
rect 34764 2832 41063 2848
rect 34764 2768 40979 2832
rect 41043 2768 41063 2832
rect 34764 2752 41063 2768
rect 34764 2688 40979 2752
rect 41043 2688 41063 2752
rect 34764 2672 41063 2688
rect 34764 2608 40979 2672
rect 41043 2608 41063 2672
rect 34764 2592 41063 2608
rect 34764 2528 40979 2592
rect 41043 2528 41063 2592
rect 34764 2512 41063 2528
rect 34764 2448 40979 2512
rect 41043 2448 41063 2512
rect 34764 2432 41063 2448
rect 34764 2368 40979 2432
rect 41043 2368 41063 2432
rect 34764 2352 41063 2368
rect 34764 2288 40979 2352
rect 41043 2288 41063 2352
rect 34764 2272 41063 2288
rect 34764 2208 40979 2272
rect 41043 2208 41063 2272
rect 34764 2192 41063 2208
rect 34764 2128 40979 2192
rect 41043 2128 41063 2192
rect 34764 2112 41063 2128
rect 34764 2048 40979 2112
rect 41043 2048 41063 2112
rect 34764 2032 41063 2048
rect 34764 1968 40979 2032
rect 41043 1968 41063 2032
rect 34764 1952 41063 1968
rect 34764 1888 40979 1952
rect 41043 1888 41063 1952
rect 34764 1872 41063 1888
rect 34764 1808 40979 1872
rect 41043 1808 41063 1872
rect 34764 1792 41063 1808
rect 34764 1728 40979 1792
rect 41043 1728 41063 1792
rect 34764 1712 41063 1728
rect 34764 1648 40979 1712
rect 41043 1648 41063 1712
rect 34764 1632 41063 1648
rect 34764 1568 40979 1632
rect 41043 1568 41063 1632
rect 34764 1552 41063 1568
rect 34764 1488 40979 1552
rect 41043 1488 41063 1552
rect 34764 1472 41063 1488
rect 34764 1408 40979 1472
rect 41043 1408 41063 1472
rect 34764 1392 41063 1408
rect 34764 1328 40979 1392
rect 41043 1328 41063 1392
rect 34764 1312 41063 1328
rect 34764 1248 40979 1312
rect 41043 1248 41063 1312
rect 34764 1232 41063 1248
rect 34764 1168 40979 1232
rect 41043 1168 41063 1232
rect 34764 1152 41063 1168
rect 34764 1088 40979 1152
rect 41043 1088 41063 1152
rect 34764 1072 41063 1088
rect 34764 1008 40979 1072
rect 41043 1008 41063 1072
rect 34764 992 41063 1008
rect 34764 928 40979 992
rect 41043 928 41063 992
rect 34764 912 41063 928
rect 34764 848 40979 912
rect 41043 848 41063 912
rect 34764 832 41063 848
rect 34764 768 40979 832
rect 41043 768 41063 832
rect 34764 752 41063 768
rect 34764 688 40979 752
rect 41043 688 41063 752
rect 34764 672 41063 688
rect 34764 608 40979 672
rect 41043 608 41063 672
rect 34764 592 41063 608
rect 34764 528 40979 592
rect 41043 528 41063 592
rect 34764 512 41063 528
rect 34764 448 40979 512
rect 41043 448 41063 512
rect 34764 432 41063 448
rect 34764 368 40979 432
rect 41043 368 41063 432
rect 34764 352 41063 368
rect 34764 288 40979 352
rect 41043 288 41063 352
rect 34764 272 41063 288
rect 34764 208 40979 272
rect 41043 208 41063 272
rect 34764 192 41063 208
rect 34764 128 40979 192
rect 41043 128 41063 192
rect 34764 112 41063 128
rect 34764 48 40979 112
rect 41043 48 41063 112
rect 34764 32 41063 48
rect 34764 -32 40979 32
rect 41043 -32 41063 32
rect 34764 -48 41063 -32
rect 34764 -112 40979 -48
rect 41043 -112 41063 -48
rect 34764 -128 41063 -112
rect 34764 -192 40979 -128
rect 41043 -192 41063 -128
rect 34764 -208 41063 -192
rect 34764 -272 40979 -208
rect 41043 -272 41063 -208
rect 34764 -288 41063 -272
rect 34764 -352 40979 -288
rect 41043 -352 41063 -288
rect 34764 -368 41063 -352
rect 34764 -432 40979 -368
rect 41043 -432 41063 -368
rect 34764 -448 41063 -432
rect 34764 -512 40979 -448
rect 41043 -512 41063 -448
rect 34764 -528 41063 -512
rect 34764 -592 40979 -528
rect 41043 -592 41063 -528
rect 34764 -608 41063 -592
rect 34764 -672 40979 -608
rect 41043 -672 41063 -608
rect 34764 -688 41063 -672
rect 34764 -752 40979 -688
rect 41043 -752 41063 -688
rect 34764 -768 41063 -752
rect 34764 -832 40979 -768
rect 41043 -832 41063 -768
rect 34764 -848 41063 -832
rect 34764 -912 40979 -848
rect 41043 -912 41063 -848
rect 34764 -928 41063 -912
rect 34764 -992 40979 -928
rect 41043 -992 41063 -928
rect 34764 -1008 41063 -992
rect 34764 -1072 40979 -1008
rect 41043 -1072 41063 -1008
rect 34764 -1088 41063 -1072
rect 34764 -1152 40979 -1088
rect 41043 -1152 41063 -1088
rect 34764 -1168 41063 -1152
rect 34764 -1232 40979 -1168
rect 41043 -1232 41063 -1168
rect 34764 -1248 41063 -1232
rect 34764 -1312 40979 -1248
rect 41043 -1312 41063 -1248
rect 34764 -1328 41063 -1312
rect 34764 -1392 40979 -1328
rect 41043 -1392 41063 -1328
rect 34764 -1408 41063 -1392
rect 34764 -1472 40979 -1408
rect 41043 -1472 41063 -1408
rect 34764 -1488 41063 -1472
rect 34764 -1552 40979 -1488
rect 41043 -1552 41063 -1488
rect 34764 -1568 41063 -1552
rect 34764 -1632 40979 -1568
rect 41043 -1632 41063 -1568
rect 34764 -1648 41063 -1632
rect 34764 -1712 40979 -1648
rect 41043 -1712 41063 -1648
rect 34764 -1728 41063 -1712
rect 34764 -1792 40979 -1728
rect 41043 -1792 41063 -1728
rect 34764 -1808 41063 -1792
rect 34764 -1872 40979 -1808
rect 41043 -1872 41063 -1808
rect 34764 -1888 41063 -1872
rect 34764 -1952 40979 -1888
rect 41043 -1952 41063 -1888
rect 34764 -1968 41063 -1952
rect 34764 -2032 40979 -1968
rect 41043 -2032 41063 -1968
rect 34764 -2048 41063 -2032
rect 34764 -2112 40979 -2048
rect 41043 -2112 41063 -2048
rect 34764 -2128 41063 -2112
rect 34764 -2192 40979 -2128
rect 41043 -2192 41063 -2128
rect 34764 -2208 41063 -2192
rect 34764 -2272 40979 -2208
rect 41043 -2272 41063 -2208
rect 34764 -2288 41063 -2272
rect 34764 -2352 40979 -2288
rect 41043 -2352 41063 -2288
rect 34764 -2368 41063 -2352
rect 34764 -2432 40979 -2368
rect 41043 -2432 41063 -2368
rect 34764 -2448 41063 -2432
rect 34764 -2512 40979 -2448
rect 41043 -2512 41063 -2448
rect 34764 -2528 41063 -2512
rect 34764 -2592 40979 -2528
rect 41043 -2592 41063 -2528
rect 34764 -2608 41063 -2592
rect 34764 -2672 40979 -2608
rect 41043 -2672 41063 -2608
rect 34764 -2688 41063 -2672
rect 34764 -2752 40979 -2688
rect 41043 -2752 41063 -2688
rect 34764 -2768 41063 -2752
rect 34764 -2832 40979 -2768
rect 41043 -2832 41063 -2768
rect 34764 -2848 41063 -2832
rect 34764 -2912 40979 -2848
rect 41043 -2912 41063 -2848
rect 34764 -2928 41063 -2912
rect 34764 -2992 40979 -2928
rect 41043 -2992 41063 -2928
rect 34764 -3008 41063 -2992
rect 34764 -3072 40979 -3008
rect 41043 -3072 41063 -3008
rect 34764 -3100 41063 -3072
rect 41083 3072 47382 3100
rect 41083 3008 47298 3072
rect 47362 3008 47382 3072
rect 41083 2992 47382 3008
rect 41083 2928 47298 2992
rect 47362 2928 47382 2992
rect 41083 2912 47382 2928
rect 41083 2848 47298 2912
rect 47362 2848 47382 2912
rect 41083 2832 47382 2848
rect 41083 2768 47298 2832
rect 47362 2768 47382 2832
rect 41083 2752 47382 2768
rect 41083 2688 47298 2752
rect 47362 2688 47382 2752
rect 41083 2672 47382 2688
rect 41083 2608 47298 2672
rect 47362 2608 47382 2672
rect 41083 2592 47382 2608
rect 41083 2528 47298 2592
rect 47362 2528 47382 2592
rect 41083 2512 47382 2528
rect 41083 2448 47298 2512
rect 47362 2448 47382 2512
rect 41083 2432 47382 2448
rect 41083 2368 47298 2432
rect 47362 2368 47382 2432
rect 41083 2352 47382 2368
rect 41083 2288 47298 2352
rect 47362 2288 47382 2352
rect 41083 2272 47382 2288
rect 41083 2208 47298 2272
rect 47362 2208 47382 2272
rect 41083 2192 47382 2208
rect 41083 2128 47298 2192
rect 47362 2128 47382 2192
rect 41083 2112 47382 2128
rect 41083 2048 47298 2112
rect 47362 2048 47382 2112
rect 41083 2032 47382 2048
rect 41083 1968 47298 2032
rect 47362 1968 47382 2032
rect 41083 1952 47382 1968
rect 41083 1888 47298 1952
rect 47362 1888 47382 1952
rect 41083 1872 47382 1888
rect 41083 1808 47298 1872
rect 47362 1808 47382 1872
rect 41083 1792 47382 1808
rect 41083 1728 47298 1792
rect 47362 1728 47382 1792
rect 41083 1712 47382 1728
rect 41083 1648 47298 1712
rect 47362 1648 47382 1712
rect 41083 1632 47382 1648
rect 41083 1568 47298 1632
rect 47362 1568 47382 1632
rect 41083 1552 47382 1568
rect 41083 1488 47298 1552
rect 47362 1488 47382 1552
rect 41083 1472 47382 1488
rect 41083 1408 47298 1472
rect 47362 1408 47382 1472
rect 41083 1392 47382 1408
rect 41083 1328 47298 1392
rect 47362 1328 47382 1392
rect 41083 1312 47382 1328
rect 41083 1248 47298 1312
rect 47362 1248 47382 1312
rect 41083 1232 47382 1248
rect 41083 1168 47298 1232
rect 47362 1168 47382 1232
rect 41083 1152 47382 1168
rect 41083 1088 47298 1152
rect 47362 1088 47382 1152
rect 41083 1072 47382 1088
rect 41083 1008 47298 1072
rect 47362 1008 47382 1072
rect 41083 992 47382 1008
rect 41083 928 47298 992
rect 47362 928 47382 992
rect 41083 912 47382 928
rect 41083 848 47298 912
rect 47362 848 47382 912
rect 41083 832 47382 848
rect 41083 768 47298 832
rect 47362 768 47382 832
rect 41083 752 47382 768
rect 41083 688 47298 752
rect 47362 688 47382 752
rect 41083 672 47382 688
rect 41083 608 47298 672
rect 47362 608 47382 672
rect 41083 592 47382 608
rect 41083 528 47298 592
rect 47362 528 47382 592
rect 41083 512 47382 528
rect 41083 448 47298 512
rect 47362 448 47382 512
rect 41083 432 47382 448
rect 41083 368 47298 432
rect 47362 368 47382 432
rect 41083 352 47382 368
rect 41083 288 47298 352
rect 47362 288 47382 352
rect 41083 272 47382 288
rect 41083 208 47298 272
rect 47362 208 47382 272
rect 41083 192 47382 208
rect 41083 128 47298 192
rect 47362 128 47382 192
rect 41083 112 47382 128
rect 41083 48 47298 112
rect 47362 48 47382 112
rect 41083 32 47382 48
rect 41083 -32 47298 32
rect 47362 -32 47382 32
rect 41083 -48 47382 -32
rect 41083 -112 47298 -48
rect 47362 -112 47382 -48
rect 41083 -128 47382 -112
rect 41083 -192 47298 -128
rect 47362 -192 47382 -128
rect 41083 -208 47382 -192
rect 41083 -272 47298 -208
rect 47362 -272 47382 -208
rect 41083 -288 47382 -272
rect 41083 -352 47298 -288
rect 47362 -352 47382 -288
rect 41083 -368 47382 -352
rect 41083 -432 47298 -368
rect 47362 -432 47382 -368
rect 41083 -448 47382 -432
rect 41083 -512 47298 -448
rect 47362 -512 47382 -448
rect 41083 -528 47382 -512
rect 41083 -592 47298 -528
rect 47362 -592 47382 -528
rect 41083 -608 47382 -592
rect 41083 -672 47298 -608
rect 47362 -672 47382 -608
rect 41083 -688 47382 -672
rect 41083 -752 47298 -688
rect 47362 -752 47382 -688
rect 41083 -768 47382 -752
rect 41083 -832 47298 -768
rect 47362 -832 47382 -768
rect 41083 -848 47382 -832
rect 41083 -912 47298 -848
rect 47362 -912 47382 -848
rect 41083 -928 47382 -912
rect 41083 -992 47298 -928
rect 47362 -992 47382 -928
rect 41083 -1008 47382 -992
rect 41083 -1072 47298 -1008
rect 47362 -1072 47382 -1008
rect 41083 -1088 47382 -1072
rect 41083 -1152 47298 -1088
rect 47362 -1152 47382 -1088
rect 41083 -1168 47382 -1152
rect 41083 -1232 47298 -1168
rect 47362 -1232 47382 -1168
rect 41083 -1248 47382 -1232
rect 41083 -1312 47298 -1248
rect 47362 -1312 47382 -1248
rect 41083 -1328 47382 -1312
rect 41083 -1392 47298 -1328
rect 47362 -1392 47382 -1328
rect 41083 -1408 47382 -1392
rect 41083 -1472 47298 -1408
rect 47362 -1472 47382 -1408
rect 41083 -1488 47382 -1472
rect 41083 -1552 47298 -1488
rect 47362 -1552 47382 -1488
rect 41083 -1568 47382 -1552
rect 41083 -1632 47298 -1568
rect 47362 -1632 47382 -1568
rect 41083 -1648 47382 -1632
rect 41083 -1712 47298 -1648
rect 47362 -1712 47382 -1648
rect 41083 -1728 47382 -1712
rect 41083 -1792 47298 -1728
rect 47362 -1792 47382 -1728
rect 41083 -1808 47382 -1792
rect 41083 -1872 47298 -1808
rect 47362 -1872 47382 -1808
rect 41083 -1888 47382 -1872
rect 41083 -1952 47298 -1888
rect 47362 -1952 47382 -1888
rect 41083 -1968 47382 -1952
rect 41083 -2032 47298 -1968
rect 47362 -2032 47382 -1968
rect 41083 -2048 47382 -2032
rect 41083 -2112 47298 -2048
rect 47362 -2112 47382 -2048
rect 41083 -2128 47382 -2112
rect 41083 -2192 47298 -2128
rect 47362 -2192 47382 -2128
rect 41083 -2208 47382 -2192
rect 41083 -2272 47298 -2208
rect 47362 -2272 47382 -2208
rect 41083 -2288 47382 -2272
rect 41083 -2352 47298 -2288
rect 47362 -2352 47382 -2288
rect 41083 -2368 47382 -2352
rect 41083 -2432 47298 -2368
rect 47362 -2432 47382 -2368
rect 41083 -2448 47382 -2432
rect 41083 -2512 47298 -2448
rect 47362 -2512 47382 -2448
rect 41083 -2528 47382 -2512
rect 41083 -2592 47298 -2528
rect 47362 -2592 47382 -2528
rect 41083 -2608 47382 -2592
rect 41083 -2672 47298 -2608
rect 47362 -2672 47382 -2608
rect 41083 -2688 47382 -2672
rect 41083 -2752 47298 -2688
rect 47362 -2752 47382 -2688
rect 41083 -2768 47382 -2752
rect 41083 -2832 47298 -2768
rect 47362 -2832 47382 -2768
rect 41083 -2848 47382 -2832
rect 41083 -2912 47298 -2848
rect 47362 -2912 47382 -2848
rect 41083 -2928 47382 -2912
rect 41083 -2992 47298 -2928
rect 47362 -2992 47382 -2928
rect 41083 -3008 47382 -2992
rect 41083 -3072 47298 -3008
rect 47362 -3072 47382 -3008
rect 41083 -3100 47382 -3072
rect -47383 -3228 -41084 -3200
rect -47383 -3292 -41168 -3228
rect -41104 -3292 -41084 -3228
rect -47383 -3308 -41084 -3292
rect -47383 -3372 -41168 -3308
rect -41104 -3372 -41084 -3308
rect -47383 -3388 -41084 -3372
rect -47383 -3452 -41168 -3388
rect -41104 -3452 -41084 -3388
rect -47383 -3468 -41084 -3452
rect -47383 -3532 -41168 -3468
rect -41104 -3532 -41084 -3468
rect -47383 -3548 -41084 -3532
rect -47383 -3612 -41168 -3548
rect -41104 -3612 -41084 -3548
rect -47383 -3628 -41084 -3612
rect -47383 -3692 -41168 -3628
rect -41104 -3692 -41084 -3628
rect -47383 -3708 -41084 -3692
rect -47383 -3772 -41168 -3708
rect -41104 -3772 -41084 -3708
rect -47383 -3788 -41084 -3772
rect -47383 -3852 -41168 -3788
rect -41104 -3852 -41084 -3788
rect -47383 -3868 -41084 -3852
rect -47383 -3932 -41168 -3868
rect -41104 -3932 -41084 -3868
rect -47383 -3948 -41084 -3932
rect -47383 -4012 -41168 -3948
rect -41104 -4012 -41084 -3948
rect -47383 -4028 -41084 -4012
rect -47383 -4092 -41168 -4028
rect -41104 -4092 -41084 -4028
rect -47383 -4108 -41084 -4092
rect -47383 -4172 -41168 -4108
rect -41104 -4172 -41084 -4108
rect -47383 -4188 -41084 -4172
rect -47383 -4252 -41168 -4188
rect -41104 -4252 -41084 -4188
rect -47383 -4268 -41084 -4252
rect -47383 -4332 -41168 -4268
rect -41104 -4332 -41084 -4268
rect -47383 -4348 -41084 -4332
rect -47383 -4412 -41168 -4348
rect -41104 -4412 -41084 -4348
rect -47383 -4428 -41084 -4412
rect -47383 -4492 -41168 -4428
rect -41104 -4492 -41084 -4428
rect -47383 -4508 -41084 -4492
rect -47383 -4572 -41168 -4508
rect -41104 -4572 -41084 -4508
rect -47383 -4588 -41084 -4572
rect -47383 -4652 -41168 -4588
rect -41104 -4652 -41084 -4588
rect -47383 -4668 -41084 -4652
rect -47383 -4732 -41168 -4668
rect -41104 -4732 -41084 -4668
rect -47383 -4748 -41084 -4732
rect -47383 -4812 -41168 -4748
rect -41104 -4812 -41084 -4748
rect -47383 -4828 -41084 -4812
rect -47383 -4892 -41168 -4828
rect -41104 -4892 -41084 -4828
rect -47383 -4908 -41084 -4892
rect -47383 -4972 -41168 -4908
rect -41104 -4972 -41084 -4908
rect -47383 -4988 -41084 -4972
rect -47383 -5052 -41168 -4988
rect -41104 -5052 -41084 -4988
rect -47383 -5068 -41084 -5052
rect -47383 -5132 -41168 -5068
rect -41104 -5132 -41084 -5068
rect -47383 -5148 -41084 -5132
rect -47383 -5212 -41168 -5148
rect -41104 -5212 -41084 -5148
rect -47383 -5228 -41084 -5212
rect -47383 -5292 -41168 -5228
rect -41104 -5292 -41084 -5228
rect -47383 -5308 -41084 -5292
rect -47383 -5372 -41168 -5308
rect -41104 -5372 -41084 -5308
rect -47383 -5388 -41084 -5372
rect -47383 -5452 -41168 -5388
rect -41104 -5452 -41084 -5388
rect -47383 -5468 -41084 -5452
rect -47383 -5532 -41168 -5468
rect -41104 -5532 -41084 -5468
rect -47383 -5548 -41084 -5532
rect -47383 -5612 -41168 -5548
rect -41104 -5612 -41084 -5548
rect -47383 -5628 -41084 -5612
rect -47383 -5692 -41168 -5628
rect -41104 -5692 -41084 -5628
rect -47383 -5708 -41084 -5692
rect -47383 -5772 -41168 -5708
rect -41104 -5772 -41084 -5708
rect -47383 -5788 -41084 -5772
rect -47383 -5852 -41168 -5788
rect -41104 -5852 -41084 -5788
rect -47383 -5868 -41084 -5852
rect -47383 -5932 -41168 -5868
rect -41104 -5932 -41084 -5868
rect -47383 -5948 -41084 -5932
rect -47383 -6012 -41168 -5948
rect -41104 -6012 -41084 -5948
rect -47383 -6028 -41084 -6012
rect -47383 -6092 -41168 -6028
rect -41104 -6092 -41084 -6028
rect -47383 -6108 -41084 -6092
rect -47383 -6172 -41168 -6108
rect -41104 -6172 -41084 -6108
rect -47383 -6188 -41084 -6172
rect -47383 -6252 -41168 -6188
rect -41104 -6252 -41084 -6188
rect -47383 -6268 -41084 -6252
rect -47383 -6332 -41168 -6268
rect -41104 -6332 -41084 -6268
rect -47383 -6348 -41084 -6332
rect -47383 -6412 -41168 -6348
rect -41104 -6412 -41084 -6348
rect -47383 -6428 -41084 -6412
rect -47383 -6492 -41168 -6428
rect -41104 -6492 -41084 -6428
rect -47383 -6508 -41084 -6492
rect -47383 -6572 -41168 -6508
rect -41104 -6572 -41084 -6508
rect -47383 -6588 -41084 -6572
rect -47383 -6652 -41168 -6588
rect -41104 -6652 -41084 -6588
rect -47383 -6668 -41084 -6652
rect -47383 -6732 -41168 -6668
rect -41104 -6732 -41084 -6668
rect -47383 -6748 -41084 -6732
rect -47383 -6812 -41168 -6748
rect -41104 -6812 -41084 -6748
rect -47383 -6828 -41084 -6812
rect -47383 -6892 -41168 -6828
rect -41104 -6892 -41084 -6828
rect -47383 -6908 -41084 -6892
rect -47383 -6972 -41168 -6908
rect -41104 -6972 -41084 -6908
rect -47383 -6988 -41084 -6972
rect -47383 -7052 -41168 -6988
rect -41104 -7052 -41084 -6988
rect -47383 -7068 -41084 -7052
rect -47383 -7132 -41168 -7068
rect -41104 -7132 -41084 -7068
rect -47383 -7148 -41084 -7132
rect -47383 -7212 -41168 -7148
rect -41104 -7212 -41084 -7148
rect -47383 -7228 -41084 -7212
rect -47383 -7292 -41168 -7228
rect -41104 -7292 -41084 -7228
rect -47383 -7308 -41084 -7292
rect -47383 -7372 -41168 -7308
rect -41104 -7372 -41084 -7308
rect -47383 -7388 -41084 -7372
rect -47383 -7452 -41168 -7388
rect -41104 -7452 -41084 -7388
rect -47383 -7468 -41084 -7452
rect -47383 -7532 -41168 -7468
rect -41104 -7532 -41084 -7468
rect -47383 -7548 -41084 -7532
rect -47383 -7612 -41168 -7548
rect -41104 -7612 -41084 -7548
rect -47383 -7628 -41084 -7612
rect -47383 -7692 -41168 -7628
rect -41104 -7692 -41084 -7628
rect -47383 -7708 -41084 -7692
rect -47383 -7772 -41168 -7708
rect -41104 -7772 -41084 -7708
rect -47383 -7788 -41084 -7772
rect -47383 -7852 -41168 -7788
rect -41104 -7852 -41084 -7788
rect -47383 -7868 -41084 -7852
rect -47383 -7932 -41168 -7868
rect -41104 -7932 -41084 -7868
rect -47383 -7948 -41084 -7932
rect -47383 -8012 -41168 -7948
rect -41104 -8012 -41084 -7948
rect -47383 -8028 -41084 -8012
rect -47383 -8092 -41168 -8028
rect -41104 -8092 -41084 -8028
rect -47383 -8108 -41084 -8092
rect -47383 -8172 -41168 -8108
rect -41104 -8172 -41084 -8108
rect -47383 -8188 -41084 -8172
rect -47383 -8252 -41168 -8188
rect -41104 -8252 -41084 -8188
rect -47383 -8268 -41084 -8252
rect -47383 -8332 -41168 -8268
rect -41104 -8332 -41084 -8268
rect -47383 -8348 -41084 -8332
rect -47383 -8412 -41168 -8348
rect -41104 -8412 -41084 -8348
rect -47383 -8428 -41084 -8412
rect -47383 -8492 -41168 -8428
rect -41104 -8492 -41084 -8428
rect -47383 -8508 -41084 -8492
rect -47383 -8572 -41168 -8508
rect -41104 -8572 -41084 -8508
rect -47383 -8588 -41084 -8572
rect -47383 -8652 -41168 -8588
rect -41104 -8652 -41084 -8588
rect -47383 -8668 -41084 -8652
rect -47383 -8732 -41168 -8668
rect -41104 -8732 -41084 -8668
rect -47383 -8748 -41084 -8732
rect -47383 -8812 -41168 -8748
rect -41104 -8812 -41084 -8748
rect -47383 -8828 -41084 -8812
rect -47383 -8892 -41168 -8828
rect -41104 -8892 -41084 -8828
rect -47383 -8908 -41084 -8892
rect -47383 -8972 -41168 -8908
rect -41104 -8972 -41084 -8908
rect -47383 -8988 -41084 -8972
rect -47383 -9052 -41168 -8988
rect -41104 -9052 -41084 -8988
rect -47383 -9068 -41084 -9052
rect -47383 -9132 -41168 -9068
rect -41104 -9132 -41084 -9068
rect -47383 -9148 -41084 -9132
rect -47383 -9212 -41168 -9148
rect -41104 -9212 -41084 -9148
rect -47383 -9228 -41084 -9212
rect -47383 -9292 -41168 -9228
rect -41104 -9292 -41084 -9228
rect -47383 -9308 -41084 -9292
rect -47383 -9372 -41168 -9308
rect -41104 -9372 -41084 -9308
rect -47383 -9400 -41084 -9372
rect -41064 -3228 -34765 -3200
rect -41064 -3292 -34849 -3228
rect -34785 -3292 -34765 -3228
rect -41064 -3308 -34765 -3292
rect -41064 -3372 -34849 -3308
rect -34785 -3372 -34765 -3308
rect -41064 -3388 -34765 -3372
rect -41064 -3452 -34849 -3388
rect -34785 -3452 -34765 -3388
rect -41064 -3468 -34765 -3452
rect -41064 -3532 -34849 -3468
rect -34785 -3532 -34765 -3468
rect -41064 -3548 -34765 -3532
rect -41064 -3612 -34849 -3548
rect -34785 -3612 -34765 -3548
rect -41064 -3628 -34765 -3612
rect -41064 -3692 -34849 -3628
rect -34785 -3692 -34765 -3628
rect -41064 -3708 -34765 -3692
rect -41064 -3772 -34849 -3708
rect -34785 -3772 -34765 -3708
rect -41064 -3788 -34765 -3772
rect -41064 -3852 -34849 -3788
rect -34785 -3852 -34765 -3788
rect -41064 -3868 -34765 -3852
rect -41064 -3932 -34849 -3868
rect -34785 -3932 -34765 -3868
rect -41064 -3948 -34765 -3932
rect -41064 -4012 -34849 -3948
rect -34785 -4012 -34765 -3948
rect -41064 -4028 -34765 -4012
rect -41064 -4092 -34849 -4028
rect -34785 -4092 -34765 -4028
rect -41064 -4108 -34765 -4092
rect -41064 -4172 -34849 -4108
rect -34785 -4172 -34765 -4108
rect -41064 -4188 -34765 -4172
rect -41064 -4252 -34849 -4188
rect -34785 -4252 -34765 -4188
rect -41064 -4268 -34765 -4252
rect -41064 -4332 -34849 -4268
rect -34785 -4332 -34765 -4268
rect -41064 -4348 -34765 -4332
rect -41064 -4412 -34849 -4348
rect -34785 -4412 -34765 -4348
rect -41064 -4428 -34765 -4412
rect -41064 -4492 -34849 -4428
rect -34785 -4492 -34765 -4428
rect -41064 -4508 -34765 -4492
rect -41064 -4572 -34849 -4508
rect -34785 -4572 -34765 -4508
rect -41064 -4588 -34765 -4572
rect -41064 -4652 -34849 -4588
rect -34785 -4652 -34765 -4588
rect -41064 -4668 -34765 -4652
rect -41064 -4732 -34849 -4668
rect -34785 -4732 -34765 -4668
rect -41064 -4748 -34765 -4732
rect -41064 -4812 -34849 -4748
rect -34785 -4812 -34765 -4748
rect -41064 -4828 -34765 -4812
rect -41064 -4892 -34849 -4828
rect -34785 -4892 -34765 -4828
rect -41064 -4908 -34765 -4892
rect -41064 -4972 -34849 -4908
rect -34785 -4972 -34765 -4908
rect -41064 -4988 -34765 -4972
rect -41064 -5052 -34849 -4988
rect -34785 -5052 -34765 -4988
rect -41064 -5068 -34765 -5052
rect -41064 -5132 -34849 -5068
rect -34785 -5132 -34765 -5068
rect -41064 -5148 -34765 -5132
rect -41064 -5212 -34849 -5148
rect -34785 -5212 -34765 -5148
rect -41064 -5228 -34765 -5212
rect -41064 -5292 -34849 -5228
rect -34785 -5292 -34765 -5228
rect -41064 -5308 -34765 -5292
rect -41064 -5372 -34849 -5308
rect -34785 -5372 -34765 -5308
rect -41064 -5388 -34765 -5372
rect -41064 -5452 -34849 -5388
rect -34785 -5452 -34765 -5388
rect -41064 -5468 -34765 -5452
rect -41064 -5532 -34849 -5468
rect -34785 -5532 -34765 -5468
rect -41064 -5548 -34765 -5532
rect -41064 -5612 -34849 -5548
rect -34785 -5612 -34765 -5548
rect -41064 -5628 -34765 -5612
rect -41064 -5692 -34849 -5628
rect -34785 -5692 -34765 -5628
rect -41064 -5708 -34765 -5692
rect -41064 -5772 -34849 -5708
rect -34785 -5772 -34765 -5708
rect -41064 -5788 -34765 -5772
rect -41064 -5852 -34849 -5788
rect -34785 -5852 -34765 -5788
rect -41064 -5868 -34765 -5852
rect -41064 -5932 -34849 -5868
rect -34785 -5932 -34765 -5868
rect -41064 -5948 -34765 -5932
rect -41064 -6012 -34849 -5948
rect -34785 -6012 -34765 -5948
rect -41064 -6028 -34765 -6012
rect -41064 -6092 -34849 -6028
rect -34785 -6092 -34765 -6028
rect -41064 -6108 -34765 -6092
rect -41064 -6172 -34849 -6108
rect -34785 -6172 -34765 -6108
rect -41064 -6188 -34765 -6172
rect -41064 -6252 -34849 -6188
rect -34785 -6252 -34765 -6188
rect -41064 -6268 -34765 -6252
rect -41064 -6332 -34849 -6268
rect -34785 -6332 -34765 -6268
rect -41064 -6348 -34765 -6332
rect -41064 -6412 -34849 -6348
rect -34785 -6412 -34765 -6348
rect -41064 -6428 -34765 -6412
rect -41064 -6492 -34849 -6428
rect -34785 -6492 -34765 -6428
rect -41064 -6508 -34765 -6492
rect -41064 -6572 -34849 -6508
rect -34785 -6572 -34765 -6508
rect -41064 -6588 -34765 -6572
rect -41064 -6652 -34849 -6588
rect -34785 -6652 -34765 -6588
rect -41064 -6668 -34765 -6652
rect -41064 -6732 -34849 -6668
rect -34785 -6732 -34765 -6668
rect -41064 -6748 -34765 -6732
rect -41064 -6812 -34849 -6748
rect -34785 -6812 -34765 -6748
rect -41064 -6828 -34765 -6812
rect -41064 -6892 -34849 -6828
rect -34785 -6892 -34765 -6828
rect -41064 -6908 -34765 -6892
rect -41064 -6972 -34849 -6908
rect -34785 -6972 -34765 -6908
rect -41064 -6988 -34765 -6972
rect -41064 -7052 -34849 -6988
rect -34785 -7052 -34765 -6988
rect -41064 -7068 -34765 -7052
rect -41064 -7132 -34849 -7068
rect -34785 -7132 -34765 -7068
rect -41064 -7148 -34765 -7132
rect -41064 -7212 -34849 -7148
rect -34785 -7212 -34765 -7148
rect -41064 -7228 -34765 -7212
rect -41064 -7292 -34849 -7228
rect -34785 -7292 -34765 -7228
rect -41064 -7308 -34765 -7292
rect -41064 -7372 -34849 -7308
rect -34785 -7372 -34765 -7308
rect -41064 -7388 -34765 -7372
rect -41064 -7452 -34849 -7388
rect -34785 -7452 -34765 -7388
rect -41064 -7468 -34765 -7452
rect -41064 -7532 -34849 -7468
rect -34785 -7532 -34765 -7468
rect -41064 -7548 -34765 -7532
rect -41064 -7612 -34849 -7548
rect -34785 -7612 -34765 -7548
rect -41064 -7628 -34765 -7612
rect -41064 -7692 -34849 -7628
rect -34785 -7692 -34765 -7628
rect -41064 -7708 -34765 -7692
rect -41064 -7772 -34849 -7708
rect -34785 -7772 -34765 -7708
rect -41064 -7788 -34765 -7772
rect -41064 -7852 -34849 -7788
rect -34785 -7852 -34765 -7788
rect -41064 -7868 -34765 -7852
rect -41064 -7932 -34849 -7868
rect -34785 -7932 -34765 -7868
rect -41064 -7948 -34765 -7932
rect -41064 -8012 -34849 -7948
rect -34785 -8012 -34765 -7948
rect -41064 -8028 -34765 -8012
rect -41064 -8092 -34849 -8028
rect -34785 -8092 -34765 -8028
rect -41064 -8108 -34765 -8092
rect -41064 -8172 -34849 -8108
rect -34785 -8172 -34765 -8108
rect -41064 -8188 -34765 -8172
rect -41064 -8252 -34849 -8188
rect -34785 -8252 -34765 -8188
rect -41064 -8268 -34765 -8252
rect -41064 -8332 -34849 -8268
rect -34785 -8332 -34765 -8268
rect -41064 -8348 -34765 -8332
rect -41064 -8412 -34849 -8348
rect -34785 -8412 -34765 -8348
rect -41064 -8428 -34765 -8412
rect -41064 -8492 -34849 -8428
rect -34785 -8492 -34765 -8428
rect -41064 -8508 -34765 -8492
rect -41064 -8572 -34849 -8508
rect -34785 -8572 -34765 -8508
rect -41064 -8588 -34765 -8572
rect -41064 -8652 -34849 -8588
rect -34785 -8652 -34765 -8588
rect -41064 -8668 -34765 -8652
rect -41064 -8732 -34849 -8668
rect -34785 -8732 -34765 -8668
rect -41064 -8748 -34765 -8732
rect -41064 -8812 -34849 -8748
rect -34785 -8812 -34765 -8748
rect -41064 -8828 -34765 -8812
rect -41064 -8892 -34849 -8828
rect -34785 -8892 -34765 -8828
rect -41064 -8908 -34765 -8892
rect -41064 -8972 -34849 -8908
rect -34785 -8972 -34765 -8908
rect -41064 -8988 -34765 -8972
rect -41064 -9052 -34849 -8988
rect -34785 -9052 -34765 -8988
rect -41064 -9068 -34765 -9052
rect -41064 -9132 -34849 -9068
rect -34785 -9132 -34765 -9068
rect -41064 -9148 -34765 -9132
rect -41064 -9212 -34849 -9148
rect -34785 -9212 -34765 -9148
rect -41064 -9228 -34765 -9212
rect -41064 -9292 -34849 -9228
rect -34785 -9292 -34765 -9228
rect -41064 -9308 -34765 -9292
rect -41064 -9372 -34849 -9308
rect -34785 -9372 -34765 -9308
rect -41064 -9400 -34765 -9372
rect -34745 -3228 -28446 -3200
rect -34745 -3292 -28530 -3228
rect -28466 -3292 -28446 -3228
rect -34745 -3308 -28446 -3292
rect -34745 -3372 -28530 -3308
rect -28466 -3372 -28446 -3308
rect -34745 -3388 -28446 -3372
rect -34745 -3452 -28530 -3388
rect -28466 -3452 -28446 -3388
rect -34745 -3468 -28446 -3452
rect -34745 -3532 -28530 -3468
rect -28466 -3532 -28446 -3468
rect -34745 -3548 -28446 -3532
rect -34745 -3612 -28530 -3548
rect -28466 -3612 -28446 -3548
rect -34745 -3628 -28446 -3612
rect -34745 -3692 -28530 -3628
rect -28466 -3692 -28446 -3628
rect -34745 -3708 -28446 -3692
rect -34745 -3772 -28530 -3708
rect -28466 -3772 -28446 -3708
rect -34745 -3788 -28446 -3772
rect -34745 -3852 -28530 -3788
rect -28466 -3852 -28446 -3788
rect -34745 -3868 -28446 -3852
rect -34745 -3932 -28530 -3868
rect -28466 -3932 -28446 -3868
rect -34745 -3948 -28446 -3932
rect -34745 -4012 -28530 -3948
rect -28466 -4012 -28446 -3948
rect -34745 -4028 -28446 -4012
rect -34745 -4092 -28530 -4028
rect -28466 -4092 -28446 -4028
rect -34745 -4108 -28446 -4092
rect -34745 -4172 -28530 -4108
rect -28466 -4172 -28446 -4108
rect -34745 -4188 -28446 -4172
rect -34745 -4252 -28530 -4188
rect -28466 -4252 -28446 -4188
rect -34745 -4268 -28446 -4252
rect -34745 -4332 -28530 -4268
rect -28466 -4332 -28446 -4268
rect -34745 -4348 -28446 -4332
rect -34745 -4412 -28530 -4348
rect -28466 -4412 -28446 -4348
rect -34745 -4428 -28446 -4412
rect -34745 -4492 -28530 -4428
rect -28466 -4492 -28446 -4428
rect -34745 -4508 -28446 -4492
rect -34745 -4572 -28530 -4508
rect -28466 -4572 -28446 -4508
rect -34745 -4588 -28446 -4572
rect -34745 -4652 -28530 -4588
rect -28466 -4652 -28446 -4588
rect -34745 -4668 -28446 -4652
rect -34745 -4732 -28530 -4668
rect -28466 -4732 -28446 -4668
rect -34745 -4748 -28446 -4732
rect -34745 -4812 -28530 -4748
rect -28466 -4812 -28446 -4748
rect -34745 -4828 -28446 -4812
rect -34745 -4892 -28530 -4828
rect -28466 -4892 -28446 -4828
rect -34745 -4908 -28446 -4892
rect -34745 -4972 -28530 -4908
rect -28466 -4972 -28446 -4908
rect -34745 -4988 -28446 -4972
rect -34745 -5052 -28530 -4988
rect -28466 -5052 -28446 -4988
rect -34745 -5068 -28446 -5052
rect -34745 -5132 -28530 -5068
rect -28466 -5132 -28446 -5068
rect -34745 -5148 -28446 -5132
rect -34745 -5212 -28530 -5148
rect -28466 -5212 -28446 -5148
rect -34745 -5228 -28446 -5212
rect -34745 -5292 -28530 -5228
rect -28466 -5292 -28446 -5228
rect -34745 -5308 -28446 -5292
rect -34745 -5372 -28530 -5308
rect -28466 -5372 -28446 -5308
rect -34745 -5388 -28446 -5372
rect -34745 -5452 -28530 -5388
rect -28466 -5452 -28446 -5388
rect -34745 -5468 -28446 -5452
rect -34745 -5532 -28530 -5468
rect -28466 -5532 -28446 -5468
rect -34745 -5548 -28446 -5532
rect -34745 -5612 -28530 -5548
rect -28466 -5612 -28446 -5548
rect -34745 -5628 -28446 -5612
rect -34745 -5692 -28530 -5628
rect -28466 -5692 -28446 -5628
rect -34745 -5708 -28446 -5692
rect -34745 -5772 -28530 -5708
rect -28466 -5772 -28446 -5708
rect -34745 -5788 -28446 -5772
rect -34745 -5852 -28530 -5788
rect -28466 -5852 -28446 -5788
rect -34745 -5868 -28446 -5852
rect -34745 -5932 -28530 -5868
rect -28466 -5932 -28446 -5868
rect -34745 -5948 -28446 -5932
rect -34745 -6012 -28530 -5948
rect -28466 -6012 -28446 -5948
rect -34745 -6028 -28446 -6012
rect -34745 -6092 -28530 -6028
rect -28466 -6092 -28446 -6028
rect -34745 -6108 -28446 -6092
rect -34745 -6172 -28530 -6108
rect -28466 -6172 -28446 -6108
rect -34745 -6188 -28446 -6172
rect -34745 -6252 -28530 -6188
rect -28466 -6252 -28446 -6188
rect -34745 -6268 -28446 -6252
rect -34745 -6332 -28530 -6268
rect -28466 -6332 -28446 -6268
rect -34745 -6348 -28446 -6332
rect -34745 -6412 -28530 -6348
rect -28466 -6412 -28446 -6348
rect -34745 -6428 -28446 -6412
rect -34745 -6492 -28530 -6428
rect -28466 -6492 -28446 -6428
rect -34745 -6508 -28446 -6492
rect -34745 -6572 -28530 -6508
rect -28466 -6572 -28446 -6508
rect -34745 -6588 -28446 -6572
rect -34745 -6652 -28530 -6588
rect -28466 -6652 -28446 -6588
rect -34745 -6668 -28446 -6652
rect -34745 -6732 -28530 -6668
rect -28466 -6732 -28446 -6668
rect -34745 -6748 -28446 -6732
rect -34745 -6812 -28530 -6748
rect -28466 -6812 -28446 -6748
rect -34745 -6828 -28446 -6812
rect -34745 -6892 -28530 -6828
rect -28466 -6892 -28446 -6828
rect -34745 -6908 -28446 -6892
rect -34745 -6972 -28530 -6908
rect -28466 -6972 -28446 -6908
rect -34745 -6988 -28446 -6972
rect -34745 -7052 -28530 -6988
rect -28466 -7052 -28446 -6988
rect -34745 -7068 -28446 -7052
rect -34745 -7132 -28530 -7068
rect -28466 -7132 -28446 -7068
rect -34745 -7148 -28446 -7132
rect -34745 -7212 -28530 -7148
rect -28466 -7212 -28446 -7148
rect -34745 -7228 -28446 -7212
rect -34745 -7292 -28530 -7228
rect -28466 -7292 -28446 -7228
rect -34745 -7308 -28446 -7292
rect -34745 -7372 -28530 -7308
rect -28466 -7372 -28446 -7308
rect -34745 -7388 -28446 -7372
rect -34745 -7452 -28530 -7388
rect -28466 -7452 -28446 -7388
rect -34745 -7468 -28446 -7452
rect -34745 -7532 -28530 -7468
rect -28466 -7532 -28446 -7468
rect -34745 -7548 -28446 -7532
rect -34745 -7612 -28530 -7548
rect -28466 -7612 -28446 -7548
rect -34745 -7628 -28446 -7612
rect -34745 -7692 -28530 -7628
rect -28466 -7692 -28446 -7628
rect -34745 -7708 -28446 -7692
rect -34745 -7772 -28530 -7708
rect -28466 -7772 -28446 -7708
rect -34745 -7788 -28446 -7772
rect -34745 -7852 -28530 -7788
rect -28466 -7852 -28446 -7788
rect -34745 -7868 -28446 -7852
rect -34745 -7932 -28530 -7868
rect -28466 -7932 -28446 -7868
rect -34745 -7948 -28446 -7932
rect -34745 -8012 -28530 -7948
rect -28466 -8012 -28446 -7948
rect -34745 -8028 -28446 -8012
rect -34745 -8092 -28530 -8028
rect -28466 -8092 -28446 -8028
rect -34745 -8108 -28446 -8092
rect -34745 -8172 -28530 -8108
rect -28466 -8172 -28446 -8108
rect -34745 -8188 -28446 -8172
rect -34745 -8252 -28530 -8188
rect -28466 -8252 -28446 -8188
rect -34745 -8268 -28446 -8252
rect -34745 -8332 -28530 -8268
rect -28466 -8332 -28446 -8268
rect -34745 -8348 -28446 -8332
rect -34745 -8412 -28530 -8348
rect -28466 -8412 -28446 -8348
rect -34745 -8428 -28446 -8412
rect -34745 -8492 -28530 -8428
rect -28466 -8492 -28446 -8428
rect -34745 -8508 -28446 -8492
rect -34745 -8572 -28530 -8508
rect -28466 -8572 -28446 -8508
rect -34745 -8588 -28446 -8572
rect -34745 -8652 -28530 -8588
rect -28466 -8652 -28446 -8588
rect -34745 -8668 -28446 -8652
rect -34745 -8732 -28530 -8668
rect -28466 -8732 -28446 -8668
rect -34745 -8748 -28446 -8732
rect -34745 -8812 -28530 -8748
rect -28466 -8812 -28446 -8748
rect -34745 -8828 -28446 -8812
rect -34745 -8892 -28530 -8828
rect -28466 -8892 -28446 -8828
rect -34745 -8908 -28446 -8892
rect -34745 -8972 -28530 -8908
rect -28466 -8972 -28446 -8908
rect -34745 -8988 -28446 -8972
rect -34745 -9052 -28530 -8988
rect -28466 -9052 -28446 -8988
rect -34745 -9068 -28446 -9052
rect -34745 -9132 -28530 -9068
rect -28466 -9132 -28446 -9068
rect -34745 -9148 -28446 -9132
rect -34745 -9212 -28530 -9148
rect -28466 -9212 -28446 -9148
rect -34745 -9228 -28446 -9212
rect -34745 -9292 -28530 -9228
rect -28466 -9292 -28446 -9228
rect -34745 -9308 -28446 -9292
rect -34745 -9372 -28530 -9308
rect -28466 -9372 -28446 -9308
rect -34745 -9400 -28446 -9372
rect -28426 -3228 -22127 -3200
rect -28426 -3292 -22211 -3228
rect -22147 -3292 -22127 -3228
rect -28426 -3308 -22127 -3292
rect -28426 -3372 -22211 -3308
rect -22147 -3372 -22127 -3308
rect -28426 -3388 -22127 -3372
rect -28426 -3452 -22211 -3388
rect -22147 -3452 -22127 -3388
rect -28426 -3468 -22127 -3452
rect -28426 -3532 -22211 -3468
rect -22147 -3532 -22127 -3468
rect -28426 -3548 -22127 -3532
rect -28426 -3612 -22211 -3548
rect -22147 -3612 -22127 -3548
rect -28426 -3628 -22127 -3612
rect -28426 -3692 -22211 -3628
rect -22147 -3692 -22127 -3628
rect -28426 -3708 -22127 -3692
rect -28426 -3772 -22211 -3708
rect -22147 -3772 -22127 -3708
rect -28426 -3788 -22127 -3772
rect -28426 -3852 -22211 -3788
rect -22147 -3852 -22127 -3788
rect -28426 -3868 -22127 -3852
rect -28426 -3932 -22211 -3868
rect -22147 -3932 -22127 -3868
rect -28426 -3948 -22127 -3932
rect -28426 -4012 -22211 -3948
rect -22147 -4012 -22127 -3948
rect -28426 -4028 -22127 -4012
rect -28426 -4092 -22211 -4028
rect -22147 -4092 -22127 -4028
rect -28426 -4108 -22127 -4092
rect -28426 -4172 -22211 -4108
rect -22147 -4172 -22127 -4108
rect -28426 -4188 -22127 -4172
rect -28426 -4252 -22211 -4188
rect -22147 -4252 -22127 -4188
rect -28426 -4268 -22127 -4252
rect -28426 -4332 -22211 -4268
rect -22147 -4332 -22127 -4268
rect -28426 -4348 -22127 -4332
rect -28426 -4412 -22211 -4348
rect -22147 -4412 -22127 -4348
rect -28426 -4428 -22127 -4412
rect -28426 -4492 -22211 -4428
rect -22147 -4492 -22127 -4428
rect -28426 -4508 -22127 -4492
rect -28426 -4572 -22211 -4508
rect -22147 -4572 -22127 -4508
rect -28426 -4588 -22127 -4572
rect -28426 -4652 -22211 -4588
rect -22147 -4652 -22127 -4588
rect -28426 -4668 -22127 -4652
rect -28426 -4732 -22211 -4668
rect -22147 -4732 -22127 -4668
rect -28426 -4748 -22127 -4732
rect -28426 -4812 -22211 -4748
rect -22147 -4812 -22127 -4748
rect -28426 -4828 -22127 -4812
rect -28426 -4892 -22211 -4828
rect -22147 -4892 -22127 -4828
rect -28426 -4908 -22127 -4892
rect -28426 -4972 -22211 -4908
rect -22147 -4972 -22127 -4908
rect -28426 -4988 -22127 -4972
rect -28426 -5052 -22211 -4988
rect -22147 -5052 -22127 -4988
rect -28426 -5068 -22127 -5052
rect -28426 -5132 -22211 -5068
rect -22147 -5132 -22127 -5068
rect -28426 -5148 -22127 -5132
rect -28426 -5212 -22211 -5148
rect -22147 -5212 -22127 -5148
rect -28426 -5228 -22127 -5212
rect -28426 -5292 -22211 -5228
rect -22147 -5292 -22127 -5228
rect -28426 -5308 -22127 -5292
rect -28426 -5372 -22211 -5308
rect -22147 -5372 -22127 -5308
rect -28426 -5388 -22127 -5372
rect -28426 -5452 -22211 -5388
rect -22147 -5452 -22127 -5388
rect -28426 -5468 -22127 -5452
rect -28426 -5532 -22211 -5468
rect -22147 -5532 -22127 -5468
rect -28426 -5548 -22127 -5532
rect -28426 -5612 -22211 -5548
rect -22147 -5612 -22127 -5548
rect -28426 -5628 -22127 -5612
rect -28426 -5692 -22211 -5628
rect -22147 -5692 -22127 -5628
rect -28426 -5708 -22127 -5692
rect -28426 -5772 -22211 -5708
rect -22147 -5772 -22127 -5708
rect -28426 -5788 -22127 -5772
rect -28426 -5852 -22211 -5788
rect -22147 -5852 -22127 -5788
rect -28426 -5868 -22127 -5852
rect -28426 -5932 -22211 -5868
rect -22147 -5932 -22127 -5868
rect -28426 -5948 -22127 -5932
rect -28426 -6012 -22211 -5948
rect -22147 -6012 -22127 -5948
rect -28426 -6028 -22127 -6012
rect -28426 -6092 -22211 -6028
rect -22147 -6092 -22127 -6028
rect -28426 -6108 -22127 -6092
rect -28426 -6172 -22211 -6108
rect -22147 -6172 -22127 -6108
rect -28426 -6188 -22127 -6172
rect -28426 -6252 -22211 -6188
rect -22147 -6252 -22127 -6188
rect -28426 -6268 -22127 -6252
rect -28426 -6332 -22211 -6268
rect -22147 -6332 -22127 -6268
rect -28426 -6348 -22127 -6332
rect -28426 -6412 -22211 -6348
rect -22147 -6412 -22127 -6348
rect -28426 -6428 -22127 -6412
rect -28426 -6492 -22211 -6428
rect -22147 -6492 -22127 -6428
rect -28426 -6508 -22127 -6492
rect -28426 -6572 -22211 -6508
rect -22147 -6572 -22127 -6508
rect -28426 -6588 -22127 -6572
rect -28426 -6652 -22211 -6588
rect -22147 -6652 -22127 -6588
rect -28426 -6668 -22127 -6652
rect -28426 -6732 -22211 -6668
rect -22147 -6732 -22127 -6668
rect -28426 -6748 -22127 -6732
rect -28426 -6812 -22211 -6748
rect -22147 -6812 -22127 -6748
rect -28426 -6828 -22127 -6812
rect -28426 -6892 -22211 -6828
rect -22147 -6892 -22127 -6828
rect -28426 -6908 -22127 -6892
rect -28426 -6972 -22211 -6908
rect -22147 -6972 -22127 -6908
rect -28426 -6988 -22127 -6972
rect -28426 -7052 -22211 -6988
rect -22147 -7052 -22127 -6988
rect -28426 -7068 -22127 -7052
rect -28426 -7132 -22211 -7068
rect -22147 -7132 -22127 -7068
rect -28426 -7148 -22127 -7132
rect -28426 -7212 -22211 -7148
rect -22147 -7212 -22127 -7148
rect -28426 -7228 -22127 -7212
rect -28426 -7292 -22211 -7228
rect -22147 -7292 -22127 -7228
rect -28426 -7308 -22127 -7292
rect -28426 -7372 -22211 -7308
rect -22147 -7372 -22127 -7308
rect -28426 -7388 -22127 -7372
rect -28426 -7452 -22211 -7388
rect -22147 -7452 -22127 -7388
rect -28426 -7468 -22127 -7452
rect -28426 -7532 -22211 -7468
rect -22147 -7532 -22127 -7468
rect -28426 -7548 -22127 -7532
rect -28426 -7612 -22211 -7548
rect -22147 -7612 -22127 -7548
rect -28426 -7628 -22127 -7612
rect -28426 -7692 -22211 -7628
rect -22147 -7692 -22127 -7628
rect -28426 -7708 -22127 -7692
rect -28426 -7772 -22211 -7708
rect -22147 -7772 -22127 -7708
rect -28426 -7788 -22127 -7772
rect -28426 -7852 -22211 -7788
rect -22147 -7852 -22127 -7788
rect -28426 -7868 -22127 -7852
rect -28426 -7932 -22211 -7868
rect -22147 -7932 -22127 -7868
rect -28426 -7948 -22127 -7932
rect -28426 -8012 -22211 -7948
rect -22147 -8012 -22127 -7948
rect -28426 -8028 -22127 -8012
rect -28426 -8092 -22211 -8028
rect -22147 -8092 -22127 -8028
rect -28426 -8108 -22127 -8092
rect -28426 -8172 -22211 -8108
rect -22147 -8172 -22127 -8108
rect -28426 -8188 -22127 -8172
rect -28426 -8252 -22211 -8188
rect -22147 -8252 -22127 -8188
rect -28426 -8268 -22127 -8252
rect -28426 -8332 -22211 -8268
rect -22147 -8332 -22127 -8268
rect -28426 -8348 -22127 -8332
rect -28426 -8412 -22211 -8348
rect -22147 -8412 -22127 -8348
rect -28426 -8428 -22127 -8412
rect -28426 -8492 -22211 -8428
rect -22147 -8492 -22127 -8428
rect -28426 -8508 -22127 -8492
rect -28426 -8572 -22211 -8508
rect -22147 -8572 -22127 -8508
rect -28426 -8588 -22127 -8572
rect -28426 -8652 -22211 -8588
rect -22147 -8652 -22127 -8588
rect -28426 -8668 -22127 -8652
rect -28426 -8732 -22211 -8668
rect -22147 -8732 -22127 -8668
rect -28426 -8748 -22127 -8732
rect -28426 -8812 -22211 -8748
rect -22147 -8812 -22127 -8748
rect -28426 -8828 -22127 -8812
rect -28426 -8892 -22211 -8828
rect -22147 -8892 -22127 -8828
rect -28426 -8908 -22127 -8892
rect -28426 -8972 -22211 -8908
rect -22147 -8972 -22127 -8908
rect -28426 -8988 -22127 -8972
rect -28426 -9052 -22211 -8988
rect -22147 -9052 -22127 -8988
rect -28426 -9068 -22127 -9052
rect -28426 -9132 -22211 -9068
rect -22147 -9132 -22127 -9068
rect -28426 -9148 -22127 -9132
rect -28426 -9212 -22211 -9148
rect -22147 -9212 -22127 -9148
rect -28426 -9228 -22127 -9212
rect -28426 -9292 -22211 -9228
rect -22147 -9292 -22127 -9228
rect -28426 -9308 -22127 -9292
rect -28426 -9372 -22211 -9308
rect -22147 -9372 -22127 -9308
rect -28426 -9400 -22127 -9372
rect -22107 -3228 -15808 -3200
rect -22107 -3292 -15892 -3228
rect -15828 -3292 -15808 -3228
rect -22107 -3308 -15808 -3292
rect -22107 -3372 -15892 -3308
rect -15828 -3372 -15808 -3308
rect -22107 -3388 -15808 -3372
rect -22107 -3452 -15892 -3388
rect -15828 -3452 -15808 -3388
rect -22107 -3468 -15808 -3452
rect -22107 -3532 -15892 -3468
rect -15828 -3532 -15808 -3468
rect -22107 -3548 -15808 -3532
rect -22107 -3612 -15892 -3548
rect -15828 -3612 -15808 -3548
rect -22107 -3628 -15808 -3612
rect -22107 -3692 -15892 -3628
rect -15828 -3692 -15808 -3628
rect -22107 -3708 -15808 -3692
rect -22107 -3772 -15892 -3708
rect -15828 -3772 -15808 -3708
rect -22107 -3788 -15808 -3772
rect -22107 -3852 -15892 -3788
rect -15828 -3852 -15808 -3788
rect -22107 -3868 -15808 -3852
rect -22107 -3932 -15892 -3868
rect -15828 -3932 -15808 -3868
rect -22107 -3948 -15808 -3932
rect -22107 -4012 -15892 -3948
rect -15828 -4012 -15808 -3948
rect -22107 -4028 -15808 -4012
rect -22107 -4092 -15892 -4028
rect -15828 -4092 -15808 -4028
rect -22107 -4108 -15808 -4092
rect -22107 -4172 -15892 -4108
rect -15828 -4172 -15808 -4108
rect -22107 -4188 -15808 -4172
rect -22107 -4252 -15892 -4188
rect -15828 -4252 -15808 -4188
rect -22107 -4268 -15808 -4252
rect -22107 -4332 -15892 -4268
rect -15828 -4332 -15808 -4268
rect -22107 -4348 -15808 -4332
rect -22107 -4412 -15892 -4348
rect -15828 -4412 -15808 -4348
rect -22107 -4428 -15808 -4412
rect -22107 -4492 -15892 -4428
rect -15828 -4492 -15808 -4428
rect -22107 -4508 -15808 -4492
rect -22107 -4572 -15892 -4508
rect -15828 -4572 -15808 -4508
rect -22107 -4588 -15808 -4572
rect -22107 -4652 -15892 -4588
rect -15828 -4652 -15808 -4588
rect -22107 -4668 -15808 -4652
rect -22107 -4732 -15892 -4668
rect -15828 -4732 -15808 -4668
rect -22107 -4748 -15808 -4732
rect -22107 -4812 -15892 -4748
rect -15828 -4812 -15808 -4748
rect -22107 -4828 -15808 -4812
rect -22107 -4892 -15892 -4828
rect -15828 -4892 -15808 -4828
rect -22107 -4908 -15808 -4892
rect -22107 -4972 -15892 -4908
rect -15828 -4972 -15808 -4908
rect -22107 -4988 -15808 -4972
rect -22107 -5052 -15892 -4988
rect -15828 -5052 -15808 -4988
rect -22107 -5068 -15808 -5052
rect -22107 -5132 -15892 -5068
rect -15828 -5132 -15808 -5068
rect -22107 -5148 -15808 -5132
rect -22107 -5212 -15892 -5148
rect -15828 -5212 -15808 -5148
rect -22107 -5228 -15808 -5212
rect -22107 -5292 -15892 -5228
rect -15828 -5292 -15808 -5228
rect -22107 -5308 -15808 -5292
rect -22107 -5372 -15892 -5308
rect -15828 -5372 -15808 -5308
rect -22107 -5388 -15808 -5372
rect -22107 -5452 -15892 -5388
rect -15828 -5452 -15808 -5388
rect -22107 -5468 -15808 -5452
rect -22107 -5532 -15892 -5468
rect -15828 -5532 -15808 -5468
rect -22107 -5548 -15808 -5532
rect -22107 -5612 -15892 -5548
rect -15828 -5612 -15808 -5548
rect -22107 -5628 -15808 -5612
rect -22107 -5692 -15892 -5628
rect -15828 -5692 -15808 -5628
rect -22107 -5708 -15808 -5692
rect -22107 -5772 -15892 -5708
rect -15828 -5772 -15808 -5708
rect -22107 -5788 -15808 -5772
rect -22107 -5852 -15892 -5788
rect -15828 -5852 -15808 -5788
rect -22107 -5868 -15808 -5852
rect -22107 -5932 -15892 -5868
rect -15828 -5932 -15808 -5868
rect -22107 -5948 -15808 -5932
rect -22107 -6012 -15892 -5948
rect -15828 -6012 -15808 -5948
rect -22107 -6028 -15808 -6012
rect -22107 -6092 -15892 -6028
rect -15828 -6092 -15808 -6028
rect -22107 -6108 -15808 -6092
rect -22107 -6172 -15892 -6108
rect -15828 -6172 -15808 -6108
rect -22107 -6188 -15808 -6172
rect -22107 -6252 -15892 -6188
rect -15828 -6252 -15808 -6188
rect -22107 -6268 -15808 -6252
rect -22107 -6332 -15892 -6268
rect -15828 -6332 -15808 -6268
rect -22107 -6348 -15808 -6332
rect -22107 -6412 -15892 -6348
rect -15828 -6412 -15808 -6348
rect -22107 -6428 -15808 -6412
rect -22107 -6492 -15892 -6428
rect -15828 -6492 -15808 -6428
rect -22107 -6508 -15808 -6492
rect -22107 -6572 -15892 -6508
rect -15828 -6572 -15808 -6508
rect -22107 -6588 -15808 -6572
rect -22107 -6652 -15892 -6588
rect -15828 -6652 -15808 -6588
rect -22107 -6668 -15808 -6652
rect -22107 -6732 -15892 -6668
rect -15828 -6732 -15808 -6668
rect -22107 -6748 -15808 -6732
rect -22107 -6812 -15892 -6748
rect -15828 -6812 -15808 -6748
rect -22107 -6828 -15808 -6812
rect -22107 -6892 -15892 -6828
rect -15828 -6892 -15808 -6828
rect -22107 -6908 -15808 -6892
rect -22107 -6972 -15892 -6908
rect -15828 -6972 -15808 -6908
rect -22107 -6988 -15808 -6972
rect -22107 -7052 -15892 -6988
rect -15828 -7052 -15808 -6988
rect -22107 -7068 -15808 -7052
rect -22107 -7132 -15892 -7068
rect -15828 -7132 -15808 -7068
rect -22107 -7148 -15808 -7132
rect -22107 -7212 -15892 -7148
rect -15828 -7212 -15808 -7148
rect -22107 -7228 -15808 -7212
rect -22107 -7292 -15892 -7228
rect -15828 -7292 -15808 -7228
rect -22107 -7308 -15808 -7292
rect -22107 -7372 -15892 -7308
rect -15828 -7372 -15808 -7308
rect -22107 -7388 -15808 -7372
rect -22107 -7452 -15892 -7388
rect -15828 -7452 -15808 -7388
rect -22107 -7468 -15808 -7452
rect -22107 -7532 -15892 -7468
rect -15828 -7532 -15808 -7468
rect -22107 -7548 -15808 -7532
rect -22107 -7612 -15892 -7548
rect -15828 -7612 -15808 -7548
rect -22107 -7628 -15808 -7612
rect -22107 -7692 -15892 -7628
rect -15828 -7692 -15808 -7628
rect -22107 -7708 -15808 -7692
rect -22107 -7772 -15892 -7708
rect -15828 -7772 -15808 -7708
rect -22107 -7788 -15808 -7772
rect -22107 -7852 -15892 -7788
rect -15828 -7852 -15808 -7788
rect -22107 -7868 -15808 -7852
rect -22107 -7932 -15892 -7868
rect -15828 -7932 -15808 -7868
rect -22107 -7948 -15808 -7932
rect -22107 -8012 -15892 -7948
rect -15828 -8012 -15808 -7948
rect -22107 -8028 -15808 -8012
rect -22107 -8092 -15892 -8028
rect -15828 -8092 -15808 -8028
rect -22107 -8108 -15808 -8092
rect -22107 -8172 -15892 -8108
rect -15828 -8172 -15808 -8108
rect -22107 -8188 -15808 -8172
rect -22107 -8252 -15892 -8188
rect -15828 -8252 -15808 -8188
rect -22107 -8268 -15808 -8252
rect -22107 -8332 -15892 -8268
rect -15828 -8332 -15808 -8268
rect -22107 -8348 -15808 -8332
rect -22107 -8412 -15892 -8348
rect -15828 -8412 -15808 -8348
rect -22107 -8428 -15808 -8412
rect -22107 -8492 -15892 -8428
rect -15828 -8492 -15808 -8428
rect -22107 -8508 -15808 -8492
rect -22107 -8572 -15892 -8508
rect -15828 -8572 -15808 -8508
rect -22107 -8588 -15808 -8572
rect -22107 -8652 -15892 -8588
rect -15828 -8652 -15808 -8588
rect -22107 -8668 -15808 -8652
rect -22107 -8732 -15892 -8668
rect -15828 -8732 -15808 -8668
rect -22107 -8748 -15808 -8732
rect -22107 -8812 -15892 -8748
rect -15828 -8812 -15808 -8748
rect -22107 -8828 -15808 -8812
rect -22107 -8892 -15892 -8828
rect -15828 -8892 -15808 -8828
rect -22107 -8908 -15808 -8892
rect -22107 -8972 -15892 -8908
rect -15828 -8972 -15808 -8908
rect -22107 -8988 -15808 -8972
rect -22107 -9052 -15892 -8988
rect -15828 -9052 -15808 -8988
rect -22107 -9068 -15808 -9052
rect -22107 -9132 -15892 -9068
rect -15828 -9132 -15808 -9068
rect -22107 -9148 -15808 -9132
rect -22107 -9212 -15892 -9148
rect -15828 -9212 -15808 -9148
rect -22107 -9228 -15808 -9212
rect -22107 -9292 -15892 -9228
rect -15828 -9292 -15808 -9228
rect -22107 -9308 -15808 -9292
rect -22107 -9372 -15892 -9308
rect -15828 -9372 -15808 -9308
rect -22107 -9400 -15808 -9372
rect -15788 -3228 -9489 -3200
rect -15788 -3292 -9573 -3228
rect -9509 -3292 -9489 -3228
rect -15788 -3308 -9489 -3292
rect -15788 -3372 -9573 -3308
rect -9509 -3372 -9489 -3308
rect -15788 -3388 -9489 -3372
rect -15788 -3452 -9573 -3388
rect -9509 -3452 -9489 -3388
rect -15788 -3468 -9489 -3452
rect -15788 -3532 -9573 -3468
rect -9509 -3532 -9489 -3468
rect -15788 -3548 -9489 -3532
rect -15788 -3612 -9573 -3548
rect -9509 -3612 -9489 -3548
rect -15788 -3628 -9489 -3612
rect -15788 -3692 -9573 -3628
rect -9509 -3692 -9489 -3628
rect -15788 -3708 -9489 -3692
rect -15788 -3772 -9573 -3708
rect -9509 -3772 -9489 -3708
rect -15788 -3788 -9489 -3772
rect -15788 -3852 -9573 -3788
rect -9509 -3852 -9489 -3788
rect -15788 -3868 -9489 -3852
rect -15788 -3932 -9573 -3868
rect -9509 -3932 -9489 -3868
rect -15788 -3948 -9489 -3932
rect -15788 -4012 -9573 -3948
rect -9509 -4012 -9489 -3948
rect -15788 -4028 -9489 -4012
rect -15788 -4092 -9573 -4028
rect -9509 -4092 -9489 -4028
rect -15788 -4108 -9489 -4092
rect -15788 -4172 -9573 -4108
rect -9509 -4172 -9489 -4108
rect -15788 -4188 -9489 -4172
rect -15788 -4252 -9573 -4188
rect -9509 -4252 -9489 -4188
rect -15788 -4268 -9489 -4252
rect -15788 -4332 -9573 -4268
rect -9509 -4332 -9489 -4268
rect -15788 -4348 -9489 -4332
rect -15788 -4412 -9573 -4348
rect -9509 -4412 -9489 -4348
rect -15788 -4428 -9489 -4412
rect -15788 -4492 -9573 -4428
rect -9509 -4492 -9489 -4428
rect -15788 -4508 -9489 -4492
rect -15788 -4572 -9573 -4508
rect -9509 -4572 -9489 -4508
rect -15788 -4588 -9489 -4572
rect -15788 -4652 -9573 -4588
rect -9509 -4652 -9489 -4588
rect -15788 -4668 -9489 -4652
rect -15788 -4732 -9573 -4668
rect -9509 -4732 -9489 -4668
rect -15788 -4748 -9489 -4732
rect -15788 -4812 -9573 -4748
rect -9509 -4812 -9489 -4748
rect -15788 -4828 -9489 -4812
rect -15788 -4892 -9573 -4828
rect -9509 -4892 -9489 -4828
rect -15788 -4908 -9489 -4892
rect -15788 -4972 -9573 -4908
rect -9509 -4972 -9489 -4908
rect -15788 -4988 -9489 -4972
rect -15788 -5052 -9573 -4988
rect -9509 -5052 -9489 -4988
rect -15788 -5068 -9489 -5052
rect -15788 -5132 -9573 -5068
rect -9509 -5132 -9489 -5068
rect -15788 -5148 -9489 -5132
rect -15788 -5212 -9573 -5148
rect -9509 -5212 -9489 -5148
rect -15788 -5228 -9489 -5212
rect -15788 -5292 -9573 -5228
rect -9509 -5292 -9489 -5228
rect -15788 -5308 -9489 -5292
rect -15788 -5372 -9573 -5308
rect -9509 -5372 -9489 -5308
rect -15788 -5388 -9489 -5372
rect -15788 -5452 -9573 -5388
rect -9509 -5452 -9489 -5388
rect -15788 -5468 -9489 -5452
rect -15788 -5532 -9573 -5468
rect -9509 -5532 -9489 -5468
rect -15788 -5548 -9489 -5532
rect -15788 -5612 -9573 -5548
rect -9509 -5612 -9489 -5548
rect -15788 -5628 -9489 -5612
rect -15788 -5692 -9573 -5628
rect -9509 -5692 -9489 -5628
rect -15788 -5708 -9489 -5692
rect -15788 -5772 -9573 -5708
rect -9509 -5772 -9489 -5708
rect -15788 -5788 -9489 -5772
rect -15788 -5852 -9573 -5788
rect -9509 -5852 -9489 -5788
rect -15788 -5868 -9489 -5852
rect -15788 -5932 -9573 -5868
rect -9509 -5932 -9489 -5868
rect -15788 -5948 -9489 -5932
rect -15788 -6012 -9573 -5948
rect -9509 -6012 -9489 -5948
rect -15788 -6028 -9489 -6012
rect -15788 -6092 -9573 -6028
rect -9509 -6092 -9489 -6028
rect -15788 -6108 -9489 -6092
rect -15788 -6172 -9573 -6108
rect -9509 -6172 -9489 -6108
rect -15788 -6188 -9489 -6172
rect -15788 -6252 -9573 -6188
rect -9509 -6252 -9489 -6188
rect -15788 -6268 -9489 -6252
rect -15788 -6332 -9573 -6268
rect -9509 -6332 -9489 -6268
rect -15788 -6348 -9489 -6332
rect -15788 -6412 -9573 -6348
rect -9509 -6412 -9489 -6348
rect -15788 -6428 -9489 -6412
rect -15788 -6492 -9573 -6428
rect -9509 -6492 -9489 -6428
rect -15788 -6508 -9489 -6492
rect -15788 -6572 -9573 -6508
rect -9509 -6572 -9489 -6508
rect -15788 -6588 -9489 -6572
rect -15788 -6652 -9573 -6588
rect -9509 -6652 -9489 -6588
rect -15788 -6668 -9489 -6652
rect -15788 -6732 -9573 -6668
rect -9509 -6732 -9489 -6668
rect -15788 -6748 -9489 -6732
rect -15788 -6812 -9573 -6748
rect -9509 -6812 -9489 -6748
rect -15788 -6828 -9489 -6812
rect -15788 -6892 -9573 -6828
rect -9509 -6892 -9489 -6828
rect -15788 -6908 -9489 -6892
rect -15788 -6972 -9573 -6908
rect -9509 -6972 -9489 -6908
rect -15788 -6988 -9489 -6972
rect -15788 -7052 -9573 -6988
rect -9509 -7052 -9489 -6988
rect -15788 -7068 -9489 -7052
rect -15788 -7132 -9573 -7068
rect -9509 -7132 -9489 -7068
rect -15788 -7148 -9489 -7132
rect -15788 -7212 -9573 -7148
rect -9509 -7212 -9489 -7148
rect -15788 -7228 -9489 -7212
rect -15788 -7292 -9573 -7228
rect -9509 -7292 -9489 -7228
rect -15788 -7308 -9489 -7292
rect -15788 -7372 -9573 -7308
rect -9509 -7372 -9489 -7308
rect -15788 -7388 -9489 -7372
rect -15788 -7452 -9573 -7388
rect -9509 -7452 -9489 -7388
rect -15788 -7468 -9489 -7452
rect -15788 -7532 -9573 -7468
rect -9509 -7532 -9489 -7468
rect -15788 -7548 -9489 -7532
rect -15788 -7612 -9573 -7548
rect -9509 -7612 -9489 -7548
rect -15788 -7628 -9489 -7612
rect -15788 -7692 -9573 -7628
rect -9509 -7692 -9489 -7628
rect -15788 -7708 -9489 -7692
rect -15788 -7772 -9573 -7708
rect -9509 -7772 -9489 -7708
rect -15788 -7788 -9489 -7772
rect -15788 -7852 -9573 -7788
rect -9509 -7852 -9489 -7788
rect -15788 -7868 -9489 -7852
rect -15788 -7932 -9573 -7868
rect -9509 -7932 -9489 -7868
rect -15788 -7948 -9489 -7932
rect -15788 -8012 -9573 -7948
rect -9509 -8012 -9489 -7948
rect -15788 -8028 -9489 -8012
rect -15788 -8092 -9573 -8028
rect -9509 -8092 -9489 -8028
rect -15788 -8108 -9489 -8092
rect -15788 -8172 -9573 -8108
rect -9509 -8172 -9489 -8108
rect -15788 -8188 -9489 -8172
rect -15788 -8252 -9573 -8188
rect -9509 -8252 -9489 -8188
rect -15788 -8268 -9489 -8252
rect -15788 -8332 -9573 -8268
rect -9509 -8332 -9489 -8268
rect -15788 -8348 -9489 -8332
rect -15788 -8412 -9573 -8348
rect -9509 -8412 -9489 -8348
rect -15788 -8428 -9489 -8412
rect -15788 -8492 -9573 -8428
rect -9509 -8492 -9489 -8428
rect -15788 -8508 -9489 -8492
rect -15788 -8572 -9573 -8508
rect -9509 -8572 -9489 -8508
rect -15788 -8588 -9489 -8572
rect -15788 -8652 -9573 -8588
rect -9509 -8652 -9489 -8588
rect -15788 -8668 -9489 -8652
rect -15788 -8732 -9573 -8668
rect -9509 -8732 -9489 -8668
rect -15788 -8748 -9489 -8732
rect -15788 -8812 -9573 -8748
rect -9509 -8812 -9489 -8748
rect -15788 -8828 -9489 -8812
rect -15788 -8892 -9573 -8828
rect -9509 -8892 -9489 -8828
rect -15788 -8908 -9489 -8892
rect -15788 -8972 -9573 -8908
rect -9509 -8972 -9489 -8908
rect -15788 -8988 -9489 -8972
rect -15788 -9052 -9573 -8988
rect -9509 -9052 -9489 -8988
rect -15788 -9068 -9489 -9052
rect -15788 -9132 -9573 -9068
rect -9509 -9132 -9489 -9068
rect -15788 -9148 -9489 -9132
rect -15788 -9212 -9573 -9148
rect -9509 -9212 -9489 -9148
rect -15788 -9228 -9489 -9212
rect -15788 -9292 -9573 -9228
rect -9509 -9292 -9489 -9228
rect -15788 -9308 -9489 -9292
rect -15788 -9372 -9573 -9308
rect -9509 -9372 -9489 -9308
rect -15788 -9400 -9489 -9372
rect -9469 -3228 -3170 -3200
rect -9469 -3292 -3254 -3228
rect -3190 -3292 -3170 -3228
rect -9469 -3308 -3170 -3292
rect -9469 -3372 -3254 -3308
rect -3190 -3372 -3170 -3308
rect -9469 -3388 -3170 -3372
rect -9469 -3452 -3254 -3388
rect -3190 -3452 -3170 -3388
rect -9469 -3468 -3170 -3452
rect -9469 -3532 -3254 -3468
rect -3190 -3532 -3170 -3468
rect -9469 -3548 -3170 -3532
rect -9469 -3612 -3254 -3548
rect -3190 -3612 -3170 -3548
rect -9469 -3628 -3170 -3612
rect -9469 -3692 -3254 -3628
rect -3190 -3692 -3170 -3628
rect -9469 -3708 -3170 -3692
rect -9469 -3772 -3254 -3708
rect -3190 -3772 -3170 -3708
rect -9469 -3788 -3170 -3772
rect -9469 -3852 -3254 -3788
rect -3190 -3852 -3170 -3788
rect -9469 -3868 -3170 -3852
rect -9469 -3932 -3254 -3868
rect -3190 -3932 -3170 -3868
rect -9469 -3948 -3170 -3932
rect -9469 -4012 -3254 -3948
rect -3190 -4012 -3170 -3948
rect -9469 -4028 -3170 -4012
rect -9469 -4092 -3254 -4028
rect -3190 -4092 -3170 -4028
rect -9469 -4108 -3170 -4092
rect -9469 -4172 -3254 -4108
rect -3190 -4172 -3170 -4108
rect -9469 -4188 -3170 -4172
rect -9469 -4252 -3254 -4188
rect -3190 -4252 -3170 -4188
rect -9469 -4268 -3170 -4252
rect -9469 -4332 -3254 -4268
rect -3190 -4332 -3170 -4268
rect -9469 -4348 -3170 -4332
rect -9469 -4412 -3254 -4348
rect -3190 -4412 -3170 -4348
rect -9469 -4428 -3170 -4412
rect -9469 -4492 -3254 -4428
rect -3190 -4492 -3170 -4428
rect -9469 -4508 -3170 -4492
rect -9469 -4572 -3254 -4508
rect -3190 -4572 -3170 -4508
rect -9469 -4588 -3170 -4572
rect -9469 -4652 -3254 -4588
rect -3190 -4652 -3170 -4588
rect -9469 -4668 -3170 -4652
rect -9469 -4732 -3254 -4668
rect -3190 -4732 -3170 -4668
rect -9469 -4748 -3170 -4732
rect -9469 -4812 -3254 -4748
rect -3190 -4812 -3170 -4748
rect -9469 -4828 -3170 -4812
rect -9469 -4892 -3254 -4828
rect -3190 -4892 -3170 -4828
rect -9469 -4908 -3170 -4892
rect -9469 -4972 -3254 -4908
rect -3190 -4972 -3170 -4908
rect -9469 -4988 -3170 -4972
rect -9469 -5052 -3254 -4988
rect -3190 -5052 -3170 -4988
rect -9469 -5068 -3170 -5052
rect -9469 -5132 -3254 -5068
rect -3190 -5132 -3170 -5068
rect -9469 -5148 -3170 -5132
rect -9469 -5212 -3254 -5148
rect -3190 -5212 -3170 -5148
rect -9469 -5228 -3170 -5212
rect -9469 -5292 -3254 -5228
rect -3190 -5292 -3170 -5228
rect -9469 -5308 -3170 -5292
rect -9469 -5372 -3254 -5308
rect -3190 -5372 -3170 -5308
rect -9469 -5388 -3170 -5372
rect -9469 -5452 -3254 -5388
rect -3190 -5452 -3170 -5388
rect -9469 -5468 -3170 -5452
rect -9469 -5532 -3254 -5468
rect -3190 -5532 -3170 -5468
rect -9469 -5548 -3170 -5532
rect -9469 -5612 -3254 -5548
rect -3190 -5612 -3170 -5548
rect -9469 -5628 -3170 -5612
rect -9469 -5692 -3254 -5628
rect -3190 -5692 -3170 -5628
rect -9469 -5708 -3170 -5692
rect -9469 -5772 -3254 -5708
rect -3190 -5772 -3170 -5708
rect -9469 -5788 -3170 -5772
rect -9469 -5852 -3254 -5788
rect -3190 -5852 -3170 -5788
rect -9469 -5868 -3170 -5852
rect -9469 -5932 -3254 -5868
rect -3190 -5932 -3170 -5868
rect -9469 -5948 -3170 -5932
rect -9469 -6012 -3254 -5948
rect -3190 -6012 -3170 -5948
rect -9469 -6028 -3170 -6012
rect -9469 -6092 -3254 -6028
rect -3190 -6092 -3170 -6028
rect -9469 -6108 -3170 -6092
rect -9469 -6172 -3254 -6108
rect -3190 -6172 -3170 -6108
rect -9469 -6188 -3170 -6172
rect -9469 -6252 -3254 -6188
rect -3190 -6252 -3170 -6188
rect -9469 -6268 -3170 -6252
rect -9469 -6332 -3254 -6268
rect -3190 -6332 -3170 -6268
rect -9469 -6348 -3170 -6332
rect -9469 -6412 -3254 -6348
rect -3190 -6412 -3170 -6348
rect -9469 -6428 -3170 -6412
rect -9469 -6492 -3254 -6428
rect -3190 -6492 -3170 -6428
rect -9469 -6508 -3170 -6492
rect -9469 -6572 -3254 -6508
rect -3190 -6572 -3170 -6508
rect -9469 -6588 -3170 -6572
rect -9469 -6652 -3254 -6588
rect -3190 -6652 -3170 -6588
rect -9469 -6668 -3170 -6652
rect -9469 -6732 -3254 -6668
rect -3190 -6732 -3170 -6668
rect -9469 -6748 -3170 -6732
rect -9469 -6812 -3254 -6748
rect -3190 -6812 -3170 -6748
rect -9469 -6828 -3170 -6812
rect -9469 -6892 -3254 -6828
rect -3190 -6892 -3170 -6828
rect -9469 -6908 -3170 -6892
rect -9469 -6972 -3254 -6908
rect -3190 -6972 -3170 -6908
rect -9469 -6988 -3170 -6972
rect -9469 -7052 -3254 -6988
rect -3190 -7052 -3170 -6988
rect -9469 -7068 -3170 -7052
rect -9469 -7132 -3254 -7068
rect -3190 -7132 -3170 -7068
rect -9469 -7148 -3170 -7132
rect -9469 -7212 -3254 -7148
rect -3190 -7212 -3170 -7148
rect -9469 -7228 -3170 -7212
rect -9469 -7292 -3254 -7228
rect -3190 -7292 -3170 -7228
rect -9469 -7308 -3170 -7292
rect -9469 -7372 -3254 -7308
rect -3190 -7372 -3170 -7308
rect -9469 -7388 -3170 -7372
rect -9469 -7452 -3254 -7388
rect -3190 -7452 -3170 -7388
rect -9469 -7468 -3170 -7452
rect -9469 -7532 -3254 -7468
rect -3190 -7532 -3170 -7468
rect -9469 -7548 -3170 -7532
rect -9469 -7612 -3254 -7548
rect -3190 -7612 -3170 -7548
rect -9469 -7628 -3170 -7612
rect -9469 -7692 -3254 -7628
rect -3190 -7692 -3170 -7628
rect -9469 -7708 -3170 -7692
rect -9469 -7772 -3254 -7708
rect -3190 -7772 -3170 -7708
rect -9469 -7788 -3170 -7772
rect -9469 -7852 -3254 -7788
rect -3190 -7852 -3170 -7788
rect -9469 -7868 -3170 -7852
rect -9469 -7932 -3254 -7868
rect -3190 -7932 -3170 -7868
rect -9469 -7948 -3170 -7932
rect -9469 -8012 -3254 -7948
rect -3190 -8012 -3170 -7948
rect -9469 -8028 -3170 -8012
rect -9469 -8092 -3254 -8028
rect -3190 -8092 -3170 -8028
rect -9469 -8108 -3170 -8092
rect -9469 -8172 -3254 -8108
rect -3190 -8172 -3170 -8108
rect -9469 -8188 -3170 -8172
rect -9469 -8252 -3254 -8188
rect -3190 -8252 -3170 -8188
rect -9469 -8268 -3170 -8252
rect -9469 -8332 -3254 -8268
rect -3190 -8332 -3170 -8268
rect -9469 -8348 -3170 -8332
rect -9469 -8412 -3254 -8348
rect -3190 -8412 -3170 -8348
rect -9469 -8428 -3170 -8412
rect -9469 -8492 -3254 -8428
rect -3190 -8492 -3170 -8428
rect -9469 -8508 -3170 -8492
rect -9469 -8572 -3254 -8508
rect -3190 -8572 -3170 -8508
rect -9469 -8588 -3170 -8572
rect -9469 -8652 -3254 -8588
rect -3190 -8652 -3170 -8588
rect -9469 -8668 -3170 -8652
rect -9469 -8732 -3254 -8668
rect -3190 -8732 -3170 -8668
rect -9469 -8748 -3170 -8732
rect -9469 -8812 -3254 -8748
rect -3190 -8812 -3170 -8748
rect -9469 -8828 -3170 -8812
rect -9469 -8892 -3254 -8828
rect -3190 -8892 -3170 -8828
rect -9469 -8908 -3170 -8892
rect -9469 -8972 -3254 -8908
rect -3190 -8972 -3170 -8908
rect -9469 -8988 -3170 -8972
rect -9469 -9052 -3254 -8988
rect -3190 -9052 -3170 -8988
rect -9469 -9068 -3170 -9052
rect -9469 -9132 -3254 -9068
rect -3190 -9132 -3170 -9068
rect -9469 -9148 -3170 -9132
rect -9469 -9212 -3254 -9148
rect -3190 -9212 -3170 -9148
rect -9469 -9228 -3170 -9212
rect -9469 -9292 -3254 -9228
rect -3190 -9292 -3170 -9228
rect -9469 -9308 -3170 -9292
rect -9469 -9372 -3254 -9308
rect -3190 -9372 -3170 -9308
rect -9469 -9400 -3170 -9372
rect -3150 -3228 3149 -3200
rect -3150 -3292 3065 -3228
rect 3129 -3292 3149 -3228
rect -3150 -3308 3149 -3292
rect -3150 -3372 3065 -3308
rect 3129 -3372 3149 -3308
rect -3150 -3388 3149 -3372
rect -3150 -3452 3065 -3388
rect 3129 -3452 3149 -3388
rect -3150 -3468 3149 -3452
rect -3150 -3532 3065 -3468
rect 3129 -3532 3149 -3468
rect -3150 -3548 3149 -3532
rect -3150 -3612 3065 -3548
rect 3129 -3612 3149 -3548
rect -3150 -3628 3149 -3612
rect -3150 -3692 3065 -3628
rect 3129 -3692 3149 -3628
rect -3150 -3708 3149 -3692
rect -3150 -3772 3065 -3708
rect 3129 -3772 3149 -3708
rect -3150 -3788 3149 -3772
rect -3150 -3852 3065 -3788
rect 3129 -3852 3149 -3788
rect -3150 -3868 3149 -3852
rect -3150 -3932 3065 -3868
rect 3129 -3932 3149 -3868
rect -3150 -3948 3149 -3932
rect -3150 -4012 3065 -3948
rect 3129 -4012 3149 -3948
rect -3150 -4028 3149 -4012
rect -3150 -4092 3065 -4028
rect 3129 -4092 3149 -4028
rect -3150 -4108 3149 -4092
rect -3150 -4172 3065 -4108
rect 3129 -4172 3149 -4108
rect -3150 -4188 3149 -4172
rect -3150 -4252 3065 -4188
rect 3129 -4252 3149 -4188
rect -3150 -4268 3149 -4252
rect -3150 -4332 3065 -4268
rect 3129 -4332 3149 -4268
rect -3150 -4348 3149 -4332
rect -3150 -4412 3065 -4348
rect 3129 -4412 3149 -4348
rect -3150 -4428 3149 -4412
rect -3150 -4492 3065 -4428
rect 3129 -4492 3149 -4428
rect -3150 -4508 3149 -4492
rect -3150 -4572 3065 -4508
rect 3129 -4572 3149 -4508
rect -3150 -4588 3149 -4572
rect -3150 -4652 3065 -4588
rect 3129 -4652 3149 -4588
rect -3150 -4668 3149 -4652
rect -3150 -4732 3065 -4668
rect 3129 -4732 3149 -4668
rect -3150 -4748 3149 -4732
rect -3150 -4812 3065 -4748
rect 3129 -4812 3149 -4748
rect -3150 -4828 3149 -4812
rect -3150 -4892 3065 -4828
rect 3129 -4892 3149 -4828
rect -3150 -4908 3149 -4892
rect -3150 -4972 3065 -4908
rect 3129 -4972 3149 -4908
rect -3150 -4988 3149 -4972
rect -3150 -5052 3065 -4988
rect 3129 -5052 3149 -4988
rect -3150 -5068 3149 -5052
rect -3150 -5132 3065 -5068
rect 3129 -5132 3149 -5068
rect -3150 -5148 3149 -5132
rect -3150 -5212 3065 -5148
rect 3129 -5212 3149 -5148
rect -3150 -5228 3149 -5212
rect -3150 -5292 3065 -5228
rect 3129 -5292 3149 -5228
rect -3150 -5308 3149 -5292
rect -3150 -5372 3065 -5308
rect 3129 -5372 3149 -5308
rect -3150 -5388 3149 -5372
rect -3150 -5452 3065 -5388
rect 3129 -5452 3149 -5388
rect -3150 -5468 3149 -5452
rect -3150 -5532 3065 -5468
rect 3129 -5532 3149 -5468
rect -3150 -5548 3149 -5532
rect -3150 -5612 3065 -5548
rect 3129 -5612 3149 -5548
rect -3150 -5628 3149 -5612
rect -3150 -5692 3065 -5628
rect 3129 -5692 3149 -5628
rect -3150 -5708 3149 -5692
rect -3150 -5772 3065 -5708
rect 3129 -5772 3149 -5708
rect -3150 -5788 3149 -5772
rect -3150 -5852 3065 -5788
rect 3129 -5852 3149 -5788
rect -3150 -5868 3149 -5852
rect -3150 -5932 3065 -5868
rect 3129 -5932 3149 -5868
rect -3150 -5948 3149 -5932
rect -3150 -6012 3065 -5948
rect 3129 -6012 3149 -5948
rect -3150 -6028 3149 -6012
rect -3150 -6092 3065 -6028
rect 3129 -6092 3149 -6028
rect -3150 -6108 3149 -6092
rect -3150 -6172 3065 -6108
rect 3129 -6172 3149 -6108
rect -3150 -6188 3149 -6172
rect -3150 -6252 3065 -6188
rect 3129 -6252 3149 -6188
rect -3150 -6268 3149 -6252
rect -3150 -6332 3065 -6268
rect 3129 -6332 3149 -6268
rect -3150 -6348 3149 -6332
rect -3150 -6412 3065 -6348
rect 3129 -6412 3149 -6348
rect -3150 -6428 3149 -6412
rect -3150 -6492 3065 -6428
rect 3129 -6492 3149 -6428
rect -3150 -6508 3149 -6492
rect -3150 -6572 3065 -6508
rect 3129 -6572 3149 -6508
rect -3150 -6588 3149 -6572
rect -3150 -6652 3065 -6588
rect 3129 -6652 3149 -6588
rect -3150 -6668 3149 -6652
rect -3150 -6732 3065 -6668
rect 3129 -6732 3149 -6668
rect -3150 -6748 3149 -6732
rect -3150 -6812 3065 -6748
rect 3129 -6812 3149 -6748
rect -3150 -6828 3149 -6812
rect -3150 -6892 3065 -6828
rect 3129 -6892 3149 -6828
rect -3150 -6908 3149 -6892
rect -3150 -6972 3065 -6908
rect 3129 -6972 3149 -6908
rect -3150 -6988 3149 -6972
rect -3150 -7052 3065 -6988
rect 3129 -7052 3149 -6988
rect -3150 -7068 3149 -7052
rect -3150 -7132 3065 -7068
rect 3129 -7132 3149 -7068
rect -3150 -7148 3149 -7132
rect -3150 -7212 3065 -7148
rect 3129 -7212 3149 -7148
rect -3150 -7228 3149 -7212
rect -3150 -7292 3065 -7228
rect 3129 -7292 3149 -7228
rect -3150 -7308 3149 -7292
rect -3150 -7372 3065 -7308
rect 3129 -7372 3149 -7308
rect -3150 -7388 3149 -7372
rect -3150 -7452 3065 -7388
rect 3129 -7452 3149 -7388
rect -3150 -7468 3149 -7452
rect -3150 -7532 3065 -7468
rect 3129 -7532 3149 -7468
rect -3150 -7548 3149 -7532
rect -3150 -7612 3065 -7548
rect 3129 -7612 3149 -7548
rect -3150 -7628 3149 -7612
rect -3150 -7692 3065 -7628
rect 3129 -7692 3149 -7628
rect -3150 -7708 3149 -7692
rect -3150 -7772 3065 -7708
rect 3129 -7772 3149 -7708
rect -3150 -7788 3149 -7772
rect -3150 -7852 3065 -7788
rect 3129 -7852 3149 -7788
rect -3150 -7868 3149 -7852
rect -3150 -7932 3065 -7868
rect 3129 -7932 3149 -7868
rect -3150 -7948 3149 -7932
rect -3150 -8012 3065 -7948
rect 3129 -8012 3149 -7948
rect -3150 -8028 3149 -8012
rect -3150 -8092 3065 -8028
rect 3129 -8092 3149 -8028
rect -3150 -8108 3149 -8092
rect -3150 -8172 3065 -8108
rect 3129 -8172 3149 -8108
rect -3150 -8188 3149 -8172
rect -3150 -8252 3065 -8188
rect 3129 -8252 3149 -8188
rect -3150 -8268 3149 -8252
rect -3150 -8332 3065 -8268
rect 3129 -8332 3149 -8268
rect -3150 -8348 3149 -8332
rect -3150 -8412 3065 -8348
rect 3129 -8412 3149 -8348
rect -3150 -8428 3149 -8412
rect -3150 -8492 3065 -8428
rect 3129 -8492 3149 -8428
rect -3150 -8508 3149 -8492
rect -3150 -8572 3065 -8508
rect 3129 -8572 3149 -8508
rect -3150 -8588 3149 -8572
rect -3150 -8652 3065 -8588
rect 3129 -8652 3149 -8588
rect -3150 -8668 3149 -8652
rect -3150 -8732 3065 -8668
rect 3129 -8732 3149 -8668
rect -3150 -8748 3149 -8732
rect -3150 -8812 3065 -8748
rect 3129 -8812 3149 -8748
rect -3150 -8828 3149 -8812
rect -3150 -8892 3065 -8828
rect 3129 -8892 3149 -8828
rect -3150 -8908 3149 -8892
rect -3150 -8972 3065 -8908
rect 3129 -8972 3149 -8908
rect -3150 -8988 3149 -8972
rect -3150 -9052 3065 -8988
rect 3129 -9052 3149 -8988
rect -3150 -9068 3149 -9052
rect -3150 -9132 3065 -9068
rect 3129 -9132 3149 -9068
rect -3150 -9148 3149 -9132
rect -3150 -9212 3065 -9148
rect 3129 -9212 3149 -9148
rect -3150 -9228 3149 -9212
rect -3150 -9292 3065 -9228
rect 3129 -9292 3149 -9228
rect -3150 -9308 3149 -9292
rect -3150 -9372 3065 -9308
rect 3129 -9372 3149 -9308
rect -3150 -9400 3149 -9372
rect 3169 -3228 9468 -3200
rect 3169 -3292 9384 -3228
rect 9448 -3292 9468 -3228
rect 3169 -3308 9468 -3292
rect 3169 -3372 9384 -3308
rect 9448 -3372 9468 -3308
rect 3169 -3388 9468 -3372
rect 3169 -3452 9384 -3388
rect 9448 -3452 9468 -3388
rect 3169 -3468 9468 -3452
rect 3169 -3532 9384 -3468
rect 9448 -3532 9468 -3468
rect 3169 -3548 9468 -3532
rect 3169 -3612 9384 -3548
rect 9448 -3612 9468 -3548
rect 3169 -3628 9468 -3612
rect 3169 -3692 9384 -3628
rect 9448 -3692 9468 -3628
rect 3169 -3708 9468 -3692
rect 3169 -3772 9384 -3708
rect 9448 -3772 9468 -3708
rect 3169 -3788 9468 -3772
rect 3169 -3852 9384 -3788
rect 9448 -3852 9468 -3788
rect 3169 -3868 9468 -3852
rect 3169 -3932 9384 -3868
rect 9448 -3932 9468 -3868
rect 3169 -3948 9468 -3932
rect 3169 -4012 9384 -3948
rect 9448 -4012 9468 -3948
rect 3169 -4028 9468 -4012
rect 3169 -4092 9384 -4028
rect 9448 -4092 9468 -4028
rect 3169 -4108 9468 -4092
rect 3169 -4172 9384 -4108
rect 9448 -4172 9468 -4108
rect 3169 -4188 9468 -4172
rect 3169 -4252 9384 -4188
rect 9448 -4252 9468 -4188
rect 3169 -4268 9468 -4252
rect 3169 -4332 9384 -4268
rect 9448 -4332 9468 -4268
rect 3169 -4348 9468 -4332
rect 3169 -4412 9384 -4348
rect 9448 -4412 9468 -4348
rect 3169 -4428 9468 -4412
rect 3169 -4492 9384 -4428
rect 9448 -4492 9468 -4428
rect 3169 -4508 9468 -4492
rect 3169 -4572 9384 -4508
rect 9448 -4572 9468 -4508
rect 3169 -4588 9468 -4572
rect 3169 -4652 9384 -4588
rect 9448 -4652 9468 -4588
rect 3169 -4668 9468 -4652
rect 3169 -4732 9384 -4668
rect 9448 -4732 9468 -4668
rect 3169 -4748 9468 -4732
rect 3169 -4812 9384 -4748
rect 9448 -4812 9468 -4748
rect 3169 -4828 9468 -4812
rect 3169 -4892 9384 -4828
rect 9448 -4892 9468 -4828
rect 3169 -4908 9468 -4892
rect 3169 -4972 9384 -4908
rect 9448 -4972 9468 -4908
rect 3169 -4988 9468 -4972
rect 3169 -5052 9384 -4988
rect 9448 -5052 9468 -4988
rect 3169 -5068 9468 -5052
rect 3169 -5132 9384 -5068
rect 9448 -5132 9468 -5068
rect 3169 -5148 9468 -5132
rect 3169 -5212 9384 -5148
rect 9448 -5212 9468 -5148
rect 3169 -5228 9468 -5212
rect 3169 -5292 9384 -5228
rect 9448 -5292 9468 -5228
rect 3169 -5308 9468 -5292
rect 3169 -5372 9384 -5308
rect 9448 -5372 9468 -5308
rect 3169 -5388 9468 -5372
rect 3169 -5452 9384 -5388
rect 9448 -5452 9468 -5388
rect 3169 -5468 9468 -5452
rect 3169 -5532 9384 -5468
rect 9448 -5532 9468 -5468
rect 3169 -5548 9468 -5532
rect 3169 -5612 9384 -5548
rect 9448 -5612 9468 -5548
rect 3169 -5628 9468 -5612
rect 3169 -5692 9384 -5628
rect 9448 -5692 9468 -5628
rect 3169 -5708 9468 -5692
rect 3169 -5772 9384 -5708
rect 9448 -5772 9468 -5708
rect 3169 -5788 9468 -5772
rect 3169 -5852 9384 -5788
rect 9448 -5852 9468 -5788
rect 3169 -5868 9468 -5852
rect 3169 -5932 9384 -5868
rect 9448 -5932 9468 -5868
rect 3169 -5948 9468 -5932
rect 3169 -6012 9384 -5948
rect 9448 -6012 9468 -5948
rect 3169 -6028 9468 -6012
rect 3169 -6092 9384 -6028
rect 9448 -6092 9468 -6028
rect 3169 -6108 9468 -6092
rect 3169 -6172 9384 -6108
rect 9448 -6172 9468 -6108
rect 3169 -6188 9468 -6172
rect 3169 -6252 9384 -6188
rect 9448 -6252 9468 -6188
rect 3169 -6268 9468 -6252
rect 3169 -6332 9384 -6268
rect 9448 -6332 9468 -6268
rect 3169 -6348 9468 -6332
rect 3169 -6412 9384 -6348
rect 9448 -6412 9468 -6348
rect 3169 -6428 9468 -6412
rect 3169 -6492 9384 -6428
rect 9448 -6492 9468 -6428
rect 3169 -6508 9468 -6492
rect 3169 -6572 9384 -6508
rect 9448 -6572 9468 -6508
rect 3169 -6588 9468 -6572
rect 3169 -6652 9384 -6588
rect 9448 -6652 9468 -6588
rect 3169 -6668 9468 -6652
rect 3169 -6732 9384 -6668
rect 9448 -6732 9468 -6668
rect 3169 -6748 9468 -6732
rect 3169 -6812 9384 -6748
rect 9448 -6812 9468 -6748
rect 3169 -6828 9468 -6812
rect 3169 -6892 9384 -6828
rect 9448 -6892 9468 -6828
rect 3169 -6908 9468 -6892
rect 3169 -6972 9384 -6908
rect 9448 -6972 9468 -6908
rect 3169 -6988 9468 -6972
rect 3169 -7052 9384 -6988
rect 9448 -7052 9468 -6988
rect 3169 -7068 9468 -7052
rect 3169 -7132 9384 -7068
rect 9448 -7132 9468 -7068
rect 3169 -7148 9468 -7132
rect 3169 -7212 9384 -7148
rect 9448 -7212 9468 -7148
rect 3169 -7228 9468 -7212
rect 3169 -7292 9384 -7228
rect 9448 -7292 9468 -7228
rect 3169 -7308 9468 -7292
rect 3169 -7372 9384 -7308
rect 9448 -7372 9468 -7308
rect 3169 -7388 9468 -7372
rect 3169 -7452 9384 -7388
rect 9448 -7452 9468 -7388
rect 3169 -7468 9468 -7452
rect 3169 -7532 9384 -7468
rect 9448 -7532 9468 -7468
rect 3169 -7548 9468 -7532
rect 3169 -7612 9384 -7548
rect 9448 -7612 9468 -7548
rect 3169 -7628 9468 -7612
rect 3169 -7692 9384 -7628
rect 9448 -7692 9468 -7628
rect 3169 -7708 9468 -7692
rect 3169 -7772 9384 -7708
rect 9448 -7772 9468 -7708
rect 3169 -7788 9468 -7772
rect 3169 -7852 9384 -7788
rect 9448 -7852 9468 -7788
rect 3169 -7868 9468 -7852
rect 3169 -7932 9384 -7868
rect 9448 -7932 9468 -7868
rect 3169 -7948 9468 -7932
rect 3169 -8012 9384 -7948
rect 9448 -8012 9468 -7948
rect 3169 -8028 9468 -8012
rect 3169 -8092 9384 -8028
rect 9448 -8092 9468 -8028
rect 3169 -8108 9468 -8092
rect 3169 -8172 9384 -8108
rect 9448 -8172 9468 -8108
rect 3169 -8188 9468 -8172
rect 3169 -8252 9384 -8188
rect 9448 -8252 9468 -8188
rect 3169 -8268 9468 -8252
rect 3169 -8332 9384 -8268
rect 9448 -8332 9468 -8268
rect 3169 -8348 9468 -8332
rect 3169 -8412 9384 -8348
rect 9448 -8412 9468 -8348
rect 3169 -8428 9468 -8412
rect 3169 -8492 9384 -8428
rect 9448 -8492 9468 -8428
rect 3169 -8508 9468 -8492
rect 3169 -8572 9384 -8508
rect 9448 -8572 9468 -8508
rect 3169 -8588 9468 -8572
rect 3169 -8652 9384 -8588
rect 9448 -8652 9468 -8588
rect 3169 -8668 9468 -8652
rect 3169 -8732 9384 -8668
rect 9448 -8732 9468 -8668
rect 3169 -8748 9468 -8732
rect 3169 -8812 9384 -8748
rect 9448 -8812 9468 -8748
rect 3169 -8828 9468 -8812
rect 3169 -8892 9384 -8828
rect 9448 -8892 9468 -8828
rect 3169 -8908 9468 -8892
rect 3169 -8972 9384 -8908
rect 9448 -8972 9468 -8908
rect 3169 -8988 9468 -8972
rect 3169 -9052 9384 -8988
rect 9448 -9052 9468 -8988
rect 3169 -9068 9468 -9052
rect 3169 -9132 9384 -9068
rect 9448 -9132 9468 -9068
rect 3169 -9148 9468 -9132
rect 3169 -9212 9384 -9148
rect 9448 -9212 9468 -9148
rect 3169 -9228 9468 -9212
rect 3169 -9292 9384 -9228
rect 9448 -9292 9468 -9228
rect 3169 -9308 9468 -9292
rect 3169 -9372 9384 -9308
rect 9448 -9372 9468 -9308
rect 3169 -9400 9468 -9372
rect 9488 -3228 15787 -3200
rect 9488 -3292 15703 -3228
rect 15767 -3292 15787 -3228
rect 9488 -3308 15787 -3292
rect 9488 -3372 15703 -3308
rect 15767 -3372 15787 -3308
rect 9488 -3388 15787 -3372
rect 9488 -3452 15703 -3388
rect 15767 -3452 15787 -3388
rect 9488 -3468 15787 -3452
rect 9488 -3532 15703 -3468
rect 15767 -3532 15787 -3468
rect 9488 -3548 15787 -3532
rect 9488 -3612 15703 -3548
rect 15767 -3612 15787 -3548
rect 9488 -3628 15787 -3612
rect 9488 -3692 15703 -3628
rect 15767 -3692 15787 -3628
rect 9488 -3708 15787 -3692
rect 9488 -3772 15703 -3708
rect 15767 -3772 15787 -3708
rect 9488 -3788 15787 -3772
rect 9488 -3852 15703 -3788
rect 15767 -3852 15787 -3788
rect 9488 -3868 15787 -3852
rect 9488 -3932 15703 -3868
rect 15767 -3932 15787 -3868
rect 9488 -3948 15787 -3932
rect 9488 -4012 15703 -3948
rect 15767 -4012 15787 -3948
rect 9488 -4028 15787 -4012
rect 9488 -4092 15703 -4028
rect 15767 -4092 15787 -4028
rect 9488 -4108 15787 -4092
rect 9488 -4172 15703 -4108
rect 15767 -4172 15787 -4108
rect 9488 -4188 15787 -4172
rect 9488 -4252 15703 -4188
rect 15767 -4252 15787 -4188
rect 9488 -4268 15787 -4252
rect 9488 -4332 15703 -4268
rect 15767 -4332 15787 -4268
rect 9488 -4348 15787 -4332
rect 9488 -4412 15703 -4348
rect 15767 -4412 15787 -4348
rect 9488 -4428 15787 -4412
rect 9488 -4492 15703 -4428
rect 15767 -4492 15787 -4428
rect 9488 -4508 15787 -4492
rect 9488 -4572 15703 -4508
rect 15767 -4572 15787 -4508
rect 9488 -4588 15787 -4572
rect 9488 -4652 15703 -4588
rect 15767 -4652 15787 -4588
rect 9488 -4668 15787 -4652
rect 9488 -4732 15703 -4668
rect 15767 -4732 15787 -4668
rect 9488 -4748 15787 -4732
rect 9488 -4812 15703 -4748
rect 15767 -4812 15787 -4748
rect 9488 -4828 15787 -4812
rect 9488 -4892 15703 -4828
rect 15767 -4892 15787 -4828
rect 9488 -4908 15787 -4892
rect 9488 -4972 15703 -4908
rect 15767 -4972 15787 -4908
rect 9488 -4988 15787 -4972
rect 9488 -5052 15703 -4988
rect 15767 -5052 15787 -4988
rect 9488 -5068 15787 -5052
rect 9488 -5132 15703 -5068
rect 15767 -5132 15787 -5068
rect 9488 -5148 15787 -5132
rect 9488 -5212 15703 -5148
rect 15767 -5212 15787 -5148
rect 9488 -5228 15787 -5212
rect 9488 -5292 15703 -5228
rect 15767 -5292 15787 -5228
rect 9488 -5308 15787 -5292
rect 9488 -5372 15703 -5308
rect 15767 -5372 15787 -5308
rect 9488 -5388 15787 -5372
rect 9488 -5452 15703 -5388
rect 15767 -5452 15787 -5388
rect 9488 -5468 15787 -5452
rect 9488 -5532 15703 -5468
rect 15767 -5532 15787 -5468
rect 9488 -5548 15787 -5532
rect 9488 -5612 15703 -5548
rect 15767 -5612 15787 -5548
rect 9488 -5628 15787 -5612
rect 9488 -5692 15703 -5628
rect 15767 -5692 15787 -5628
rect 9488 -5708 15787 -5692
rect 9488 -5772 15703 -5708
rect 15767 -5772 15787 -5708
rect 9488 -5788 15787 -5772
rect 9488 -5852 15703 -5788
rect 15767 -5852 15787 -5788
rect 9488 -5868 15787 -5852
rect 9488 -5932 15703 -5868
rect 15767 -5932 15787 -5868
rect 9488 -5948 15787 -5932
rect 9488 -6012 15703 -5948
rect 15767 -6012 15787 -5948
rect 9488 -6028 15787 -6012
rect 9488 -6092 15703 -6028
rect 15767 -6092 15787 -6028
rect 9488 -6108 15787 -6092
rect 9488 -6172 15703 -6108
rect 15767 -6172 15787 -6108
rect 9488 -6188 15787 -6172
rect 9488 -6252 15703 -6188
rect 15767 -6252 15787 -6188
rect 9488 -6268 15787 -6252
rect 9488 -6332 15703 -6268
rect 15767 -6332 15787 -6268
rect 9488 -6348 15787 -6332
rect 9488 -6412 15703 -6348
rect 15767 -6412 15787 -6348
rect 9488 -6428 15787 -6412
rect 9488 -6492 15703 -6428
rect 15767 -6492 15787 -6428
rect 9488 -6508 15787 -6492
rect 9488 -6572 15703 -6508
rect 15767 -6572 15787 -6508
rect 9488 -6588 15787 -6572
rect 9488 -6652 15703 -6588
rect 15767 -6652 15787 -6588
rect 9488 -6668 15787 -6652
rect 9488 -6732 15703 -6668
rect 15767 -6732 15787 -6668
rect 9488 -6748 15787 -6732
rect 9488 -6812 15703 -6748
rect 15767 -6812 15787 -6748
rect 9488 -6828 15787 -6812
rect 9488 -6892 15703 -6828
rect 15767 -6892 15787 -6828
rect 9488 -6908 15787 -6892
rect 9488 -6972 15703 -6908
rect 15767 -6972 15787 -6908
rect 9488 -6988 15787 -6972
rect 9488 -7052 15703 -6988
rect 15767 -7052 15787 -6988
rect 9488 -7068 15787 -7052
rect 9488 -7132 15703 -7068
rect 15767 -7132 15787 -7068
rect 9488 -7148 15787 -7132
rect 9488 -7212 15703 -7148
rect 15767 -7212 15787 -7148
rect 9488 -7228 15787 -7212
rect 9488 -7292 15703 -7228
rect 15767 -7292 15787 -7228
rect 9488 -7308 15787 -7292
rect 9488 -7372 15703 -7308
rect 15767 -7372 15787 -7308
rect 9488 -7388 15787 -7372
rect 9488 -7452 15703 -7388
rect 15767 -7452 15787 -7388
rect 9488 -7468 15787 -7452
rect 9488 -7532 15703 -7468
rect 15767 -7532 15787 -7468
rect 9488 -7548 15787 -7532
rect 9488 -7612 15703 -7548
rect 15767 -7612 15787 -7548
rect 9488 -7628 15787 -7612
rect 9488 -7692 15703 -7628
rect 15767 -7692 15787 -7628
rect 9488 -7708 15787 -7692
rect 9488 -7772 15703 -7708
rect 15767 -7772 15787 -7708
rect 9488 -7788 15787 -7772
rect 9488 -7852 15703 -7788
rect 15767 -7852 15787 -7788
rect 9488 -7868 15787 -7852
rect 9488 -7932 15703 -7868
rect 15767 -7932 15787 -7868
rect 9488 -7948 15787 -7932
rect 9488 -8012 15703 -7948
rect 15767 -8012 15787 -7948
rect 9488 -8028 15787 -8012
rect 9488 -8092 15703 -8028
rect 15767 -8092 15787 -8028
rect 9488 -8108 15787 -8092
rect 9488 -8172 15703 -8108
rect 15767 -8172 15787 -8108
rect 9488 -8188 15787 -8172
rect 9488 -8252 15703 -8188
rect 15767 -8252 15787 -8188
rect 9488 -8268 15787 -8252
rect 9488 -8332 15703 -8268
rect 15767 -8332 15787 -8268
rect 9488 -8348 15787 -8332
rect 9488 -8412 15703 -8348
rect 15767 -8412 15787 -8348
rect 9488 -8428 15787 -8412
rect 9488 -8492 15703 -8428
rect 15767 -8492 15787 -8428
rect 9488 -8508 15787 -8492
rect 9488 -8572 15703 -8508
rect 15767 -8572 15787 -8508
rect 9488 -8588 15787 -8572
rect 9488 -8652 15703 -8588
rect 15767 -8652 15787 -8588
rect 9488 -8668 15787 -8652
rect 9488 -8732 15703 -8668
rect 15767 -8732 15787 -8668
rect 9488 -8748 15787 -8732
rect 9488 -8812 15703 -8748
rect 15767 -8812 15787 -8748
rect 9488 -8828 15787 -8812
rect 9488 -8892 15703 -8828
rect 15767 -8892 15787 -8828
rect 9488 -8908 15787 -8892
rect 9488 -8972 15703 -8908
rect 15767 -8972 15787 -8908
rect 9488 -8988 15787 -8972
rect 9488 -9052 15703 -8988
rect 15767 -9052 15787 -8988
rect 9488 -9068 15787 -9052
rect 9488 -9132 15703 -9068
rect 15767 -9132 15787 -9068
rect 9488 -9148 15787 -9132
rect 9488 -9212 15703 -9148
rect 15767 -9212 15787 -9148
rect 9488 -9228 15787 -9212
rect 9488 -9292 15703 -9228
rect 15767 -9292 15787 -9228
rect 9488 -9308 15787 -9292
rect 9488 -9372 15703 -9308
rect 15767 -9372 15787 -9308
rect 9488 -9400 15787 -9372
rect 15807 -3228 22106 -3200
rect 15807 -3292 22022 -3228
rect 22086 -3292 22106 -3228
rect 15807 -3308 22106 -3292
rect 15807 -3372 22022 -3308
rect 22086 -3372 22106 -3308
rect 15807 -3388 22106 -3372
rect 15807 -3452 22022 -3388
rect 22086 -3452 22106 -3388
rect 15807 -3468 22106 -3452
rect 15807 -3532 22022 -3468
rect 22086 -3532 22106 -3468
rect 15807 -3548 22106 -3532
rect 15807 -3612 22022 -3548
rect 22086 -3612 22106 -3548
rect 15807 -3628 22106 -3612
rect 15807 -3692 22022 -3628
rect 22086 -3692 22106 -3628
rect 15807 -3708 22106 -3692
rect 15807 -3772 22022 -3708
rect 22086 -3772 22106 -3708
rect 15807 -3788 22106 -3772
rect 15807 -3852 22022 -3788
rect 22086 -3852 22106 -3788
rect 15807 -3868 22106 -3852
rect 15807 -3932 22022 -3868
rect 22086 -3932 22106 -3868
rect 15807 -3948 22106 -3932
rect 15807 -4012 22022 -3948
rect 22086 -4012 22106 -3948
rect 15807 -4028 22106 -4012
rect 15807 -4092 22022 -4028
rect 22086 -4092 22106 -4028
rect 15807 -4108 22106 -4092
rect 15807 -4172 22022 -4108
rect 22086 -4172 22106 -4108
rect 15807 -4188 22106 -4172
rect 15807 -4252 22022 -4188
rect 22086 -4252 22106 -4188
rect 15807 -4268 22106 -4252
rect 15807 -4332 22022 -4268
rect 22086 -4332 22106 -4268
rect 15807 -4348 22106 -4332
rect 15807 -4412 22022 -4348
rect 22086 -4412 22106 -4348
rect 15807 -4428 22106 -4412
rect 15807 -4492 22022 -4428
rect 22086 -4492 22106 -4428
rect 15807 -4508 22106 -4492
rect 15807 -4572 22022 -4508
rect 22086 -4572 22106 -4508
rect 15807 -4588 22106 -4572
rect 15807 -4652 22022 -4588
rect 22086 -4652 22106 -4588
rect 15807 -4668 22106 -4652
rect 15807 -4732 22022 -4668
rect 22086 -4732 22106 -4668
rect 15807 -4748 22106 -4732
rect 15807 -4812 22022 -4748
rect 22086 -4812 22106 -4748
rect 15807 -4828 22106 -4812
rect 15807 -4892 22022 -4828
rect 22086 -4892 22106 -4828
rect 15807 -4908 22106 -4892
rect 15807 -4972 22022 -4908
rect 22086 -4972 22106 -4908
rect 15807 -4988 22106 -4972
rect 15807 -5052 22022 -4988
rect 22086 -5052 22106 -4988
rect 15807 -5068 22106 -5052
rect 15807 -5132 22022 -5068
rect 22086 -5132 22106 -5068
rect 15807 -5148 22106 -5132
rect 15807 -5212 22022 -5148
rect 22086 -5212 22106 -5148
rect 15807 -5228 22106 -5212
rect 15807 -5292 22022 -5228
rect 22086 -5292 22106 -5228
rect 15807 -5308 22106 -5292
rect 15807 -5372 22022 -5308
rect 22086 -5372 22106 -5308
rect 15807 -5388 22106 -5372
rect 15807 -5452 22022 -5388
rect 22086 -5452 22106 -5388
rect 15807 -5468 22106 -5452
rect 15807 -5532 22022 -5468
rect 22086 -5532 22106 -5468
rect 15807 -5548 22106 -5532
rect 15807 -5612 22022 -5548
rect 22086 -5612 22106 -5548
rect 15807 -5628 22106 -5612
rect 15807 -5692 22022 -5628
rect 22086 -5692 22106 -5628
rect 15807 -5708 22106 -5692
rect 15807 -5772 22022 -5708
rect 22086 -5772 22106 -5708
rect 15807 -5788 22106 -5772
rect 15807 -5852 22022 -5788
rect 22086 -5852 22106 -5788
rect 15807 -5868 22106 -5852
rect 15807 -5932 22022 -5868
rect 22086 -5932 22106 -5868
rect 15807 -5948 22106 -5932
rect 15807 -6012 22022 -5948
rect 22086 -6012 22106 -5948
rect 15807 -6028 22106 -6012
rect 15807 -6092 22022 -6028
rect 22086 -6092 22106 -6028
rect 15807 -6108 22106 -6092
rect 15807 -6172 22022 -6108
rect 22086 -6172 22106 -6108
rect 15807 -6188 22106 -6172
rect 15807 -6252 22022 -6188
rect 22086 -6252 22106 -6188
rect 15807 -6268 22106 -6252
rect 15807 -6332 22022 -6268
rect 22086 -6332 22106 -6268
rect 15807 -6348 22106 -6332
rect 15807 -6412 22022 -6348
rect 22086 -6412 22106 -6348
rect 15807 -6428 22106 -6412
rect 15807 -6492 22022 -6428
rect 22086 -6492 22106 -6428
rect 15807 -6508 22106 -6492
rect 15807 -6572 22022 -6508
rect 22086 -6572 22106 -6508
rect 15807 -6588 22106 -6572
rect 15807 -6652 22022 -6588
rect 22086 -6652 22106 -6588
rect 15807 -6668 22106 -6652
rect 15807 -6732 22022 -6668
rect 22086 -6732 22106 -6668
rect 15807 -6748 22106 -6732
rect 15807 -6812 22022 -6748
rect 22086 -6812 22106 -6748
rect 15807 -6828 22106 -6812
rect 15807 -6892 22022 -6828
rect 22086 -6892 22106 -6828
rect 15807 -6908 22106 -6892
rect 15807 -6972 22022 -6908
rect 22086 -6972 22106 -6908
rect 15807 -6988 22106 -6972
rect 15807 -7052 22022 -6988
rect 22086 -7052 22106 -6988
rect 15807 -7068 22106 -7052
rect 15807 -7132 22022 -7068
rect 22086 -7132 22106 -7068
rect 15807 -7148 22106 -7132
rect 15807 -7212 22022 -7148
rect 22086 -7212 22106 -7148
rect 15807 -7228 22106 -7212
rect 15807 -7292 22022 -7228
rect 22086 -7292 22106 -7228
rect 15807 -7308 22106 -7292
rect 15807 -7372 22022 -7308
rect 22086 -7372 22106 -7308
rect 15807 -7388 22106 -7372
rect 15807 -7452 22022 -7388
rect 22086 -7452 22106 -7388
rect 15807 -7468 22106 -7452
rect 15807 -7532 22022 -7468
rect 22086 -7532 22106 -7468
rect 15807 -7548 22106 -7532
rect 15807 -7612 22022 -7548
rect 22086 -7612 22106 -7548
rect 15807 -7628 22106 -7612
rect 15807 -7692 22022 -7628
rect 22086 -7692 22106 -7628
rect 15807 -7708 22106 -7692
rect 15807 -7772 22022 -7708
rect 22086 -7772 22106 -7708
rect 15807 -7788 22106 -7772
rect 15807 -7852 22022 -7788
rect 22086 -7852 22106 -7788
rect 15807 -7868 22106 -7852
rect 15807 -7932 22022 -7868
rect 22086 -7932 22106 -7868
rect 15807 -7948 22106 -7932
rect 15807 -8012 22022 -7948
rect 22086 -8012 22106 -7948
rect 15807 -8028 22106 -8012
rect 15807 -8092 22022 -8028
rect 22086 -8092 22106 -8028
rect 15807 -8108 22106 -8092
rect 15807 -8172 22022 -8108
rect 22086 -8172 22106 -8108
rect 15807 -8188 22106 -8172
rect 15807 -8252 22022 -8188
rect 22086 -8252 22106 -8188
rect 15807 -8268 22106 -8252
rect 15807 -8332 22022 -8268
rect 22086 -8332 22106 -8268
rect 15807 -8348 22106 -8332
rect 15807 -8412 22022 -8348
rect 22086 -8412 22106 -8348
rect 15807 -8428 22106 -8412
rect 15807 -8492 22022 -8428
rect 22086 -8492 22106 -8428
rect 15807 -8508 22106 -8492
rect 15807 -8572 22022 -8508
rect 22086 -8572 22106 -8508
rect 15807 -8588 22106 -8572
rect 15807 -8652 22022 -8588
rect 22086 -8652 22106 -8588
rect 15807 -8668 22106 -8652
rect 15807 -8732 22022 -8668
rect 22086 -8732 22106 -8668
rect 15807 -8748 22106 -8732
rect 15807 -8812 22022 -8748
rect 22086 -8812 22106 -8748
rect 15807 -8828 22106 -8812
rect 15807 -8892 22022 -8828
rect 22086 -8892 22106 -8828
rect 15807 -8908 22106 -8892
rect 15807 -8972 22022 -8908
rect 22086 -8972 22106 -8908
rect 15807 -8988 22106 -8972
rect 15807 -9052 22022 -8988
rect 22086 -9052 22106 -8988
rect 15807 -9068 22106 -9052
rect 15807 -9132 22022 -9068
rect 22086 -9132 22106 -9068
rect 15807 -9148 22106 -9132
rect 15807 -9212 22022 -9148
rect 22086 -9212 22106 -9148
rect 15807 -9228 22106 -9212
rect 15807 -9292 22022 -9228
rect 22086 -9292 22106 -9228
rect 15807 -9308 22106 -9292
rect 15807 -9372 22022 -9308
rect 22086 -9372 22106 -9308
rect 15807 -9400 22106 -9372
rect 22126 -3228 28425 -3200
rect 22126 -3292 28341 -3228
rect 28405 -3292 28425 -3228
rect 22126 -3308 28425 -3292
rect 22126 -3372 28341 -3308
rect 28405 -3372 28425 -3308
rect 22126 -3388 28425 -3372
rect 22126 -3452 28341 -3388
rect 28405 -3452 28425 -3388
rect 22126 -3468 28425 -3452
rect 22126 -3532 28341 -3468
rect 28405 -3532 28425 -3468
rect 22126 -3548 28425 -3532
rect 22126 -3612 28341 -3548
rect 28405 -3612 28425 -3548
rect 22126 -3628 28425 -3612
rect 22126 -3692 28341 -3628
rect 28405 -3692 28425 -3628
rect 22126 -3708 28425 -3692
rect 22126 -3772 28341 -3708
rect 28405 -3772 28425 -3708
rect 22126 -3788 28425 -3772
rect 22126 -3852 28341 -3788
rect 28405 -3852 28425 -3788
rect 22126 -3868 28425 -3852
rect 22126 -3932 28341 -3868
rect 28405 -3932 28425 -3868
rect 22126 -3948 28425 -3932
rect 22126 -4012 28341 -3948
rect 28405 -4012 28425 -3948
rect 22126 -4028 28425 -4012
rect 22126 -4092 28341 -4028
rect 28405 -4092 28425 -4028
rect 22126 -4108 28425 -4092
rect 22126 -4172 28341 -4108
rect 28405 -4172 28425 -4108
rect 22126 -4188 28425 -4172
rect 22126 -4252 28341 -4188
rect 28405 -4252 28425 -4188
rect 22126 -4268 28425 -4252
rect 22126 -4332 28341 -4268
rect 28405 -4332 28425 -4268
rect 22126 -4348 28425 -4332
rect 22126 -4412 28341 -4348
rect 28405 -4412 28425 -4348
rect 22126 -4428 28425 -4412
rect 22126 -4492 28341 -4428
rect 28405 -4492 28425 -4428
rect 22126 -4508 28425 -4492
rect 22126 -4572 28341 -4508
rect 28405 -4572 28425 -4508
rect 22126 -4588 28425 -4572
rect 22126 -4652 28341 -4588
rect 28405 -4652 28425 -4588
rect 22126 -4668 28425 -4652
rect 22126 -4732 28341 -4668
rect 28405 -4732 28425 -4668
rect 22126 -4748 28425 -4732
rect 22126 -4812 28341 -4748
rect 28405 -4812 28425 -4748
rect 22126 -4828 28425 -4812
rect 22126 -4892 28341 -4828
rect 28405 -4892 28425 -4828
rect 22126 -4908 28425 -4892
rect 22126 -4972 28341 -4908
rect 28405 -4972 28425 -4908
rect 22126 -4988 28425 -4972
rect 22126 -5052 28341 -4988
rect 28405 -5052 28425 -4988
rect 22126 -5068 28425 -5052
rect 22126 -5132 28341 -5068
rect 28405 -5132 28425 -5068
rect 22126 -5148 28425 -5132
rect 22126 -5212 28341 -5148
rect 28405 -5212 28425 -5148
rect 22126 -5228 28425 -5212
rect 22126 -5292 28341 -5228
rect 28405 -5292 28425 -5228
rect 22126 -5308 28425 -5292
rect 22126 -5372 28341 -5308
rect 28405 -5372 28425 -5308
rect 22126 -5388 28425 -5372
rect 22126 -5452 28341 -5388
rect 28405 -5452 28425 -5388
rect 22126 -5468 28425 -5452
rect 22126 -5532 28341 -5468
rect 28405 -5532 28425 -5468
rect 22126 -5548 28425 -5532
rect 22126 -5612 28341 -5548
rect 28405 -5612 28425 -5548
rect 22126 -5628 28425 -5612
rect 22126 -5692 28341 -5628
rect 28405 -5692 28425 -5628
rect 22126 -5708 28425 -5692
rect 22126 -5772 28341 -5708
rect 28405 -5772 28425 -5708
rect 22126 -5788 28425 -5772
rect 22126 -5852 28341 -5788
rect 28405 -5852 28425 -5788
rect 22126 -5868 28425 -5852
rect 22126 -5932 28341 -5868
rect 28405 -5932 28425 -5868
rect 22126 -5948 28425 -5932
rect 22126 -6012 28341 -5948
rect 28405 -6012 28425 -5948
rect 22126 -6028 28425 -6012
rect 22126 -6092 28341 -6028
rect 28405 -6092 28425 -6028
rect 22126 -6108 28425 -6092
rect 22126 -6172 28341 -6108
rect 28405 -6172 28425 -6108
rect 22126 -6188 28425 -6172
rect 22126 -6252 28341 -6188
rect 28405 -6252 28425 -6188
rect 22126 -6268 28425 -6252
rect 22126 -6332 28341 -6268
rect 28405 -6332 28425 -6268
rect 22126 -6348 28425 -6332
rect 22126 -6412 28341 -6348
rect 28405 -6412 28425 -6348
rect 22126 -6428 28425 -6412
rect 22126 -6492 28341 -6428
rect 28405 -6492 28425 -6428
rect 22126 -6508 28425 -6492
rect 22126 -6572 28341 -6508
rect 28405 -6572 28425 -6508
rect 22126 -6588 28425 -6572
rect 22126 -6652 28341 -6588
rect 28405 -6652 28425 -6588
rect 22126 -6668 28425 -6652
rect 22126 -6732 28341 -6668
rect 28405 -6732 28425 -6668
rect 22126 -6748 28425 -6732
rect 22126 -6812 28341 -6748
rect 28405 -6812 28425 -6748
rect 22126 -6828 28425 -6812
rect 22126 -6892 28341 -6828
rect 28405 -6892 28425 -6828
rect 22126 -6908 28425 -6892
rect 22126 -6972 28341 -6908
rect 28405 -6972 28425 -6908
rect 22126 -6988 28425 -6972
rect 22126 -7052 28341 -6988
rect 28405 -7052 28425 -6988
rect 22126 -7068 28425 -7052
rect 22126 -7132 28341 -7068
rect 28405 -7132 28425 -7068
rect 22126 -7148 28425 -7132
rect 22126 -7212 28341 -7148
rect 28405 -7212 28425 -7148
rect 22126 -7228 28425 -7212
rect 22126 -7292 28341 -7228
rect 28405 -7292 28425 -7228
rect 22126 -7308 28425 -7292
rect 22126 -7372 28341 -7308
rect 28405 -7372 28425 -7308
rect 22126 -7388 28425 -7372
rect 22126 -7452 28341 -7388
rect 28405 -7452 28425 -7388
rect 22126 -7468 28425 -7452
rect 22126 -7532 28341 -7468
rect 28405 -7532 28425 -7468
rect 22126 -7548 28425 -7532
rect 22126 -7612 28341 -7548
rect 28405 -7612 28425 -7548
rect 22126 -7628 28425 -7612
rect 22126 -7692 28341 -7628
rect 28405 -7692 28425 -7628
rect 22126 -7708 28425 -7692
rect 22126 -7772 28341 -7708
rect 28405 -7772 28425 -7708
rect 22126 -7788 28425 -7772
rect 22126 -7852 28341 -7788
rect 28405 -7852 28425 -7788
rect 22126 -7868 28425 -7852
rect 22126 -7932 28341 -7868
rect 28405 -7932 28425 -7868
rect 22126 -7948 28425 -7932
rect 22126 -8012 28341 -7948
rect 28405 -8012 28425 -7948
rect 22126 -8028 28425 -8012
rect 22126 -8092 28341 -8028
rect 28405 -8092 28425 -8028
rect 22126 -8108 28425 -8092
rect 22126 -8172 28341 -8108
rect 28405 -8172 28425 -8108
rect 22126 -8188 28425 -8172
rect 22126 -8252 28341 -8188
rect 28405 -8252 28425 -8188
rect 22126 -8268 28425 -8252
rect 22126 -8332 28341 -8268
rect 28405 -8332 28425 -8268
rect 22126 -8348 28425 -8332
rect 22126 -8412 28341 -8348
rect 28405 -8412 28425 -8348
rect 22126 -8428 28425 -8412
rect 22126 -8492 28341 -8428
rect 28405 -8492 28425 -8428
rect 22126 -8508 28425 -8492
rect 22126 -8572 28341 -8508
rect 28405 -8572 28425 -8508
rect 22126 -8588 28425 -8572
rect 22126 -8652 28341 -8588
rect 28405 -8652 28425 -8588
rect 22126 -8668 28425 -8652
rect 22126 -8732 28341 -8668
rect 28405 -8732 28425 -8668
rect 22126 -8748 28425 -8732
rect 22126 -8812 28341 -8748
rect 28405 -8812 28425 -8748
rect 22126 -8828 28425 -8812
rect 22126 -8892 28341 -8828
rect 28405 -8892 28425 -8828
rect 22126 -8908 28425 -8892
rect 22126 -8972 28341 -8908
rect 28405 -8972 28425 -8908
rect 22126 -8988 28425 -8972
rect 22126 -9052 28341 -8988
rect 28405 -9052 28425 -8988
rect 22126 -9068 28425 -9052
rect 22126 -9132 28341 -9068
rect 28405 -9132 28425 -9068
rect 22126 -9148 28425 -9132
rect 22126 -9212 28341 -9148
rect 28405 -9212 28425 -9148
rect 22126 -9228 28425 -9212
rect 22126 -9292 28341 -9228
rect 28405 -9292 28425 -9228
rect 22126 -9308 28425 -9292
rect 22126 -9372 28341 -9308
rect 28405 -9372 28425 -9308
rect 22126 -9400 28425 -9372
rect 28445 -3228 34744 -3200
rect 28445 -3292 34660 -3228
rect 34724 -3292 34744 -3228
rect 28445 -3308 34744 -3292
rect 28445 -3372 34660 -3308
rect 34724 -3372 34744 -3308
rect 28445 -3388 34744 -3372
rect 28445 -3452 34660 -3388
rect 34724 -3452 34744 -3388
rect 28445 -3468 34744 -3452
rect 28445 -3532 34660 -3468
rect 34724 -3532 34744 -3468
rect 28445 -3548 34744 -3532
rect 28445 -3612 34660 -3548
rect 34724 -3612 34744 -3548
rect 28445 -3628 34744 -3612
rect 28445 -3692 34660 -3628
rect 34724 -3692 34744 -3628
rect 28445 -3708 34744 -3692
rect 28445 -3772 34660 -3708
rect 34724 -3772 34744 -3708
rect 28445 -3788 34744 -3772
rect 28445 -3852 34660 -3788
rect 34724 -3852 34744 -3788
rect 28445 -3868 34744 -3852
rect 28445 -3932 34660 -3868
rect 34724 -3932 34744 -3868
rect 28445 -3948 34744 -3932
rect 28445 -4012 34660 -3948
rect 34724 -4012 34744 -3948
rect 28445 -4028 34744 -4012
rect 28445 -4092 34660 -4028
rect 34724 -4092 34744 -4028
rect 28445 -4108 34744 -4092
rect 28445 -4172 34660 -4108
rect 34724 -4172 34744 -4108
rect 28445 -4188 34744 -4172
rect 28445 -4252 34660 -4188
rect 34724 -4252 34744 -4188
rect 28445 -4268 34744 -4252
rect 28445 -4332 34660 -4268
rect 34724 -4332 34744 -4268
rect 28445 -4348 34744 -4332
rect 28445 -4412 34660 -4348
rect 34724 -4412 34744 -4348
rect 28445 -4428 34744 -4412
rect 28445 -4492 34660 -4428
rect 34724 -4492 34744 -4428
rect 28445 -4508 34744 -4492
rect 28445 -4572 34660 -4508
rect 34724 -4572 34744 -4508
rect 28445 -4588 34744 -4572
rect 28445 -4652 34660 -4588
rect 34724 -4652 34744 -4588
rect 28445 -4668 34744 -4652
rect 28445 -4732 34660 -4668
rect 34724 -4732 34744 -4668
rect 28445 -4748 34744 -4732
rect 28445 -4812 34660 -4748
rect 34724 -4812 34744 -4748
rect 28445 -4828 34744 -4812
rect 28445 -4892 34660 -4828
rect 34724 -4892 34744 -4828
rect 28445 -4908 34744 -4892
rect 28445 -4972 34660 -4908
rect 34724 -4972 34744 -4908
rect 28445 -4988 34744 -4972
rect 28445 -5052 34660 -4988
rect 34724 -5052 34744 -4988
rect 28445 -5068 34744 -5052
rect 28445 -5132 34660 -5068
rect 34724 -5132 34744 -5068
rect 28445 -5148 34744 -5132
rect 28445 -5212 34660 -5148
rect 34724 -5212 34744 -5148
rect 28445 -5228 34744 -5212
rect 28445 -5292 34660 -5228
rect 34724 -5292 34744 -5228
rect 28445 -5308 34744 -5292
rect 28445 -5372 34660 -5308
rect 34724 -5372 34744 -5308
rect 28445 -5388 34744 -5372
rect 28445 -5452 34660 -5388
rect 34724 -5452 34744 -5388
rect 28445 -5468 34744 -5452
rect 28445 -5532 34660 -5468
rect 34724 -5532 34744 -5468
rect 28445 -5548 34744 -5532
rect 28445 -5612 34660 -5548
rect 34724 -5612 34744 -5548
rect 28445 -5628 34744 -5612
rect 28445 -5692 34660 -5628
rect 34724 -5692 34744 -5628
rect 28445 -5708 34744 -5692
rect 28445 -5772 34660 -5708
rect 34724 -5772 34744 -5708
rect 28445 -5788 34744 -5772
rect 28445 -5852 34660 -5788
rect 34724 -5852 34744 -5788
rect 28445 -5868 34744 -5852
rect 28445 -5932 34660 -5868
rect 34724 -5932 34744 -5868
rect 28445 -5948 34744 -5932
rect 28445 -6012 34660 -5948
rect 34724 -6012 34744 -5948
rect 28445 -6028 34744 -6012
rect 28445 -6092 34660 -6028
rect 34724 -6092 34744 -6028
rect 28445 -6108 34744 -6092
rect 28445 -6172 34660 -6108
rect 34724 -6172 34744 -6108
rect 28445 -6188 34744 -6172
rect 28445 -6252 34660 -6188
rect 34724 -6252 34744 -6188
rect 28445 -6268 34744 -6252
rect 28445 -6332 34660 -6268
rect 34724 -6332 34744 -6268
rect 28445 -6348 34744 -6332
rect 28445 -6412 34660 -6348
rect 34724 -6412 34744 -6348
rect 28445 -6428 34744 -6412
rect 28445 -6492 34660 -6428
rect 34724 -6492 34744 -6428
rect 28445 -6508 34744 -6492
rect 28445 -6572 34660 -6508
rect 34724 -6572 34744 -6508
rect 28445 -6588 34744 -6572
rect 28445 -6652 34660 -6588
rect 34724 -6652 34744 -6588
rect 28445 -6668 34744 -6652
rect 28445 -6732 34660 -6668
rect 34724 -6732 34744 -6668
rect 28445 -6748 34744 -6732
rect 28445 -6812 34660 -6748
rect 34724 -6812 34744 -6748
rect 28445 -6828 34744 -6812
rect 28445 -6892 34660 -6828
rect 34724 -6892 34744 -6828
rect 28445 -6908 34744 -6892
rect 28445 -6972 34660 -6908
rect 34724 -6972 34744 -6908
rect 28445 -6988 34744 -6972
rect 28445 -7052 34660 -6988
rect 34724 -7052 34744 -6988
rect 28445 -7068 34744 -7052
rect 28445 -7132 34660 -7068
rect 34724 -7132 34744 -7068
rect 28445 -7148 34744 -7132
rect 28445 -7212 34660 -7148
rect 34724 -7212 34744 -7148
rect 28445 -7228 34744 -7212
rect 28445 -7292 34660 -7228
rect 34724 -7292 34744 -7228
rect 28445 -7308 34744 -7292
rect 28445 -7372 34660 -7308
rect 34724 -7372 34744 -7308
rect 28445 -7388 34744 -7372
rect 28445 -7452 34660 -7388
rect 34724 -7452 34744 -7388
rect 28445 -7468 34744 -7452
rect 28445 -7532 34660 -7468
rect 34724 -7532 34744 -7468
rect 28445 -7548 34744 -7532
rect 28445 -7612 34660 -7548
rect 34724 -7612 34744 -7548
rect 28445 -7628 34744 -7612
rect 28445 -7692 34660 -7628
rect 34724 -7692 34744 -7628
rect 28445 -7708 34744 -7692
rect 28445 -7772 34660 -7708
rect 34724 -7772 34744 -7708
rect 28445 -7788 34744 -7772
rect 28445 -7852 34660 -7788
rect 34724 -7852 34744 -7788
rect 28445 -7868 34744 -7852
rect 28445 -7932 34660 -7868
rect 34724 -7932 34744 -7868
rect 28445 -7948 34744 -7932
rect 28445 -8012 34660 -7948
rect 34724 -8012 34744 -7948
rect 28445 -8028 34744 -8012
rect 28445 -8092 34660 -8028
rect 34724 -8092 34744 -8028
rect 28445 -8108 34744 -8092
rect 28445 -8172 34660 -8108
rect 34724 -8172 34744 -8108
rect 28445 -8188 34744 -8172
rect 28445 -8252 34660 -8188
rect 34724 -8252 34744 -8188
rect 28445 -8268 34744 -8252
rect 28445 -8332 34660 -8268
rect 34724 -8332 34744 -8268
rect 28445 -8348 34744 -8332
rect 28445 -8412 34660 -8348
rect 34724 -8412 34744 -8348
rect 28445 -8428 34744 -8412
rect 28445 -8492 34660 -8428
rect 34724 -8492 34744 -8428
rect 28445 -8508 34744 -8492
rect 28445 -8572 34660 -8508
rect 34724 -8572 34744 -8508
rect 28445 -8588 34744 -8572
rect 28445 -8652 34660 -8588
rect 34724 -8652 34744 -8588
rect 28445 -8668 34744 -8652
rect 28445 -8732 34660 -8668
rect 34724 -8732 34744 -8668
rect 28445 -8748 34744 -8732
rect 28445 -8812 34660 -8748
rect 34724 -8812 34744 -8748
rect 28445 -8828 34744 -8812
rect 28445 -8892 34660 -8828
rect 34724 -8892 34744 -8828
rect 28445 -8908 34744 -8892
rect 28445 -8972 34660 -8908
rect 34724 -8972 34744 -8908
rect 28445 -8988 34744 -8972
rect 28445 -9052 34660 -8988
rect 34724 -9052 34744 -8988
rect 28445 -9068 34744 -9052
rect 28445 -9132 34660 -9068
rect 34724 -9132 34744 -9068
rect 28445 -9148 34744 -9132
rect 28445 -9212 34660 -9148
rect 34724 -9212 34744 -9148
rect 28445 -9228 34744 -9212
rect 28445 -9292 34660 -9228
rect 34724 -9292 34744 -9228
rect 28445 -9308 34744 -9292
rect 28445 -9372 34660 -9308
rect 34724 -9372 34744 -9308
rect 28445 -9400 34744 -9372
rect 34764 -3228 41063 -3200
rect 34764 -3292 40979 -3228
rect 41043 -3292 41063 -3228
rect 34764 -3308 41063 -3292
rect 34764 -3372 40979 -3308
rect 41043 -3372 41063 -3308
rect 34764 -3388 41063 -3372
rect 34764 -3452 40979 -3388
rect 41043 -3452 41063 -3388
rect 34764 -3468 41063 -3452
rect 34764 -3532 40979 -3468
rect 41043 -3532 41063 -3468
rect 34764 -3548 41063 -3532
rect 34764 -3612 40979 -3548
rect 41043 -3612 41063 -3548
rect 34764 -3628 41063 -3612
rect 34764 -3692 40979 -3628
rect 41043 -3692 41063 -3628
rect 34764 -3708 41063 -3692
rect 34764 -3772 40979 -3708
rect 41043 -3772 41063 -3708
rect 34764 -3788 41063 -3772
rect 34764 -3852 40979 -3788
rect 41043 -3852 41063 -3788
rect 34764 -3868 41063 -3852
rect 34764 -3932 40979 -3868
rect 41043 -3932 41063 -3868
rect 34764 -3948 41063 -3932
rect 34764 -4012 40979 -3948
rect 41043 -4012 41063 -3948
rect 34764 -4028 41063 -4012
rect 34764 -4092 40979 -4028
rect 41043 -4092 41063 -4028
rect 34764 -4108 41063 -4092
rect 34764 -4172 40979 -4108
rect 41043 -4172 41063 -4108
rect 34764 -4188 41063 -4172
rect 34764 -4252 40979 -4188
rect 41043 -4252 41063 -4188
rect 34764 -4268 41063 -4252
rect 34764 -4332 40979 -4268
rect 41043 -4332 41063 -4268
rect 34764 -4348 41063 -4332
rect 34764 -4412 40979 -4348
rect 41043 -4412 41063 -4348
rect 34764 -4428 41063 -4412
rect 34764 -4492 40979 -4428
rect 41043 -4492 41063 -4428
rect 34764 -4508 41063 -4492
rect 34764 -4572 40979 -4508
rect 41043 -4572 41063 -4508
rect 34764 -4588 41063 -4572
rect 34764 -4652 40979 -4588
rect 41043 -4652 41063 -4588
rect 34764 -4668 41063 -4652
rect 34764 -4732 40979 -4668
rect 41043 -4732 41063 -4668
rect 34764 -4748 41063 -4732
rect 34764 -4812 40979 -4748
rect 41043 -4812 41063 -4748
rect 34764 -4828 41063 -4812
rect 34764 -4892 40979 -4828
rect 41043 -4892 41063 -4828
rect 34764 -4908 41063 -4892
rect 34764 -4972 40979 -4908
rect 41043 -4972 41063 -4908
rect 34764 -4988 41063 -4972
rect 34764 -5052 40979 -4988
rect 41043 -5052 41063 -4988
rect 34764 -5068 41063 -5052
rect 34764 -5132 40979 -5068
rect 41043 -5132 41063 -5068
rect 34764 -5148 41063 -5132
rect 34764 -5212 40979 -5148
rect 41043 -5212 41063 -5148
rect 34764 -5228 41063 -5212
rect 34764 -5292 40979 -5228
rect 41043 -5292 41063 -5228
rect 34764 -5308 41063 -5292
rect 34764 -5372 40979 -5308
rect 41043 -5372 41063 -5308
rect 34764 -5388 41063 -5372
rect 34764 -5452 40979 -5388
rect 41043 -5452 41063 -5388
rect 34764 -5468 41063 -5452
rect 34764 -5532 40979 -5468
rect 41043 -5532 41063 -5468
rect 34764 -5548 41063 -5532
rect 34764 -5612 40979 -5548
rect 41043 -5612 41063 -5548
rect 34764 -5628 41063 -5612
rect 34764 -5692 40979 -5628
rect 41043 -5692 41063 -5628
rect 34764 -5708 41063 -5692
rect 34764 -5772 40979 -5708
rect 41043 -5772 41063 -5708
rect 34764 -5788 41063 -5772
rect 34764 -5852 40979 -5788
rect 41043 -5852 41063 -5788
rect 34764 -5868 41063 -5852
rect 34764 -5932 40979 -5868
rect 41043 -5932 41063 -5868
rect 34764 -5948 41063 -5932
rect 34764 -6012 40979 -5948
rect 41043 -6012 41063 -5948
rect 34764 -6028 41063 -6012
rect 34764 -6092 40979 -6028
rect 41043 -6092 41063 -6028
rect 34764 -6108 41063 -6092
rect 34764 -6172 40979 -6108
rect 41043 -6172 41063 -6108
rect 34764 -6188 41063 -6172
rect 34764 -6252 40979 -6188
rect 41043 -6252 41063 -6188
rect 34764 -6268 41063 -6252
rect 34764 -6332 40979 -6268
rect 41043 -6332 41063 -6268
rect 34764 -6348 41063 -6332
rect 34764 -6412 40979 -6348
rect 41043 -6412 41063 -6348
rect 34764 -6428 41063 -6412
rect 34764 -6492 40979 -6428
rect 41043 -6492 41063 -6428
rect 34764 -6508 41063 -6492
rect 34764 -6572 40979 -6508
rect 41043 -6572 41063 -6508
rect 34764 -6588 41063 -6572
rect 34764 -6652 40979 -6588
rect 41043 -6652 41063 -6588
rect 34764 -6668 41063 -6652
rect 34764 -6732 40979 -6668
rect 41043 -6732 41063 -6668
rect 34764 -6748 41063 -6732
rect 34764 -6812 40979 -6748
rect 41043 -6812 41063 -6748
rect 34764 -6828 41063 -6812
rect 34764 -6892 40979 -6828
rect 41043 -6892 41063 -6828
rect 34764 -6908 41063 -6892
rect 34764 -6972 40979 -6908
rect 41043 -6972 41063 -6908
rect 34764 -6988 41063 -6972
rect 34764 -7052 40979 -6988
rect 41043 -7052 41063 -6988
rect 34764 -7068 41063 -7052
rect 34764 -7132 40979 -7068
rect 41043 -7132 41063 -7068
rect 34764 -7148 41063 -7132
rect 34764 -7212 40979 -7148
rect 41043 -7212 41063 -7148
rect 34764 -7228 41063 -7212
rect 34764 -7292 40979 -7228
rect 41043 -7292 41063 -7228
rect 34764 -7308 41063 -7292
rect 34764 -7372 40979 -7308
rect 41043 -7372 41063 -7308
rect 34764 -7388 41063 -7372
rect 34764 -7452 40979 -7388
rect 41043 -7452 41063 -7388
rect 34764 -7468 41063 -7452
rect 34764 -7532 40979 -7468
rect 41043 -7532 41063 -7468
rect 34764 -7548 41063 -7532
rect 34764 -7612 40979 -7548
rect 41043 -7612 41063 -7548
rect 34764 -7628 41063 -7612
rect 34764 -7692 40979 -7628
rect 41043 -7692 41063 -7628
rect 34764 -7708 41063 -7692
rect 34764 -7772 40979 -7708
rect 41043 -7772 41063 -7708
rect 34764 -7788 41063 -7772
rect 34764 -7852 40979 -7788
rect 41043 -7852 41063 -7788
rect 34764 -7868 41063 -7852
rect 34764 -7932 40979 -7868
rect 41043 -7932 41063 -7868
rect 34764 -7948 41063 -7932
rect 34764 -8012 40979 -7948
rect 41043 -8012 41063 -7948
rect 34764 -8028 41063 -8012
rect 34764 -8092 40979 -8028
rect 41043 -8092 41063 -8028
rect 34764 -8108 41063 -8092
rect 34764 -8172 40979 -8108
rect 41043 -8172 41063 -8108
rect 34764 -8188 41063 -8172
rect 34764 -8252 40979 -8188
rect 41043 -8252 41063 -8188
rect 34764 -8268 41063 -8252
rect 34764 -8332 40979 -8268
rect 41043 -8332 41063 -8268
rect 34764 -8348 41063 -8332
rect 34764 -8412 40979 -8348
rect 41043 -8412 41063 -8348
rect 34764 -8428 41063 -8412
rect 34764 -8492 40979 -8428
rect 41043 -8492 41063 -8428
rect 34764 -8508 41063 -8492
rect 34764 -8572 40979 -8508
rect 41043 -8572 41063 -8508
rect 34764 -8588 41063 -8572
rect 34764 -8652 40979 -8588
rect 41043 -8652 41063 -8588
rect 34764 -8668 41063 -8652
rect 34764 -8732 40979 -8668
rect 41043 -8732 41063 -8668
rect 34764 -8748 41063 -8732
rect 34764 -8812 40979 -8748
rect 41043 -8812 41063 -8748
rect 34764 -8828 41063 -8812
rect 34764 -8892 40979 -8828
rect 41043 -8892 41063 -8828
rect 34764 -8908 41063 -8892
rect 34764 -8972 40979 -8908
rect 41043 -8972 41063 -8908
rect 34764 -8988 41063 -8972
rect 34764 -9052 40979 -8988
rect 41043 -9052 41063 -8988
rect 34764 -9068 41063 -9052
rect 34764 -9132 40979 -9068
rect 41043 -9132 41063 -9068
rect 34764 -9148 41063 -9132
rect 34764 -9212 40979 -9148
rect 41043 -9212 41063 -9148
rect 34764 -9228 41063 -9212
rect 34764 -9292 40979 -9228
rect 41043 -9292 41063 -9228
rect 34764 -9308 41063 -9292
rect 34764 -9372 40979 -9308
rect 41043 -9372 41063 -9308
rect 34764 -9400 41063 -9372
rect 41083 -3228 47382 -3200
rect 41083 -3292 47298 -3228
rect 47362 -3292 47382 -3228
rect 41083 -3308 47382 -3292
rect 41083 -3372 47298 -3308
rect 47362 -3372 47382 -3308
rect 41083 -3388 47382 -3372
rect 41083 -3452 47298 -3388
rect 47362 -3452 47382 -3388
rect 41083 -3468 47382 -3452
rect 41083 -3532 47298 -3468
rect 47362 -3532 47382 -3468
rect 41083 -3548 47382 -3532
rect 41083 -3612 47298 -3548
rect 47362 -3612 47382 -3548
rect 41083 -3628 47382 -3612
rect 41083 -3692 47298 -3628
rect 47362 -3692 47382 -3628
rect 41083 -3708 47382 -3692
rect 41083 -3772 47298 -3708
rect 47362 -3772 47382 -3708
rect 41083 -3788 47382 -3772
rect 41083 -3852 47298 -3788
rect 47362 -3852 47382 -3788
rect 41083 -3868 47382 -3852
rect 41083 -3932 47298 -3868
rect 47362 -3932 47382 -3868
rect 41083 -3948 47382 -3932
rect 41083 -4012 47298 -3948
rect 47362 -4012 47382 -3948
rect 41083 -4028 47382 -4012
rect 41083 -4092 47298 -4028
rect 47362 -4092 47382 -4028
rect 41083 -4108 47382 -4092
rect 41083 -4172 47298 -4108
rect 47362 -4172 47382 -4108
rect 41083 -4188 47382 -4172
rect 41083 -4252 47298 -4188
rect 47362 -4252 47382 -4188
rect 41083 -4268 47382 -4252
rect 41083 -4332 47298 -4268
rect 47362 -4332 47382 -4268
rect 41083 -4348 47382 -4332
rect 41083 -4412 47298 -4348
rect 47362 -4412 47382 -4348
rect 41083 -4428 47382 -4412
rect 41083 -4492 47298 -4428
rect 47362 -4492 47382 -4428
rect 41083 -4508 47382 -4492
rect 41083 -4572 47298 -4508
rect 47362 -4572 47382 -4508
rect 41083 -4588 47382 -4572
rect 41083 -4652 47298 -4588
rect 47362 -4652 47382 -4588
rect 41083 -4668 47382 -4652
rect 41083 -4732 47298 -4668
rect 47362 -4732 47382 -4668
rect 41083 -4748 47382 -4732
rect 41083 -4812 47298 -4748
rect 47362 -4812 47382 -4748
rect 41083 -4828 47382 -4812
rect 41083 -4892 47298 -4828
rect 47362 -4892 47382 -4828
rect 41083 -4908 47382 -4892
rect 41083 -4972 47298 -4908
rect 47362 -4972 47382 -4908
rect 41083 -4988 47382 -4972
rect 41083 -5052 47298 -4988
rect 47362 -5052 47382 -4988
rect 41083 -5068 47382 -5052
rect 41083 -5132 47298 -5068
rect 47362 -5132 47382 -5068
rect 41083 -5148 47382 -5132
rect 41083 -5212 47298 -5148
rect 47362 -5212 47382 -5148
rect 41083 -5228 47382 -5212
rect 41083 -5292 47298 -5228
rect 47362 -5292 47382 -5228
rect 41083 -5308 47382 -5292
rect 41083 -5372 47298 -5308
rect 47362 -5372 47382 -5308
rect 41083 -5388 47382 -5372
rect 41083 -5452 47298 -5388
rect 47362 -5452 47382 -5388
rect 41083 -5468 47382 -5452
rect 41083 -5532 47298 -5468
rect 47362 -5532 47382 -5468
rect 41083 -5548 47382 -5532
rect 41083 -5612 47298 -5548
rect 47362 -5612 47382 -5548
rect 41083 -5628 47382 -5612
rect 41083 -5692 47298 -5628
rect 47362 -5692 47382 -5628
rect 41083 -5708 47382 -5692
rect 41083 -5772 47298 -5708
rect 47362 -5772 47382 -5708
rect 41083 -5788 47382 -5772
rect 41083 -5852 47298 -5788
rect 47362 -5852 47382 -5788
rect 41083 -5868 47382 -5852
rect 41083 -5932 47298 -5868
rect 47362 -5932 47382 -5868
rect 41083 -5948 47382 -5932
rect 41083 -6012 47298 -5948
rect 47362 -6012 47382 -5948
rect 41083 -6028 47382 -6012
rect 41083 -6092 47298 -6028
rect 47362 -6092 47382 -6028
rect 41083 -6108 47382 -6092
rect 41083 -6172 47298 -6108
rect 47362 -6172 47382 -6108
rect 41083 -6188 47382 -6172
rect 41083 -6252 47298 -6188
rect 47362 -6252 47382 -6188
rect 41083 -6268 47382 -6252
rect 41083 -6332 47298 -6268
rect 47362 -6332 47382 -6268
rect 41083 -6348 47382 -6332
rect 41083 -6412 47298 -6348
rect 47362 -6412 47382 -6348
rect 41083 -6428 47382 -6412
rect 41083 -6492 47298 -6428
rect 47362 -6492 47382 -6428
rect 41083 -6508 47382 -6492
rect 41083 -6572 47298 -6508
rect 47362 -6572 47382 -6508
rect 41083 -6588 47382 -6572
rect 41083 -6652 47298 -6588
rect 47362 -6652 47382 -6588
rect 41083 -6668 47382 -6652
rect 41083 -6732 47298 -6668
rect 47362 -6732 47382 -6668
rect 41083 -6748 47382 -6732
rect 41083 -6812 47298 -6748
rect 47362 -6812 47382 -6748
rect 41083 -6828 47382 -6812
rect 41083 -6892 47298 -6828
rect 47362 -6892 47382 -6828
rect 41083 -6908 47382 -6892
rect 41083 -6972 47298 -6908
rect 47362 -6972 47382 -6908
rect 41083 -6988 47382 -6972
rect 41083 -7052 47298 -6988
rect 47362 -7052 47382 -6988
rect 41083 -7068 47382 -7052
rect 41083 -7132 47298 -7068
rect 47362 -7132 47382 -7068
rect 41083 -7148 47382 -7132
rect 41083 -7212 47298 -7148
rect 47362 -7212 47382 -7148
rect 41083 -7228 47382 -7212
rect 41083 -7292 47298 -7228
rect 47362 -7292 47382 -7228
rect 41083 -7308 47382 -7292
rect 41083 -7372 47298 -7308
rect 47362 -7372 47382 -7308
rect 41083 -7388 47382 -7372
rect 41083 -7452 47298 -7388
rect 47362 -7452 47382 -7388
rect 41083 -7468 47382 -7452
rect 41083 -7532 47298 -7468
rect 47362 -7532 47382 -7468
rect 41083 -7548 47382 -7532
rect 41083 -7612 47298 -7548
rect 47362 -7612 47382 -7548
rect 41083 -7628 47382 -7612
rect 41083 -7692 47298 -7628
rect 47362 -7692 47382 -7628
rect 41083 -7708 47382 -7692
rect 41083 -7772 47298 -7708
rect 47362 -7772 47382 -7708
rect 41083 -7788 47382 -7772
rect 41083 -7852 47298 -7788
rect 47362 -7852 47382 -7788
rect 41083 -7868 47382 -7852
rect 41083 -7932 47298 -7868
rect 47362 -7932 47382 -7868
rect 41083 -7948 47382 -7932
rect 41083 -8012 47298 -7948
rect 47362 -8012 47382 -7948
rect 41083 -8028 47382 -8012
rect 41083 -8092 47298 -8028
rect 47362 -8092 47382 -8028
rect 41083 -8108 47382 -8092
rect 41083 -8172 47298 -8108
rect 47362 -8172 47382 -8108
rect 41083 -8188 47382 -8172
rect 41083 -8252 47298 -8188
rect 47362 -8252 47382 -8188
rect 41083 -8268 47382 -8252
rect 41083 -8332 47298 -8268
rect 47362 -8332 47382 -8268
rect 41083 -8348 47382 -8332
rect 41083 -8412 47298 -8348
rect 47362 -8412 47382 -8348
rect 41083 -8428 47382 -8412
rect 41083 -8492 47298 -8428
rect 47362 -8492 47382 -8428
rect 41083 -8508 47382 -8492
rect 41083 -8572 47298 -8508
rect 47362 -8572 47382 -8508
rect 41083 -8588 47382 -8572
rect 41083 -8652 47298 -8588
rect 47362 -8652 47382 -8588
rect 41083 -8668 47382 -8652
rect 41083 -8732 47298 -8668
rect 47362 -8732 47382 -8668
rect 41083 -8748 47382 -8732
rect 41083 -8812 47298 -8748
rect 47362 -8812 47382 -8748
rect 41083 -8828 47382 -8812
rect 41083 -8892 47298 -8828
rect 47362 -8892 47382 -8828
rect 41083 -8908 47382 -8892
rect 41083 -8972 47298 -8908
rect 47362 -8972 47382 -8908
rect 41083 -8988 47382 -8972
rect 41083 -9052 47298 -8988
rect 47362 -9052 47382 -8988
rect 41083 -9068 47382 -9052
rect 41083 -9132 47298 -9068
rect 47362 -9132 47382 -9068
rect 41083 -9148 47382 -9132
rect 41083 -9212 47298 -9148
rect 47362 -9212 47382 -9148
rect 41083 -9228 47382 -9212
rect 41083 -9292 47298 -9228
rect 47362 -9292 47382 -9228
rect 41083 -9308 47382 -9292
rect 41083 -9372 47298 -9308
rect 47362 -9372 47382 -9308
rect 41083 -9400 47382 -9372
rect -47383 -9528 -41084 -9500
rect -47383 -9592 -41168 -9528
rect -41104 -9592 -41084 -9528
rect -47383 -9608 -41084 -9592
rect -47383 -9672 -41168 -9608
rect -41104 -9672 -41084 -9608
rect -47383 -9688 -41084 -9672
rect -47383 -9752 -41168 -9688
rect -41104 -9752 -41084 -9688
rect -47383 -9768 -41084 -9752
rect -47383 -9832 -41168 -9768
rect -41104 -9832 -41084 -9768
rect -47383 -9848 -41084 -9832
rect -47383 -9912 -41168 -9848
rect -41104 -9912 -41084 -9848
rect -47383 -9928 -41084 -9912
rect -47383 -9992 -41168 -9928
rect -41104 -9992 -41084 -9928
rect -47383 -10008 -41084 -9992
rect -47383 -10072 -41168 -10008
rect -41104 -10072 -41084 -10008
rect -47383 -10088 -41084 -10072
rect -47383 -10152 -41168 -10088
rect -41104 -10152 -41084 -10088
rect -47383 -10168 -41084 -10152
rect -47383 -10232 -41168 -10168
rect -41104 -10232 -41084 -10168
rect -47383 -10248 -41084 -10232
rect -47383 -10312 -41168 -10248
rect -41104 -10312 -41084 -10248
rect -47383 -10328 -41084 -10312
rect -47383 -10392 -41168 -10328
rect -41104 -10392 -41084 -10328
rect -47383 -10408 -41084 -10392
rect -47383 -10472 -41168 -10408
rect -41104 -10472 -41084 -10408
rect -47383 -10488 -41084 -10472
rect -47383 -10552 -41168 -10488
rect -41104 -10552 -41084 -10488
rect -47383 -10568 -41084 -10552
rect -47383 -10632 -41168 -10568
rect -41104 -10632 -41084 -10568
rect -47383 -10648 -41084 -10632
rect -47383 -10712 -41168 -10648
rect -41104 -10712 -41084 -10648
rect -47383 -10728 -41084 -10712
rect -47383 -10792 -41168 -10728
rect -41104 -10792 -41084 -10728
rect -47383 -10808 -41084 -10792
rect -47383 -10872 -41168 -10808
rect -41104 -10872 -41084 -10808
rect -47383 -10888 -41084 -10872
rect -47383 -10952 -41168 -10888
rect -41104 -10952 -41084 -10888
rect -47383 -10968 -41084 -10952
rect -47383 -11032 -41168 -10968
rect -41104 -11032 -41084 -10968
rect -47383 -11048 -41084 -11032
rect -47383 -11112 -41168 -11048
rect -41104 -11112 -41084 -11048
rect -47383 -11128 -41084 -11112
rect -47383 -11192 -41168 -11128
rect -41104 -11192 -41084 -11128
rect -47383 -11208 -41084 -11192
rect -47383 -11272 -41168 -11208
rect -41104 -11272 -41084 -11208
rect -47383 -11288 -41084 -11272
rect -47383 -11352 -41168 -11288
rect -41104 -11352 -41084 -11288
rect -47383 -11368 -41084 -11352
rect -47383 -11432 -41168 -11368
rect -41104 -11432 -41084 -11368
rect -47383 -11448 -41084 -11432
rect -47383 -11512 -41168 -11448
rect -41104 -11512 -41084 -11448
rect -47383 -11528 -41084 -11512
rect -47383 -11592 -41168 -11528
rect -41104 -11592 -41084 -11528
rect -47383 -11608 -41084 -11592
rect -47383 -11672 -41168 -11608
rect -41104 -11672 -41084 -11608
rect -47383 -11688 -41084 -11672
rect -47383 -11752 -41168 -11688
rect -41104 -11752 -41084 -11688
rect -47383 -11768 -41084 -11752
rect -47383 -11832 -41168 -11768
rect -41104 -11832 -41084 -11768
rect -47383 -11848 -41084 -11832
rect -47383 -11912 -41168 -11848
rect -41104 -11912 -41084 -11848
rect -47383 -11928 -41084 -11912
rect -47383 -11992 -41168 -11928
rect -41104 -11992 -41084 -11928
rect -47383 -12008 -41084 -11992
rect -47383 -12072 -41168 -12008
rect -41104 -12072 -41084 -12008
rect -47383 -12088 -41084 -12072
rect -47383 -12152 -41168 -12088
rect -41104 -12152 -41084 -12088
rect -47383 -12168 -41084 -12152
rect -47383 -12232 -41168 -12168
rect -41104 -12232 -41084 -12168
rect -47383 -12248 -41084 -12232
rect -47383 -12312 -41168 -12248
rect -41104 -12312 -41084 -12248
rect -47383 -12328 -41084 -12312
rect -47383 -12392 -41168 -12328
rect -41104 -12392 -41084 -12328
rect -47383 -12408 -41084 -12392
rect -47383 -12472 -41168 -12408
rect -41104 -12472 -41084 -12408
rect -47383 -12488 -41084 -12472
rect -47383 -12552 -41168 -12488
rect -41104 -12552 -41084 -12488
rect -47383 -12568 -41084 -12552
rect -47383 -12632 -41168 -12568
rect -41104 -12632 -41084 -12568
rect -47383 -12648 -41084 -12632
rect -47383 -12712 -41168 -12648
rect -41104 -12712 -41084 -12648
rect -47383 -12728 -41084 -12712
rect -47383 -12792 -41168 -12728
rect -41104 -12792 -41084 -12728
rect -47383 -12808 -41084 -12792
rect -47383 -12872 -41168 -12808
rect -41104 -12872 -41084 -12808
rect -47383 -12888 -41084 -12872
rect -47383 -12952 -41168 -12888
rect -41104 -12952 -41084 -12888
rect -47383 -12968 -41084 -12952
rect -47383 -13032 -41168 -12968
rect -41104 -13032 -41084 -12968
rect -47383 -13048 -41084 -13032
rect -47383 -13112 -41168 -13048
rect -41104 -13112 -41084 -13048
rect -47383 -13128 -41084 -13112
rect -47383 -13192 -41168 -13128
rect -41104 -13192 -41084 -13128
rect -47383 -13208 -41084 -13192
rect -47383 -13272 -41168 -13208
rect -41104 -13272 -41084 -13208
rect -47383 -13288 -41084 -13272
rect -47383 -13352 -41168 -13288
rect -41104 -13352 -41084 -13288
rect -47383 -13368 -41084 -13352
rect -47383 -13432 -41168 -13368
rect -41104 -13432 -41084 -13368
rect -47383 -13448 -41084 -13432
rect -47383 -13512 -41168 -13448
rect -41104 -13512 -41084 -13448
rect -47383 -13528 -41084 -13512
rect -47383 -13592 -41168 -13528
rect -41104 -13592 -41084 -13528
rect -47383 -13608 -41084 -13592
rect -47383 -13672 -41168 -13608
rect -41104 -13672 -41084 -13608
rect -47383 -13688 -41084 -13672
rect -47383 -13752 -41168 -13688
rect -41104 -13752 -41084 -13688
rect -47383 -13768 -41084 -13752
rect -47383 -13832 -41168 -13768
rect -41104 -13832 -41084 -13768
rect -47383 -13848 -41084 -13832
rect -47383 -13912 -41168 -13848
rect -41104 -13912 -41084 -13848
rect -47383 -13928 -41084 -13912
rect -47383 -13992 -41168 -13928
rect -41104 -13992 -41084 -13928
rect -47383 -14008 -41084 -13992
rect -47383 -14072 -41168 -14008
rect -41104 -14072 -41084 -14008
rect -47383 -14088 -41084 -14072
rect -47383 -14152 -41168 -14088
rect -41104 -14152 -41084 -14088
rect -47383 -14168 -41084 -14152
rect -47383 -14232 -41168 -14168
rect -41104 -14232 -41084 -14168
rect -47383 -14248 -41084 -14232
rect -47383 -14312 -41168 -14248
rect -41104 -14312 -41084 -14248
rect -47383 -14328 -41084 -14312
rect -47383 -14392 -41168 -14328
rect -41104 -14392 -41084 -14328
rect -47383 -14408 -41084 -14392
rect -47383 -14472 -41168 -14408
rect -41104 -14472 -41084 -14408
rect -47383 -14488 -41084 -14472
rect -47383 -14552 -41168 -14488
rect -41104 -14552 -41084 -14488
rect -47383 -14568 -41084 -14552
rect -47383 -14632 -41168 -14568
rect -41104 -14632 -41084 -14568
rect -47383 -14648 -41084 -14632
rect -47383 -14712 -41168 -14648
rect -41104 -14712 -41084 -14648
rect -47383 -14728 -41084 -14712
rect -47383 -14792 -41168 -14728
rect -41104 -14792 -41084 -14728
rect -47383 -14808 -41084 -14792
rect -47383 -14872 -41168 -14808
rect -41104 -14872 -41084 -14808
rect -47383 -14888 -41084 -14872
rect -47383 -14952 -41168 -14888
rect -41104 -14952 -41084 -14888
rect -47383 -14968 -41084 -14952
rect -47383 -15032 -41168 -14968
rect -41104 -15032 -41084 -14968
rect -47383 -15048 -41084 -15032
rect -47383 -15112 -41168 -15048
rect -41104 -15112 -41084 -15048
rect -47383 -15128 -41084 -15112
rect -47383 -15192 -41168 -15128
rect -41104 -15192 -41084 -15128
rect -47383 -15208 -41084 -15192
rect -47383 -15272 -41168 -15208
rect -41104 -15272 -41084 -15208
rect -47383 -15288 -41084 -15272
rect -47383 -15352 -41168 -15288
rect -41104 -15352 -41084 -15288
rect -47383 -15368 -41084 -15352
rect -47383 -15432 -41168 -15368
rect -41104 -15432 -41084 -15368
rect -47383 -15448 -41084 -15432
rect -47383 -15512 -41168 -15448
rect -41104 -15512 -41084 -15448
rect -47383 -15528 -41084 -15512
rect -47383 -15592 -41168 -15528
rect -41104 -15592 -41084 -15528
rect -47383 -15608 -41084 -15592
rect -47383 -15672 -41168 -15608
rect -41104 -15672 -41084 -15608
rect -47383 -15700 -41084 -15672
rect -41064 -9528 -34765 -9500
rect -41064 -9592 -34849 -9528
rect -34785 -9592 -34765 -9528
rect -41064 -9608 -34765 -9592
rect -41064 -9672 -34849 -9608
rect -34785 -9672 -34765 -9608
rect -41064 -9688 -34765 -9672
rect -41064 -9752 -34849 -9688
rect -34785 -9752 -34765 -9688
rect -41064 -9768 -34765 -9752
rect -41064 -9832 -34849 -9768
rect -34785 -9832 -34765 -9768
rect -41064 -9848 -34765 -9832
rect -41064 -9912 -34849 -9848
rect -34785 -9912 -34765 -9848
rect -41064 -9928 -34765 -9912
rect -41064 -9992 -34849 -9928
rect -34785 -9992 -34765 -9928
rect -41064 -10008 -34765 -9992
rect -41064 -10072 -34849 -10008
rect -34785 -10072 -34765 -10008
rect -41064 -10088 -34765 -10072
rect -41064 -10152 -34849 -10088
rect -34785 -10152 -34765 -10088
rect -41064 -10168 -34765 -10152
rect -41064 -10232 -34849 -10168
rect -34785 -10232 -34765 -10168
rect -41064 -10248 -34765 -10232
rect -41064 -10312 -34849 -10248
rect -34785 -10312 -34765 -10248
rect -41064 -10328 -34765 -10312
rect -41064 -10392 -34849 -10328
rect -34785 -10392 -34765 -10328
rect -41064 -10408 -34765 -10392
rect -41064 -10472 -34849 -10408
rect -34785 -10472 -34765 -10408
rect -41064 -10488 -34765 -10472
rect -41064 -10552 -34849 -10488
rect -34785 -10552 -34765 -10488
rect -41064 -10568 -34765 -10552
rect -41064 -10632 -34849 -10568
rect -34785 -10632 -34765 -10568
rect -41064 -10648 -34765 -10632
rect -41064 -10712 -34849 -10648
rect -34785 -10712 -34765 -10648
rect -41064 -10728 -34765 -10712
rect -41064 -10792 -34849 -10728
rect -34785 -10792 -34765 -10728
rect -41064 -10808 -34765 -10792
rect -41064 -10872 -34849 -10808
rect -34785 -10872 -34765 -10808
rect -41064 -10888 -34765 -10872
rect -41064 -10952 -34849 -10888
rect -34785 -10952 -34765 -10888
rect -41064 -10968 -34765 -10952
rect -41064 -11032 -34849 -10968
rect -34785 -11032 -34765 -10968
rect -41064 -11048 -34765 -11032
rect -41064 -11112 -34849 -11048
rect -34785 -11112 -34765 -11048
rect -41064 -11128 -34765 -11112
rect -41064 -11192 -34849 -11128
rect -34785 -11192 -34765 -11128
rect -41064 -11208 -34765 -11192
rect -41064 -11272 -34849 -11208
rect -34785 -11272 -34765 -11208
rect -41064 -11288 -34765 -11272
rect -41064 -11352 -34849 -11288
rect -34785 -11352 -34765 -11288
rect -41064 -11368 -34765 -11352
rect -41064 -11432 -34849 -11368
rect -34785 -11432 -34765 -11368
rect -41064 -11448 -34765 -11432
rect -41064 -11512 -34849 -11448
rect -34785 -11512 -34765 -11448
rect -41064 -11528 -34765 -11512
rect -41064 -11592 -34849 -11528
rect -34785 -11592 -34765 -11528
rect -41064 -11608 -34765 -11592
rect -41064 -11672 -34849 -11608
rect -34785 -11672 -34765 -11608
rect -41064 -11688 -34765 -11672
rect -41064 -11752 -34849 -11688
rect -34785 -11752 -34765 -11688
rect -41064 -11768 -34765 -11752
rect -41064 -11832 -34849 -11768
rect -34785 -11832 -34765 -11768
rect -41064 -11848 -34765 -11832
rect -41064 -11912 -34849 -11848
rect -34785 -11912 -34765 -11848
rect -41064 -11928 -34765 -11912
rect -41064 -11992 -34849 -11928
rect -34785 -11992 -34765 -11928
rect -41064 -12008 -34765 -11992
rect -41064 -12072 -34849 -12008
rect -34785 -12072 -34765 -12008
rect -41064 -12088 -34765 -12072
rect -41064 -12152 -34849 -12088
rect -34785 -12152 -34765 -12088
rect -41064 -12168 -34765 -12152
rect -41064 -12232 -34849 -12168
rect -34785 -12232 -34765 -12168
rect -41064 -12248 -34765 -12232
rect -41064 -12312 -34849 -12248
rect -34785 -12312 -34765 -12248
rect -41064 -12328 -34765 -12312
rect -41064 -12392 -34849 -12328
rect -34785 -12392 -34765 -12328
rect -41064 -12408 -34765 -12392
rect -41064 -12472 -34849 -12408
rect -34785 -12472 -34765 -12408
rect -41064 -12488 -34765 -12472
rect -41064 -12552 -34849 -12488
rect -34785 -12552 -34765 -12488
rect -41064 -12568 -34765 -12552
rect -41064 -12632 -34849 -12568
rect -34785 -12632 -34765 -12568
rect -41064 -12648 -34765 -12632
rect -41064 -12712 -34849 -12648
rect -34785 -12712 -34765 -12648
rect -41064 -12728 -34765 -12712
rect -41064 -12792 -34849 -12728
rect -34785 -12792 -34765 -12728
rect -41064 -12808 -34765 -12792
rect -41064 -12872 -34849 -12808
rect -34785 -12872 -34765 -12808
rect -41064 -12888 -34765 -12872
rect -41064 -12952 -34849 -12888
rect -34785 -12952 -34765 -12888
rect -41064 -12968 -34765 -12952
rect -41064 -13032 -34849 -12968
rect -34785 -13032 -34765 -12968
rect -41064 -13048 -34765 -13032
rect -41064 -13112 -34849 -13048
rect -34785 -13112 -34765 -13048
rect -41064 -13128 -34765 -13112
rect -41064 -13192 -34849 -13128
rect -34785 -13192 -34765 -13128
rect -41064 -13208 -34765 -13192
rect -41064 -13272 -34849 -13208
rect -34785 -13272 -34765 -13208
rect -41064 -13288 -34765 -13272
rect -41064 -13352 -34849 -13288
rect -34785 -13352 -34765 -13288
rect -41064 -13368 -34765 -13352
rect -41064 -13432 -34849 -13368
rect -34785 -13432 -34765 -13368
rect -41064 -13448 -34765 -13432
rect -41064 -13512 -34849 -13448
rect -34785 -13512 -34765 -13448
rect -41064 -13528 -34765 -13512
rect -41064 -13592 -34849 -13528
rect -34785 -13592 -34765 -13528
rect -41064 -13608 -34765 -13592
rect -41064 -13672 -34849 -13608
rect -34785 -13672 -34765 -13608
rect -41064 -13688 -34765 -13672
rect -41064 -13752 -34849 -13688
rect -34785 -13752 -34765 -13688
rect -41064 -13768 -34765 -13752
rect -41064 -13832 -34849 -13768
rect -34785 -13832 -34765 -13768
rect -41064 -13848 -34765 -13832
rect -41064 -13912 -34849 -13848
rect -34785 -13912 -34765 -13848
rect -41064 -13928 -34765 -13912
rect -41064 -13992 -34849 -13928
rect -34785 -13992 -34765 -13928
rect -41064 -14008 -34765 -13992
rect -41064 -14072 -34849 -14008
rect -34785 -14072 -34765 -14008
rect -41064 -14088 -34765 -14072
rect -41064 -14152 -34849 -14088
rect -34785 -14152 -34765 -14088
rect -41064 -14168 -34765 -14152
rect -41064 -14232 -34849 -14168
rect -34785 -14232 -34765 -14168
rect -41064 -14248 -34765 -14232
rect -41064 -14312 -34849 -14248
rect -34785 -14312 -34765 -14248
rect -41064 -14328 -34765 -14312
rect -41064 -14392 -34849 -14328
rect -34785 -14392 -34765 -14328
rect -41064 -14408 -34765 -14392
rect -41064 -14472 -34849 -14408
rect -34785 -14472 -34765 -14408
rect -41064 -14488 -34765 -14472
rect -41064 -14552 -34849 -14488
rect -34785 -14552 -34765 -14488
rect -41064 -14568 -34765 -14552
rect -41064 -14632 -34849 -14568
rect -34785 -14632 -34765 -14568
rect -41064 -14648 -34765 -14632
rect -41064 -14712 -34849 -14648
rect -34785 -14712 -34765 -14648
rect -41064 -14728 -34765 -14712
rect -41064 -14792 -34849 -14728
rect -34785 -14792 -34765 -14728
rect -41064 -14808 -34765 -14792
rect -41064 -14872 -34849 -14808
rect -34785 -14872 -34765 -14808
rect -41064 -14888 -34765 -14872
rect -41064 -14952 -34849 -14888
rect -34785 -14952 -34765 -14888
rect -41064 -14968 -34765 -14952
rect -41064 -15032 -34849 -14968
rect -34785 -15032 -34765 -14968
rect -41064 -15048 -34765 -15032
rect -41064 -15112 -34849 -15048
rect -34785 -15112 -34765 -15048
rect -41064 -15128 -34765 -15112
rect -41064 -15192 -34849 -15128
rect -34785 -15192 -34765 -15128
rect -41064 -15208 -34765 -15192
rect -41064 -15272 -34849 -15208
rect -34785 -15272 -34765 -15208
rect -41064 -15288 -34765 -15272
rect -41064 -15352 -34849 -15288
rect -34785 -15352 -34765 -15288
rect -41064 -15368 -34765 -15352
rect -41064 -15432 -34849 -15368
rect -34785 -15432 -34765 -15368
rect -41064 -15448 -34765 -15432
rect -41064 -15512 -34849 -15448
rect -34785 -15512 -34765 -15448
rect -41064 -15528 -34765 -15512
rect -41064 -15592 -34849 -15528
rect -34785 -15592 -34765 -15528
rect -41064 -15608 -34765 -15592
rect -41064 -15672 -34849 -15608
rect -34785 -15672 -34765 -15608
rect -41064 -15700 -34765 -15672
rect -34745 -9528 -28446 -9500
rect -34745 -9592 -28530 -9528
rect -28466 -9592 -28446 -9528
rect -34745 -9608 -28446 -9592
rect -34745 -9672 -28530 -9608
rect -28466 -9672 -28446 -9608
rect -34745 -9688 -28446 -9672
rect -34745 -9752 -28530 -9688
rect -28466 -9752 -28446 -9688
rect -34745 -9768 -28446 -9752
rect -34745 -9832 -28530 -9768
rect -28466 -9832 -28446 -9768
rect -34745 -9848 -28446 -9832
rect -34745 -9912 -28530 -9848
rect -28466 -9912 -28446 -9848
rect -34745 -9928 -28446 -9912
rect -34745 -9992 -28530 -9928
rect -28466 -9992 -28446 -9928
rect -34745 -10008 -28446 -9992
rect -34745 -10072 -28530 -10008
rect -28466 -10072 -28446 -10008
rect -34745 -10088 -28446 -10072
rect -34745 -10152 -28530 -10088
rect -28466 -10152 -28446 -10088
rect -34745 -10168 -28446 -10152
rect -34745 -10232 -28530 -10168
rect -28466 -10232 -28446 -10168
rect -34745 -10248 -28446 -10232
rect -34745 -10312 -28530 -10248
rect -28466 -10312 -28446 -10248
rect -34745 -10328 -28446 -10312
rect -34745 -10392 -28530 -10328
rect -28466 -10392 -28446 -10328
rect -34745 -10408 -28446 -10392
rect -34745 -10472 -28530 -10408
rect -28466 -10472 -28446 -10408
rect -34745 -10488 -28446 -10472
rect -34745 -10552 -28530 -10488
rect -28466 -10552 -28446 -10488
rect -34745 -10568 -28446 -10552
rect -34745 -10632 -28530 -10568
rect -28466 -10632 -28446 -10568
rect -34745 -10648 -28446 -10632
rect -34745 -10712 -28530 -10648
rect -28466 -10712 -28446 -10648
rect -34745 -10728 -28446 -10712
rect -34745 -10792 -28530 -10728
rect -28466 -10792 -28446 -10728
rect -34745 -10808 -28446 -10792
rect -34745 -10872 -28530 -10808
rect -28466 -10872 -28446 -10808
rect -34745 -10888 -28446 -10872
rect -34745 -10952 -28530 -10888
rect -28466 -10952 -28446 -10888
rect -34745 -10968 -28446 -10952
rect -34745 -11032 -28530 -10968
rect -28466 -11032 -28446 -10968
rect -34745 -11048 -28446 -11032
rect -34745 -11112 -28530 -11048
rect -28466 -11112 -28446 -11048
rect -34745 -11128 -28446 -11112
rect -34745 -11192 -28530 -11128
rect -28466 -11192 -28446 -11128
rect -34745 -11208 -28446 -11192
rect -34745 -11272 -28530 -11208
rect -28466 -11272 -28446 -11208
rect -34745 -11288 -28446 -11272
rect -34745 -11352 -28530 -11288
rect -28466 -11352 -28446 -11288
rect -34745 -11368 -28446 -11352
rect -34745 -11432 -28530 -11368
rect -28466 -11432 -28446 -11368
rect -34745 -11448 -28446 -11432
rect -34745 -11512 -28530 -11448
rect -28466 -11512 -28446 -11448
rect -34745 -11528 -28446 -11512
rect -34745 -11592 -28530 -11528
rect -28466 -11592 -28446 -11528
rect -34745 -11608 -28446 -11592
rect -34745 -11672 -28530 -11608
rect -28466 -11672 -28446 -11608
rect -34745 -11688 -28446 -11672
rect -34745 -11752 -28530 -11688
rect -28466 -11752 -28446 -11688
rect -34745 -11768 -28446 -11752
rect -34745 -11832 -28530 -11768
rect -28466 -11832 -28446 -11768
rect -34745 -11848 -28446 -11832
rect -34745 -11912 -28530 -11848
rect -28466 -11912 -28446 -11848
rect -34745 -11928 -28446 -11912
rect -34745 -11992 -28530 -11928
rect -28466 -11992 -28446 -11928
rect -34745 -12008 -28446 -11992
rect -34745 -12072 -28530 -12008
rect -28466 -12072 -28446 -12008
rect -34745 -12088 -28446 -12072
rect -34745 -12152 -28530 -12088
rect -28466 -12152 -28446 -12088
rect -34745 -12168 -28446 -12152
rect -34745 -12232 -28530 -12168
rect -28466 -12232 -28446 -12168
rect -34745 -12248 -28446 -12232
rect -34745 -12312 -28530 -12248
rect -28466 -12312 -28446 -12248
rect -34745 -12328 -28446 -12312
rect -34745 -12392 -28530 -12328
rect -28466 -12392 -28446 -12328
rect -34745 -12408 -28446 -12392
rect -34745 -12472 -28530 -12408
rect -28466 -12472 -28446 -12408
rect -34745 -12488 -28446 -12472
rect -34745 -12552 -28530 -12488
rect -28466 -12552 -28446 -12488
rect -34745 -12568 -28446 -12552
rect -34745 -12632 -28530 -12568
rect -28466 -12632 -28446 -12568
rect -34745 -12648 -28446 -12632
rect -34745 -12712 -28530 -12648
rect -28466 -12712 -28446 -12648
rect -34745 -12728 -28446 -12712
rect -34745 -12792 -28530 -12728
rect -28466 -12792 -28446 -12728
rect -34745 -12808 -28446 -12792
rect -34745 -12872 -28530 -12808
rect -28466 -12872 -28446 -12808
rect -34745 -12888 -28446 -12872
rect -34745 -12952 -28530 -12888
rect -28466 -12952 -28446 -12888
rect -34745 -12968 -28446 -12952
rect -34745 -13032 -28530 -12968
rect -28466 -13032 -28446 -12968
rect -34745 -13048 -28446 -13032
rect -34745 -13112 -28530 -13048
rect -28466 -13112 -28446 -13048
rect -34745 -13128 -28446 -13112
rect -34745 -13192 -28530 -13128
rect -28466 -13192 -28446 -13128
rect -34745 -13208 -28446 -13192
rect -34745 -13272 -28530 -13208
rect -28466 -13272 -28446 -13208
rect -34745 -13288 -28446 -13272
rect -34745 -13352 -28530 -13288
rect -28466 -13352 -28446 -13288
rect -34745 -13368 -28446 -13352
rect -34745 -13432 -28530 -13368
rect -28466 -13432 -28446 -13368
rect -34745 -13448 -28446 -13432
rect -34745 -13512 -28530 -13448
rect -28466 -13512 -28446 -13448
rect -34745 -13528 -28446 -13512
rect -34745 -13592 -28530 -13528
rect -28466 -13592 -28446 -13528
rect -34745 -13608 -28446 -13592
rect -34745 -13672 -28530 -13608
rect -28466 -13672 -28446 -13608
rect -34745 -13688 -28446 -13672
rect -34745 -13752 -28530 -13688
rect -28466 -13752 -28446 -13688
rect -34745 -13768 -28446 -13752
rect -34745 -13832 -28530 -13768
rect -28466 -13832 -28446 -13768
rect -34745 -13848 -28446 -13832
rect -34745 -13912 -28530 -13848
rect -28466 -13912 -28446 -13848
rect -34745 -13928 -28446 -13912
rect -34745 -13992 -28530 -13928
rect -28466 -13992 -28446 -13928
rect -34745 -14008 -28446 -13992
rect -34745 -14072 -28530 -14008
rect -28466 -14072 -28446 -14008
rect -34745 -14088 -28446 -14072
rect -34745 -14152 -28530 -14088
rect -28466 -14152 -28446 -14088
rect -34745 -14168 -28446 -14152
rect -34745 -14232 -28530 -14168
rect -28466 -14232 -28446 -14168
rect -34745 -14248 -28446 -14232
rect -34745 -14312 -28530 -14248
rect -28466 -14312 -28446 -14248
rect -34745 -14328 -28446 -14312
rect -34745 -14392 -28530 -14328
rect -28466 -14392 -28446 -14328
rect -34745 -14408 -28446 -14392
rect -34745 -14472 -28530 -14408
rect -28466 -14472 -28446 -14408
rect -34745 -14488 -28446 -14472
rect -34745 -14552 -28530 -14488
rect -28466 -14552 -28446 -14488
rect -34745 -14568 -28446 -14552
rect -34745 -14632 -28530 -14568
rect -28466 -14632 -28446 -14568
rect -34745 -14648 -28446 -14632
rect -34745 -14712 -28530 -14648
rect -28466 -14712 -28446 -14648
rect -34745 -14728 -28446 -14712
rect -34745 -14792 -28530 -14728
rect -28466 -14792 -28446 -14728
rect -34745 -14808 -28446 -14792
rect -34745 -14872 -28530 -14808
rect -28466 -14872 -28446 -14808
rect -34745 -14888 -28446 -14872
rect -34745 -14952 -28530 -14888
rect -28466 -14952 -28446 -14888
rect -34745 -14968 -28446 -14952
rect -34745 -15032 -28530 -14968
rect -28466 -15032 -28446 -14968
rect -34745 -15048 -28446 -15032
rect -34745 -15112 -28530 -15048
rect -28466 -15112 -28446 -15048
rect -34745 -15128 -28446 -15112
rect -34745 -15192 -28530 -15128
rect -28466 -15192 -28446 -15128
rect -34745 -15208 -28446 -15192
rect -34745 -15272 -28530 -15208
rect -28466 -15272 -28446 -15208
rect -34745 -15288 -28446 -15272
rect -34745 -15352 -28530 -15288
rect -28466 -15352 -28446 -15288
rect -34745 -15368 -28446 -15352
rect -34745 -15432 -28530 -15368
rect -28466 -15432 -28446 -15368
rect -34745 -15448 -28446 -15432
rect -34745 -15512 -28530 -15448
rect -28466 -15512 -28446 -15448
rect -34745 -15528 -28446 -15512
rect -34745 -15592 -28530 -15528
rect -28466 -15592 -28446 -15528
rect -34745 -15608 -28446 -15592
rect -34745 -15672 -28530 -15608
rect -28466 -15672 -28446 -15608
rect -34745 -15700 -28446 -15672
rect -28426 -9528 -22127 -9500
rect -28426 -9592 -22211 -9528
rect -22147 -9592 -22127 -9528
rect -28426 -9608 -22127 -9592
rect -28426 -9672 -22211 -9608
rect -22147 -9672 -22127 -9608
rect -28426 -9688 -22127 -9672
rect -28426 -9752 -22211 -9688
rect -22147 -9752 -22127 -9688
rect -28426 -9768 -22127 -9752
rect -28426 -9832 -22211 -9768
rect -22147 -9832 -22127 -9768
rect -28426 -9848 -22127 -9832
rect -28426 -9912 -22211 -9848
rect -22147 -9912 -22127 -9848
rect -28426 -9928 -22127 -9912
rect -28426 -9992 -22211 -9928
rect -22147 -9992 -22127 -9928
rect -28426 -10008 -22127 -9992
rect -28426 -10072 -22211 -10008
rect -22147 -10072 -22127 -10008
rect -28426 -10088 -22127 -10072
rect -28426 -10152 -22211 -10088
rect -22147 -10152 -22127 -10088
rect -28426 -10168 -22127 -10152
rect -28426 -10232 -22211 -10168
rect -22147 -10232 -22127 -10168
rect -28426 -10248 -22127 -10232
rect -28426 -10312 -22211 -10248
rect -22147 -10312 -22127 -10248
rect -28426 -10328 -22127 -10312
rect -28426 -10392 -22211 -10328
rect -22147 -10392 -22127 -10328
rect -28426 -10408 -22127 -10392
rect -28426 -10472 -22211 -10408
rect -22147 -10472 -22127 -10408
rect -28426 -10488 -22127 -10472
rect -28426 -10552 -22211 -10488
rect -22147 -10552 -22127 -10488
rect -28426 -10568 -22127 -10552
rect -28426 -10632 -22211 -10568
rect -22147 -10632 -22127 -10568
rect -28426 -10648 -22127 -10632
rect -28426 -10712 -22211 -10648
rect -22147 -10712 -22127 -10648
rect -28426 -10728 -22127 -10712
rect -28426 -10792 -22211 -10728
rect -22147 -10792 -22127 -10728
rect -28426 -10808 -22127 -10792
rect -28426 -10872 -22211 -10808
rect -22147 -10872 -22127 -10808
rect -28426 -10888 -22127 -10872
rect -28426 -10952 -22211 -10888
rect -22147 -10952 -22127 -10888
rect -28426 -10968 -22127 -10952
rect -28426 -11032 -22211 -10968
rect -22147 -11032 -22127 -10968
rect -28426 -11048 -22127 -11032
rect -28426 -11112 -22211 -11048
rect -22147 -11112 -22127 -11048
rect -28426 -11128 -22127 -11112
rect -28426 -11192 -22211 -11128
rect -22147 -11192 -22127 -11128
rect -28426 -11208 -22127 -11192
rect -28426 -11272 -22211 -11208
rect -22147 -11272 -22127 -11208
rect -28426 -11288 -22127 -11272
rect -28426 -11352 -22211 -11288
rect -22147 -11352 -22127 -11288
rect -28426 -11368 -22127 -11352
rect -28426 -11432 -22211 -11368
rect -22147 -11432 -22127 -11368
rect -28426 -11448 -22127 -11432
rect -28426 -11512 -22211 -11448
rect -22147 -11512 -22127 -11448
rect -28426 -11528 -22127 -11512
rect -28426 -11592 -22211 -11528
rect -22147 -11592 -22127 -11528
rect -28426 -11608 -22127 -11592
rect -28426 -11672 -22211 -11608
rect -22147 -11672 -22127 -11608
rect -28426 -11688 -22127 -11672
rect -28426 -11752 -22211 -11688
rect -22147 -11752 -22127 -11688
rect -28426 -11768 -22127 -11752
rect -28426 -11832 -22211 -11768
rect -22147 -11832 -22127 -11768
rect -28426 -11848 -22127 -11832
rect -28426 -11912 -22211 -11848
rect -22147 -11912 -22127 -11848
rect -28426 -11928 -22127 -11912
rect -28426 -11992 -22211 -11928
rect -22147 -11992 -22127 -11928
rect -28426 -12008 -22127 -11992
rect -28426 -12072 -22211 -12008
rect -22147 -12072 -22127 -12008
rect -28426 -12088 -22127 -12072
rect -28426 -12152 -22211 -12088
rect -22147 -12152 -22127 -12088
rect -28426 -12168 -22127 -12152
rect -28426 -12232 -22211 -12168
rect -22147 -12232 -22127 -12168
rect -28426 -12248 -22127 -12232
rect -28426 -12312 -22211 -12248
rect -22147 -12312 -22127 -12248
rect -28426 -12328 -22127 -12312
rect -28426 -12392 -22211 -12328
rect -22147 -12392 -22127 -12328
rect -28426 -12408 -22127 -12392
rect -28426 -12472 -22211 -12408
rect -22147 -12472 -22127 -12408
rect -28426 -12488 -22127 -12472
rect -28426 -12552 -22211 -12488
rect -22147 -12552 -22127 -12488
rect -28426 -12568 -22127 -12552
rect -28426 -12632 -22211 -12568
rect -22147 -12632 -22127 -12568
rect -28426 -12648 -22127 -12632
rect -28426 -12712 -22211 -12648
rect -22147 -12712 -22127 -12648
rect -28426 -12728 -22127 -12712
rect -28426 -12792 -22211 -12728
rect -22147 -12792 -22127 -12728
rect -28426 -12808 -22127 -12792
rect -28426 -12872 -22211 -12808
rect -22147 -12872 -22127 -12808
rect -28426 -12888 -22127 -12872
rect -28426 -12952 -22211 -12888
rect -22147 -12952 -22127 -12888
rect -28426 -12968 -22127 -12952
rect -28426 -13032 -22211 -12968
rect -22147 -13032 -22127 -12968
rect -28426 -13048 -22127 -13032
rect -28426 -13112 -22211 -13048
rect -22147 -13112 -22127 -13048
rect -28426 -13128 -22127 -13112
rect -28426 -13192 -22211 -13128
rect -22147 -13192 -22127 -13128
rect -28426 -13208 -22127 -13192
rect -28426 -13272 -22211 -13208
rect -22147 -13272 -22127 -13208
rect -28426 -13288 -22127 -13272
rect -28426 -13352 -22211 -13288
rect -22147 -13352 -22127 -13288
rect -28426 -13368 -22127 -13352
rect -28426 -13432 -22211 -13368
rect -22147 -13432 -22127 -13368
rect -28426 -13448 -22127 -13432
rect -28426 -13512 -22211 -13448
rect -22147 -13512 -22127 -13448
rect -28426 -13528 -22127 -13512
rect -28426 -13592 -22211 -13528
rect -22147 -13592 -22127 -13528
rect -28426 -13608 -22127 -13592
rect -28426 -13672 -22211 -13608
rect -22147 -13672 -22127 -13608
rect -28426 -13688 -22127 -13672
rect -28426 -13752 -22211 -13688
rect -22147 -13752 -22127 -13688
rect -28426 -13768 -22127 -13752
rect -28426 -13832 -22211 -13768
rect -22147 -13832 -22127 -13768
rect -28426 -13848 -22127 -13832
rect -28426 -13912 -22211 -13848
rect -22147 -13912 -22127 -13848
rect -28426 -13928 -22127 -13912
rect -28426 -13992 -22211 -13928
rect -22147 -13992 -22127 -13928
rect -28426 -14008 -22127 -13992
rect -28426 -14072 -22211 -14008
rect -22147 -14072 -22127 -14008
rect -28426 -14088 -22127 -14072
rect -28426 -14152 -22211 -14088
rect -22147 -14152 -22127 -14088
rect -28426 -14168 -22127 -14152
rect -28426 -14232 -22211 -14168
rect -22147 -14232 -22127 -14168
rect -28426 -14248 -22127 -14232
rect -28426 -14312 -22211 -14248
rect -22147 -14312 -22127 -14248
rect -28426 -14328 -22127 -14312
rect -28426 -14392 -22211 -14328
rect -22147 -14392 -22127 -14328
rect -28426 -14408 -22127 -14392
rect -28426 -14472 -22211 -14408
rect -22147 -14472 -22127 -14408
rect -28426 -14488 -22127 -14472
rect -28426 -14552 -22211 -14488
rect -22147 -14552 -22127 -14488
rect -28426 -14568 -22127 -14552
rect -28426 -14632 -22211 -14568
rect -22147 -14632 -22127 -14568
rect -28426 -14648 -22127 -14632
rect -28426 -14712 -22211 -14648
rect -22147 -14712 -22127 -14648
rect -28426 -14728 -22127 -14712
rect -28426 -14792 -22211 -14728
rect -22147 -14792 -22127 -14728
rect -28426 -14808 -22127 -14792
rect -28426 -14872 -22211 -14808
rect -22147 -14872 -22127 -14808
rect -28426 -14888 -22127 -14872
rect -28426 -14952 -22211 -14888
rect -22147 -14952 -22127 -14888
rect -28426 -14968 -22127 -14952
rect -28426 -15032 -22211 -14968
rect -22147 -15032 -22127 -14968
rect -28426 -15048 -22127 -15032
rect -28426 -15112 -22211 -15048
rect -22147 -15112 -22127 -15048
rect -28426 -15128 -22127 -15112
rect -28426 -15192 -22211 -15128
rect -22147 -15192 -22127 -15128
rect -28426 -15208 -22127 -15192
rect -28426 -15272 -22211 -15208
rect -22147 -15272 -22127 -15208
rect -28426 -15288 -22127 -15272
rect -28426 -15352 -22211 -15288
rect -22147 -15352 -22127 -15288
rect -28426 -15368 -22127 -15352
rect -28426 -15432 -22211 -15368
rect -22147 -15432 -22127 -15368
rect -28426 -15448 -22127 -15432
rect -28426 -15512 -22211 -15448
rect -22147 -15512 -22127 -15448
rect -28426 -15528 -22127 -15512
rect -28426 -15592 -22211 -15528
rect -22147 -15592 -22127 -15528
rect -28426 -15608 -22127 -15592
rect -28426 -15672 -22211 -15608
rect -22147 -15672 -22127 -15608
rect -28426 -15700 -22127 -15672
rect -22107 -9528 -15808 -9500
rect -22107 -9592 -15892 -9528
rect -15828 -9592 -15808 -9528
rect -22107 -9608 -15808 -9592
rect -22107 -9672 -15892 -9608
rect -15828 -9672 -15808 -9608
rect -22107 -9688 -15808 -9672
rect -22107 -9752 -15892 -9688
rect -15828 -9752 -15808 -9688
rect -22107 -9768 -15808 -9752
rect -22107 -9832 -15892 -9768
rect -15828 -9832 -15808 -9768
rect -22107 -9848 -15808 -9832
rect -22107 -9912 -15892 -9848
rect -15828 -9912 -15808 -9848
rect -22107 -9928 -15808 -9912
rect -22107 -9992 -15892 -9928
rect -15828 -9992 -15808 -9928
rect -22107 -10008 -15808 -9992
rect -22107 -10072 -15892 -10008
rect -15828 -10072 -15808 -10008
rect -22107 -10088 -15808 -10072
rect -22107 -10152 -15892 -10088
rect -15828 -10152 -15808 -10088
rect -22107 -10168 -15808 -10152
rect -22107 -10232 -15892 -10168
rect -15828 -10232 -15808 -10168
rect -22107 -10248 -15808 -10232
rect -22107 -10312 -15892 -10248
rect -15828 -10312 -15808 -10248
rect -22107 -10328 -15808 -10312
rect -22107 -10392 -15892 -10328
rect -15828 -10392 -15808 -10328
rect -22107 -10408 -15808 -10392
rect -22107 -10472 -15892 -10408
rect -15828 -10472 -15808 -10408
rect -22107 -10488 -15808 -10472
rect -22107 -10552 -15892 -10488
rect -15828 -10552 -15808 -10488
rect -22107 -10568 -15808 -10552
rect -22107 -10632 -15892 -10568
rect -15828 -10632 -15808 -10568
rect -22107 -10648 -15808 -10632
rect -22107 -10712 -15892 -10648
rect -15828 -10712 -15808 -10648
rect -22107 -10728 -15808 -10712
rect -22107 -10792 -15892 -10728
rect -15828 -10792 -15808 -10728
rect -22107 -10808 -15808 -10792
rect -22107 -10872 -15892 -10808
rect -15828 -10872 -15808 -10808
rect -22107 -10888 -15808 -10872
rect -22107 -10952 -15892 -10888
rect -15828 -10952 -15808 -10888
rect -22107 -10968 -15808 -10952
rect -22107 -11032 -15892 -10968
rect -15828 -11032 -15808 -10968
rect -22107 -11048 -15808 -11032
rect -22107 -11112 -15892 -11048
rect -15828 -11112 -15808 -11048
rect -22107 -11128 -15808 -11112
rect -22107 -11192 -15892 -11128
rect -15828 -11192 -15808 -11128
rect -22107 -11208 -15808 -11192
rect -22107 -11272 -15892 -11208
rect -15828 -11272 -15808 -11208
rect -22107 -11288 -15808 -11272
rect -22107 -11352 -15892 -11288
rect -15828 -11352 -15808 -11288
rect -22107 -11368 -15808 -11352
rect -22107 -11432 -15892 -11368
rect -15828 -11432 -15808 -11368
rect -22107 -11448 -15808 -11432
rect -22107 -11512 -15892 -11448
rect -15828 -11512 -15808 -11448
rect -22107 -11528 -15808 -11512
rect -22107 -11592 -15892 -11528
rect -15828 -11592 -15808 -11528
rect -22107 -11608 -15808 -11592
rect -22107 -11672 -15892 -11608
rect -15828 -11672 -15808 -11608
rect -22107 -11688 -15808 -11672
rect -22107 -11752 -15892 -11688
rect -15828 -11752 -15808 -11688
rect -22107 -11768 -15808 -11752
rect -22107 -11832 -15892 -11768
rect -15828 -11832 -15808 -11768
rect -22107 -11848 -15808 -11832
rect -22107 -11912 -15892 -11848
rect -15828 -11912 -15808 -11848
rect -22107 -11928 -15808 -11912
rect -22107 -11992 -15892 -11928
rect -15828 -11992 -15808 -11928
rect -22107 -12008 -15808 -11992
rect -22107 -12072 -15892 -12008
rect -15828 -12072 -15808 -12008
rect -22107 -12088 -15808 -12072
rect -22107 -12152 -15892 -12088
rect -15828 -12152 -15808 -12088
rect -22107 -12168 -15808 -12152
rect -22107 -12232 -15892 -12168
rect -15828 -12232 -15808 -12168
rect -22107 -12248 -15808 -12232
rect -22107 -12312 -15892 -12248
rect -15828 -12312 -15808 -12248
rect -22107 -12328 -15808 -12312
rect -22107 -12392 -15892 -12328
rect -15828 -12392 -15808 -12328
rect -22107 -12408 -15808 -12392
rect -22107 -12472 -15892 -12408
rect -15828 -12472 -15808 -12408
rect -22107 -12488 -15808 -12472
rect -22107 -12552 -15892 -12488
rect -15828 -12552 -15808 -12488
rect -22107 -12568 -15808 -12552
rect -22107 -12632 -15892 -12568
rect -15828 -12632 -15808 -12568
rect -22107 -12648 -15808 -12632
rect -22107 -12712 -15892 -12648
rect -15828 -12712 -15808 -12648
rect -22107 -12728 -15808 -12712
rect -22107 -12792 -15892 -12728
rect -15828 -12792 -15808 -12728
rect -22107 -12808 -15808 -12792
rect -22107 -12872 -15892 -12808
rect -15828 -12872 -15808 -12808
rect -22107 -12888 -15808 -12872
rect -22107 -12952 -15892 -12888
rect -15828 -12952 -15808 -12888
rect -22107 -12968 -15808 -12952
rect -22107 -13032 -15892 -12968
rect -15828 -13032 -15808 -12968
rect -22107 -13048 -15808 -13032
rect -22107 -13112 -15892 -13048
rect -15828 -13112 -15808 -13048
rect -22107 -13128 -15808 -13112
rect -22107 -13192 -15892 -13128
rect -15828 -13192 -15808 -13128
rect -22107 -13208 -15808 -13192
rect -22107 -13272 -15892 -13208
rect -15828 -13272 -15808 -13208
rect -22107 -13288 -15808 -13272
rect -22107 -13352 -15892 -13288
rect -15828 -13352 -15808 -13288
rect -22107 -13368 -15808 -13352
rect -22107 -13432 -15892 -13368
rect -15828 -13432 -15808 -13368
rect -22107 -13448 -15808 -13432
rect -22107 -13512 -15892 -13448
rect -15828 -13512 -15808 -13448
rect -22107 -13528 -15808 -13512
rect -22107 -13592 -15892 -13528
rect -15828 -13592 -15808 -13528
rect -22107 -13608 -15808 -13592
rect -22107 -13672 -15892 -13608
rect -15828 -13672 -15808 -13608
rect -22107 -13688 -15808 -13672
rect -22107 -13752 -15892 -13688
rect -15828 -13752 -15808 -13688
rect -22107 -13768 -15808 -13752
rect -22107 -13832 -15892 -13768
rect -15828 -13832 -15808 -13768
rect -22107 -13848 -15808 -13832
rect -22107 -13912 -15892 -13848
rect -15828 -13912 -15808 -13848
rect -22107 -13928 -15808 -13912
rect -22107 -13992 -15892 -13928
rect -15828 -13992 -15808 -13928
rect -22107 -14008 -15808 -13992
rect -22107 -14072 -15892 -14008
rect -15828 -14072 -15808 -14008
rect -22107 -14088 -15808 -14072
rect -22107 -14152 -15892 -14088
rect -15828 -14152 -15808 -14088
rect -22107 -14168 -15808 -14152
rect -22107 -14232 -15892 -14168
rect -15828 -14232 -15808 -14168
rect -22107 -14248 -15808 -14232
rect -22107 -14312 -15892 -14248
rect -15828 -14312 -15808 -14248
rect -22107 -14328 -15808 -14312
rect -22107 -14392 -15892 -14328
rect -15828 -14392 -15808 -14328
rect -22107 -14408 -15808 -14392
rect -22107 -14472 -15892 -14408
rect -15828 -14472 -15808 -14408
rect -22107 -14488 -15808 -14472
rect -22107 -14552 -15892 -14488
rect -15828 -14552 -15808 -14488
rect -22107 -14568 -15808 -14552
rect -22107 -14632 -15892 -14568
rect -15828 -14632 -15808 -14568
rect -22107 -14648 -15808 -14632
rect -22107 -14712 -15892 -14648
rect -15828 -14712 -15808 -14648
rect -22107 -14728 -15808 -14712
rect -22107 -14792 -15892 -14728
rect -15828 -14792 -15808 -14728
rect -22107 -14808 -15808 -14792
rect -22107 -14872 -15892 -14808
rect -15828 -14872 -15808 -14808
rect -22107 -14888 -15808 -14872
rect -22107 -14952 -15892 -14888
rect -15828 -14952 -15808 -14888
rect -22107 -14968 -15808 -14952
rect -22107 -15032 -15892 -14968
rect -15828 -15032 -15808 -14968
rect -22107 -15048 -15808 -15032
rect -22107 -15112 -15892 -15048
rect -15828 -15112 -15808 -15048
rect -22107 -15128 -15808 -15112
rect -22107 -15192 -15892 -15128
rect -15828 -15192 -15808 -15128
rect -22107 -15208 -15808 -15192
rect -22107 -15272 -15892 -15208
rect -15828 -15272 -15808 -15208
rect -22107 -15288 -15808 -15272
rect -22107 -15352 -15892 -15288
rect -15828 -15352 -15808 -15288
rect -22107 -15368 -15808 -15352
rect -22107 -15432 -15892 -15368
rect -15828 -15432 -15808 -15368
rect -22107 -15448 -15808 -15432
rect -22107 -15512 -15892 -15448
rect -15828 -15512 -15808 -15448
rect -22107 -15528 -15808 -15512
rect -22107 -15592 -15892 -15528
rect -15828 -15592 -15808 -15528
rect -22107 -15608 -15808 -15592
rect -22107 -15672 -15892 -15608
rect -15828 -15672 -15808 -15608
rect -22107 -15700 -15808 -15672
rect -15788 -9528 -9489 -9500
rect -15788 -9592 -9573 -9528
rect -9509 -9592 -9489 -9528
rect -15788 -9608 -9489 -9592
rect -15788 -9672 -9573 -9608
rect -9509 -9672 -9489 -9608
rect -15788 -9688 -9489 -9672
rect -15788 -9752 -9573 -9688
rect -9509 -9752 -9489 -9688
rect -15788 -9768 -9489 -9752
rect -15788 -9832 -9573 -9768
rect -9509 -9832 -9489 -9768
rect -15788 -9848 -9489 -9832
rect -15788 -9912 -9573 -9848
rect -9509 -9912 -9489 -9848
rect -15788 -9928 -9489 -9912
rect -15788 -9992 -9573 -9928
rect -9509 -9992 -9489 -9928
rect -15788 -10008 -9489 -9992
rect -15788 -10072 -9573 -10008
rect -9509 -10072 -9489 -10008
rect -15788 -10088 -9489 -10072
rect -15788 -10152 -9573 -10088
rect -9509 -10152 -9489 -10088
rect -15788 -10168 -9489 -10152
rect -15788 -10232 -9573 -10168
rect -9509 -10232 -9489 -10168
rect -15788 -10248 -9489 -10232
rect -15788 -10312 -9573 -10248
rect -9509 -10312 -9489 -10248
rect -15788 -10328 -9489 -10312
rect -15788 -10392 -9573 -10328
rect -9509 -10392 -9489 -10328
rect -15788 -10408 -9489 -10392
rect -15788 -10472 -9573 -10408
rect -9509 -10472 -9489 -10408
rect -15788 -10488 -9489 -10472
rect -15788 -10552 -9573 -10488
rect -9509 -10552 -9489 -10488
rect -15788 -10568 -9489 -10552
rect -15788 -10632 -9573 -10568
rect -9509 -10632 -9489 -10568
rect -15788 -10648 -9489 -10632
rect -15788 -10712 -9573 -10648
rect -9509 -10712 -9489 -10648
rect -15788 -10728 -9489 -10712
rect -15788 -10792 -9573 -10728
rect -9509 -10792 -9489 -10728
rect -15788 -10808 -9489 -10792
rect -15788 -10872 -9573 -10808
rect -9509 -10872 -9489 -10808
rect -15788 -10888 -9489 -10872
rect -15788 -10952 -9573 -10888
rect -9509 -10952 -9489 -10888
rect -15788 -10968 -9489 -10952
rect -15788 -11032 -9573 -10968
rect -9509 -11032 -9489 -10968
rect -15788 -11048 -9489 -11032
rect -15788 -11112 -9573 -11048
rect -9509 -11112 -9489 -11048
rect -15788 -11128 -9489 -11112
rect -15788 -11192 -9573 -11128
rect -9509 -11192 -9489 -11128
rect -15788 -11208 -9489 -11192
rect -15788 -11272 -9573 -11208
rect -9509 -11272 -9489 -11208
rect -15788 -11288 -9489 -11272
rect -15788 -11352 -9573 -11288
rect -9509 -11352 -9489 -11288
rect -15788 -11368 -9489 -11352
rect -15788 -11432 -9573 -11368
rect -9509 -11432 -9489 -11368
rect -15788 -11448 -9489 -11432
rect -15788 -11512 -9573 -11448
rect -9509 -11512 -9489 -11448
rect -15788 -11528 -9489 -11512
rect -15788 -11592 -9573 -11528
rect -9509 -11592 -9489 -11528
rect -15788 -11608 -9489 -11592
rect -15788 -11672 -9573 -11608
rect -9509 -11672 -9489 -11608
rect -15788 -11688 -9489 -11672
rect -15788 -11752 -9573 -11688
rect -9509 -11752 -9489 -11688
rect -15788 -11768 -9489 -11752
rect -15788 -11832 -9573 -11768
rect -9509 -11832 -9489 -11768
rect -15788 -11848 -9489 -11832
rect -15788 -11912 -9573 -11848
rect -9509 -11912 -9489 -11848
rect -15788 -11928 -9489 -11912
rect -15788 -11992 -9573 -11928
rect -9509 -11992 -9489 -11928
rect -15788 -12008 -9489 -11992
rect -15788 -12072 -9573 -12008
rect -9509 -12072 -9489 -12008
rect -15788 -12088 -9489 -12072
rect -15788 -12152 -9573 -12088
rect -9509 -12152 -9489 -12088
rect -15788 -12168 -9489 -12152
rect -15788 -12232 -9573 -12168
rect -9509 -12232 -9489 -12168
rect -15788 -12248 -9489 -12232
rect -15788 -12312 -9573 -12248
rect -9509 -12312 -9489 -12248
rect -15788 -12328 -9489 -12312
rect -15788 -12392 -9573 -12328
rect -9509 -12392 -9489 -12328
rect -15788 -12408 -9489 -12392
rect -15788 -12472 -9573 -12408
rect -9509 -12472 -9489 -12408
rect -15788 -12488 -9489 -12472
rect -15788 -12552 -9573 -12488
rect -9509 -12552 -9489 -12488
rect -15788 -12568 -9489 -12552
rect -15788 -12632 -9573 -12568
rect -9509 -12632 -9489 -12568
rect -15788 -12648 -9489 -12632
rect -15788 -12712 -9573 -12648
rect -9509 -12712 -9489 -12648
rect -15788 -12728 -9489 -12712
rect -15788 -12792 -9573 -12728
rect -9509 -12792 -9489 -12728
rect -15788 -12808 -9489 -12792
rect -15788 -12872 -9573 -12808
rect -9509 -12872 -9489 -12808
rect -15788 -12888 -9489 -12872
rect -15788 -12952 -9573 -12888
rect -9509 -12952 -9489 -12888
rect -15788 -12968 -9489 -12952
rect -15788 -13032 -9573 -12968
rect -9509 -13032 -9489 -12968
rect -15788 -13048 -9489 -13032
rect -15788 -13112 -9573 -13048
rect -9509 -13112 -9489 -13048
rect -15788 -13128 -9489 -13112
rect -15788 -13192 -9573 -13128
rect -9509 -13192 -9489 -13128
rect -15788 -13208 -9489 -13192
rect -15788 -13272 -9573 -13208
rect -9509 -13272 -9489 -13208
rect -15788 -13288 -9489 -13272
rect -15788 -13352 -9573 -13288
rect -9509 -13352 -9489 -13288
rect -15788 -13368 -9489 -13352
rect -15788 -13432 -9573 -13368
rect -9509 -13432 -9489 -13368
rect -15788 -13448 -9489 -13432
rect -15788 -13512 -9573 -13448
rect -9509 -13512 -9489 -13448
rect -15788 -13528 -9489 -13512
rect -15788 -13592 -9573 -13528
rect -9509 -13592 -9489 -13528
rect -15788 -13608 -9489 -13592
rect -15788 -13672 -9573 -13608
rect -9509 -13672 -9489 -13608
rect -15788 -13688 -9489 -13672
rect -15788 -13752 -9573 -13688
rect -9509 -13752 -9489 -13688
rect -15788 -13768 -9489 -13752
rect -15788 -13832 -9573 -13768
rect -9509 -13832 -9489 -13768
rect -15788 -13848 -9489 -13832
rect -15788 -13912 -9573 -13848
rect -9509 -13912 -9489 -13848
rect -15788 -13928 -9489 -13912
rect -15788 -13992 -9573 -13928
rect -9509 -13992 -9489 -13928
rect -15788 -14008 -9489 -13992
rect -15788 -14072 -9573 -14008
rect -9509 -14072 -9489 -14008
rect -15788 -14088 -9489 -14072
rect -15788 -14152 -9573 -14088
rect -9509 -14152 -9489 -14088
rect -15788 -14168 -9489 -14152
rect -15788 -14232 -9573 -14168
rect -9509 -14232 -9489 -14168
rect -15788 -14248 -9489 -14232
rect -15788 -14312 -9573 -14248
rect -9509 -14312 -9489 -14248
rect -15788 -14328 -9489 -14312
rect -15788 -14392 -9573 -14328
rect -9509 -14392 -9489 -14328
rect -15788 -14408 -9489 -14392
rect -15788 -14472 -9573 -14408
rect -9509 -14472 -9489 -14408
rect -15788 -14488 -9489 -14472
rect -15788 -14552 -9573 -14488
rect -9509 -14552 -9489 -14488
rect -15788 -14568 -9489 -14552
rect -15788 -14632 -9573 -14568
rect -9509 -14632 -9489 -14568
rect -15788 -14648 -9489 -14632
rect -15788 -14712 -9573 -14648
rect -9509 -14712 -9489 -14648
rect -15788 -14728 -9489 -14712
rect -15788 -14792 -9573 -14728
rect -9509 -14792 -9489 -14728
rect -15788 -14808 -9489 -14792
rect -15788 -14872 -9573 -14808
rect -9509 -14872 -9489 -14808
rect -15788 -14888 -9489 -14872
rect -15788 -14952 -9573 -14888
rect -9509 -14952 -9489 -14888
rect -15788 -14968 -9489 -14952
rect -15788 -15032 -9573 -14968
rect -9509 -15032 -9489 -14968
rect -15788 -15048 -9489 -15032
rect -15788 -15112 -9573 -15048
rect -9509 -15112 -9489 -15048
rect -15788 -15128 -9489 -15112
rect -15788 -15192 -9573 -15128
rect -9509 -15192 -9489 -15128
rect -15788 -15208 -9489 -15192
rect -15788 -15272 -9573 -15208
rect -9509 -15272 -9489 -15208
rect -15788 -15288 -9489 -15272
rect -15788 -15352 -9573 -15288
rect -9509 -15352 -9489 -15288
rect -15788 -15368 -9489 -15352
rect -15788 -15432 -9573 -15368
rect -9509 -15432 -9489 -15368
rect -15788 -15448 -9489 -15432
rect -15788 -15512 -9573 -15448
rect -9509 -15512 -9489 -15448
rect -15788 -15528 -9489 -15512
rect -15788 -15592 -9573 -15528
rect -9509 -15592 -9489 -15528
rect -15788 -15608 -9489 -15592
rect -15788 -15672 -9573 -15608
rect -9509 -15672 -9489 -15608
rect -15788 -15700 -9489 -15672
rect -9469 -9528 -3170 -9500
rect -9469 -9592 -3254 -9528
rect -3190 -9592 -3170 -9528
rect -9469 -9608 -3170 -9592
rect -9469 -9672 -3254 -9608
rect -3190 -9672 -3170 -9608
rect -9469 -9688 -3170 -9672
rect -9469 -9752 -3254 -9688
rect -3190 -9752 -3170 -9688
rect -9469 -9768 -3170 -9752
rect -9469 -9832 -3254 -9768
rect -3190 -9832 -3170 -9768
rect -9469 -9848 -3170 -9832
rect -9469 -9912 -3254 -9848
rect -3190 -9912 -3170 -9848
rect -9469 -9928 -3170 -9912
rect -9469 -9992 -3254 -9928
rect -3190 -9992 -3170 -9928
rect -9469 -10008 -3170 -9992
rect -9469 -10072 -3254 -10008
rect -3190 -10072 -3170 -10008
rect -9469 -10088 -3170 -10072
rect -9469 -10152 -3254 -10088
rect -3190 -10152 -3170 -10088
rect -9469 -10168 -3170 -10152
rect -9469 -10232 -3254 -10168
rect -3190 -10232 -3170 -10168
rect -9469 -10248 -3170 -10232
rect -9469 -10312 -3254 -10248
rect -3190 -10312 -3170 -10248
rect -9469 -10328 -3170 -10312
rect -9469 -10392 -3254 -10328
rect -3190 -10392 -3170 -10328
rect -9469 -10408 -3170 -10392
rect -9469 -10472 -3254 -10408
rect -3190 -10472 -3170 -10408
rect -9469 -10488 -3170 -10472
rect -9469 -10552 -3254 -10488
rect -3190 -10552 -3170 -10488
rect -9469 -10568 -3170 -10552
rect -9469 -10632 -3254 -10568
rect -3190 -10632 -3170 -10568
rect -9469 -10648 -3170 -10632
rect -9469 -10712 -3254 -10648
rect -3190 -10712 -3170 -10648
rect -9469 -10728 -3170 -10712
rect -9469 -10792 -3254 -10728
rect -3190 -10792 -3170 -10728
rect -9469 -10808 -3170 -10792
rect -9469 -10872 -3254 -10808
rect -3190 -10872 -3170 -10808
rect -9469 -10888 -3170 -10872
rect -9469 -10952 -3254 -10888
rect -3190 -10952 -3170 -10888
rect -9469 -10968 -3170 -10952
rect -9469 -11032 -3254 -10968
rect -3190 -11032 -3170 -10968
rect -9469 -11048 -3170 -11032
rect -9469 -11112 -3254 -11048
rect -3190 -11112 -3170 -11048
rect -9469 -11128 -3170 -11112
rect -9469 -11192 -3254 -11128
rect -3190 -11192 -3170 -11128
rect -9469 -11208 -3170 -11192
rect -9469 -11272 -3254 -11208
rect -3190 -11272 -3170 -11208
rect -9469 -11288 -3170 -11272
rect -9469 -11352 -3254 -11288
rect -3190 -11352 -3170 -11288
rect -9469 -11368 -3170 -11352
rect -9469 -11432 -3254 -11368
rect -3190 -11432 -3170 -11368
rect -9469 -11448 -3170 -11432
rect -9469 -11512 -3254 -11448
rect -3190 -11512 -3170 -11448
rect -9469 -11528 -3170 -11512
rect -9469 -11592 -3254 -11528
rect -3190 -11592 -3170 -11528
rect -9469 -11608 -3170 -11592
rect -9469 -11672 -3254 -11608
rect -3190 -11672 -3170 -11608
rect -9469 -11688 -3170 -11672
rect -9469 -11752 -3254 -11688
rect -3190 -11752 -3170 -11688
rect -9469 -11768 -3170 -11752
rect -9469 -11832 -3254 -11768
rect -3190 -11832 -3170 -11768
rect -9469 -11848 -3170 -11832
rect -9469 -11912 -3254 -11848
rect -3190 -11912 -3170 -11848
rect -9469 -11928 -3170 -11912
rect -9469 -11992 -3254 -11928
rect -3190 -11992 -3170 -11928
rect -9469 -12008 -3170 -11992
rect -9469 -12072 -3254 -12008
rect -3190 -12072 -3170 -12008
rect -9469 -12088 -3170 -12072
rect -9469 -12152 -3254 -12088
rect -3190 -12152 -3170 -12088
rect -9469 -12168 -3170 -12152
rect -9469 -12232 -3254 -12168
rect -3190 -12232 -3170 -12168
rect -9469 -12248 -3170 -12232
rect -9469 -12312 -3254 -12248
rect -3190 -12312 -3170 -12248
rect -9469 -12328 -3170 -12312
rect -9469 -12392 -3254 -12328
rect -3190 -12392 -3170 -12328
rect -9469 -12408 -3170 -12392
rect -9469 -12472 -3254 -12408
rect -3190 -12472 -3170 -12408
rect -9469 -12488 -3170 -12472
rect -9469 -12552 -3254 -12488
rect -3190 -12552 -3170 -12488
rect -9469 -12568 -3170 -12552
rect -9469 -12632 -3254 -12568
rect -3190 -12632 -3170 -12568
rect -9469 -12648 -3170 -12632
rect -9469 -12712 -3254 -12648
rect -3190 -12712 -3170 -12648
rect -9469 -12728 -3170 -12712
rect -9469 -12792 -3254 -12728
rect -3190 -12792 -3170 -12728
rect -9469 -12808 -3170 -12792
rect -9469 -12872 -3254 -12808
rect -3190 -12872 -3170 -12808
rect -9469 -12888 -3170 -12872
rect -9469 -12952 -3254 -12888
rect -3190 -12952 -3170 -12888
rect -9469 -12968 -3170 -12952
rect -9469 -13032 -3254 -12968
rect -3190 -13032 -3170 -12968
rect -9469 -13048 -3170 -13032
rect -9469 -13112 -3254 -13048
rect -3190 -13112 -3170 -13048
rect -9469 -13128 -3170 -13112
rect -9469 -13192 -3254 -13128
rect -3190 -13192 -3170 -13128
rect -9469 -13208 -3170 -13192
rect -9469 -13272 -3254 -13208
rect -3190 -13272 -3170 -13208
rect -9469 -13288 -3170 -13272
rect -9469 -13352 -3254 -13288
rect -3190 -13352 -3170 -13288
rect -9469 -13368 -3170 -13352
rect -9469 -13432 -3254 -13368
rect -3190 -13432 -3170 -13368
rect -9469 -13448 -3170 -13432
rect -9469 -13512 -3254 -13448
rect -3190 -13512 -3170 -13448
rect -9469 -13528 -3170 -13512
rect -9469 -13592 -3254 -13528
rect -3190 -13592 -3170 -13528
rect -9469 -13608 -3170 -13592
rect -9469 -13672 -3254 -13608
rect -3190 -13672 -3170 -13608
rect -9469 -13688 -3170 -13672
rect -9469 -13752 -3254 -13688
rect -3190 -13752 -3170 -13688
rect -9469 -13768 -3170 -13752
rect -9469 -13832 -3254 -13768
rect -3190 -13832 -3170 -13768
rect -9469 -13848 -3170 -13832
rect -9469 -13912 -3254 -13848
rect -3190 -13912 -3170 -13848
rect -9469 -13928 -3170 -13912
rect -9469 -13992 -3254 -13928
rect -3190 -13992 -3170 -13928
rect -9469 -14008 -3170 -13992
rect -9469 -14072 -3254 -14008
rect -3190 -14072 -3170 -14008
rect -9469 -14088 -3170 -14072
rect -9469 -14152 -3254 -14088
rect -3190 -14152 -3170 -14088
rect -9469 -14168 -3170 -14152
rect -9469 -14232 -3254 -14168
rect -3190 -14232 -3170 -14168
rect -9469 -14248 -3170 -14232
rect -9469 -14312 -3254 -14248
rect -3190 -14312 -3170 -14248
rect -9469 -14328 -3170 -14312
rect -9469 -14392 -3254 -14328
rect -3190 -14392 -3170 -14328
rect -9469 -14408 -3170 -14392
rect -9469 -14472 -3254 -14408
rect -3190 -14472 -3170 -14408
rect -9469 -14488 -3170 -14472
rect -9469 -14552 -3254 -14488
rect -3190 -14552 -3170 -14488
rect -9469 -14568 -3170 -14552
rect -9469 -14632 -3254 -14568
rect -3190 -14632 -3170 -14568
rect -9469 -14648 -3170 -14632
rect -9469 -14712 -3254 -14648
rect -3190 -14712 -3170 -14648
rect -9469 -14728 -3170 -14712
rect -9469 -14792 -3254 -14728
rect -3190 -14792 -3170 -14728
rect -9469 -14808 -3170 -14792
rect -9469 -14872 -3254 -14808
rect -3190 -14872 -3170 -14808
rect -9469 -14888 -3170 -14872
rect -9469 -14952 -3254 -14888
rect -3190 -14952 -3170 -14888
rect -9469 -14968 -3170 -14952
rect -9469 -15032 -3254 -14968
rect -3190 -15032 -3170 -14968
rect -9469 -15048 -3170 -15032
rect -9469 -15112 -3254 -15048
rect -3190 -15112 -3170 -15048
rect -9469 -15128 -3170 -15112
rect -9469 -15192 -3254 -15128
rect -3190 -15192 -3170 -15128
rect -9469 -15208 -3170 -15192
rect -9469 -15272 -3254 -15208
rect -3190 -15272 -3170 -15208
rect -9469 -15288 -3170 -15272
rect -9469 -15352 -3254 -15288
rect -3190 -15352 -3170 -15288
rect -9469 -15368 -3170 -15352
rect -9469 -15432 -3254 -15368
rect -3190 -15432 -3170 -15368
rect -9469 -15448 -3170 -15432
rect -9469 -15512 -3254 -15448
rect -3190 -15512 -3170 -15448
rect -9469 -15528 -3170 -15512
rect -9469 -15592 -3254 -15528
rect -3190 -15592 -3170 -15528
rect -9469 -15608 -3170 -15592
rect -9469 -15672 -3254 -15608
rect -3190 -15672 -3170 -15608
rect -9469 -15700 -3170 -15672
rect -3150 -9528 3149 -9500
rect -3150 -9592 3065 -9528
rect 3129 -9592 3149 -9528
rect -3150 -9608 3149 -9592
rect -3150 -9672 3065 -9608
rect 3129 -9672 3149 -9608
rect -3150 -9688 3149 -9672
rect -3150 -9752 3065 -9688
rect 3129 -9752 3149 -9688
rect -3150 -9768 3149 -9752
rect -3150 -9832 3065 -9768
rect 3129 -9832 3149 -9768
rect -3150 -9848 3149 -9832
rect -3150 -9912 3065 -9848
rect 3129 -9912 3149 -9848
rect -3150 -9928 3149 -9912
rect -3150 -9992 3065 -9928
rect 3129 -9992 3149 -9928
rect -3150 -10008 3149 -9992
rect -3150 -10072 3065 -10008
rect 3129 -10072 3149 -10008
rect -3150 -10088 3149 -10072
rect -3150 -10152 3065 -10088
rect 3129 -10152 3149 -10088
rect -3150 -10168 3149 -10152
rect -3150 -10232 3065 -10168
rect 3129 -10232 3149 -10168
rect -3150 -10248 3149 -10232
rect -3150 -10312 3065 -10248
rect 3129 -10312 3149 -10248
rect -3150 -10328 3149 -10312
rect -3150 -10392 3065 -10328
rect 3129 -10392 3149 -10328
rect -3150 -10408 3149 -10392
rect -3150 -10472 3065 -10408
rect 3129 -10472 3149 -10408
rect -3150 -10488 3149 -10472
rect -3150 -10552 3065 -10488
rect 3129 -10552 3149 -10488
rect -3150 -10568 3149 -10552
rect -3150 -10632 3065 -10568
rect 3129 -10632 3149 -10568
rect -3150 -10648 3149 -10632
rect -3150 -10712 3065 -10648
rect 3129 -10712 3149 -10648
rect -3150 -10728 3149 -10712
rect -3150 -10792 3065 -10728
rect 3129 -10792 3149 -10728
rect -3150 -10808 3149 -10792
rect -3150 -10872 3065 -10808
rect 3129 -10872 3149 -10808
rect -3150 -10888 3149 -10872
rect -3150 -10952 3065 -10888
rect 3129 -10952 3149 -10888
rect -3150 -10968 3149 -10952
rect -3150 -11032 3065 -10968
rect 3129 -11032 3149 -10968
rect -3150 -11048 3149 -11032
rect -3150 -11112 3065 -11048
rect 3129 -11112 3149 -11048
rect -3150 -11128 3149 -11112
rect -3150 -11192 3065 -11128
rect 3129 -11192 3149 -11128
rect -3150 -11208 3149 -11192
rect -3150 -11272 3065 -11208
rect 3129 -11272 3149 -11208
rect -3150 -11288 3149 -11272
rect -3150 -11352 3065 -11288
rect 3129 -11352 3149 -11288
rect -3150 -11368 3149 -11352
rect -3150 -11432 3065 -11368
rect 3129 -11432 3149 -11368
rect -3150 -11448 3149 -11432
rect -3150 -11512 3065 -11448
rect 3129 -11512 3149 -11448
rect -3150 -11528 3149 -11512
rect -3150 -11592 3065 -11528
rect 3129 -11592 3149 -11528
rect -3150 -11608 3149 -11592
rect -3150 -11672 3065 -11608
rect 3129 -11672 3149 -11608
rect -3150 -11688 3149 -11672
rect -3150 -11752 3065 -11688
rect 3129 -11752 3149 -11688
rect -3150 -11768 3149 -11752
rect -3150 -11832 3065 -11768
rect 3129 -11832 3149 -11768
rect -3150 -11848 3149 -11832
rect -3150 -11912 3065 -11848
rect 3129 -11912 3149 -11848
rect -3150 -11928 3149 -11912
rect -3150 -11992 3065 -11928
rect 3129 -11992 3149 -11928
rect -3150 -12008 3149 -11992
rect -3150 -12072 3065 -12008
rect 3129 -12072 3149 -12008
rect -3150 -12088 3149 -12072
rect -3150 -12152 3065 -12088
rect 3129 -12152 3149 -12088
rect -3150 -12168 3149 -12152
rect -3150 -12232 3065 -12168
rect 3129 -12232 3149 -12168
rect -3150 -12248 3149 -12232
rect -3150 -12312 3065 -12248
rect 3129 -12312 3149 -12248
rect -3150 -12328 3149 -12312
rect -3150 -12392 3065 -12328
rect 3129 -12392 3149 -12328
rect -3150 -12408 3149 -12392
rect -3150 -12472 3065 -12408
rect 3129 -12472 3149 -12408
rect -3150 -12488 3149 -12472
rect -3150 -12552 3065 -12488
rect 3129 -12552 3149 -12488
rect -3150 -12568 3149 -12552
rect -3150 -12632 3065 -12568
rect 3129 -12632 3149 -12568
rect -3150 -12648 3149 -12632
rect -3150 -12712 3065 -12648
rect 3129 -12712 3149 -12648
rect -3150 -12728 3149 -12712
rect -3150 -12792 3065 -12728
rect 3129 -12792 3149 -12728
rect -3150 -12808 3149 -12792
rect -3150 -12872 3065 -12808
rect 3129 -12872 3149 -12808
rect -3150 -12888 3149 -12872
rect -3150 -12952 3065 -12888
rect 3129 -12952 3149 -12888
rect -3150 -12968 3149 -12952
rect -3150 -13032 3065 -12968
rect 3129 -13032 3149 -12968
rect -3150 -13048 3149 -13032
rect -3150 -13112 3065 -13048
rect 3129 -13112 3149 -13048
rect -3150 -13128 3149 -13112
rect -3150 -13192 3065 -13128
rect 3129 -13192 3149 -13128
rect -3150 -13208 3149 -13192
rect -3150 -13272 3065 -13208
rect 3129 -13272 3149 -13208
rect -3150 -13288 3149 -13272
rect -3150 -13352 3065 -13288
rect 3129 -13352 3149 -13288
rect -3150 -13368 3149 -13352
rect -3150 -13432 3065 -13368
rect 3129 -13432 3149 -13368
rect -3150 -13448 3149 -13432
rect -3150 -13512 3065 -13448
rect 3129 -13512 3149 -13448
rect -3150 -13528 3149 -13512
rect -3150 -13592 3065 -13528
rect 3129 -13592 3149 -13528
rect -3150 -13608 3149 -13592
rect -3150 -13672 3065 -13608
rect 3129 -13672 3149 -13608
rect -3150 -13688 3149 -13672
rect -3150 -13752 3065 -13688
rect 3129 -13752 3149 -13688
rect -3150 -13768 3149 -13752
rect -3150 -13832 3065 -13768
rect 3129 -13832 3149 -13768
rect -3150 -13848 3149 -13832
rect -3150 -13912 3065 -13848
rect 3129 -13912 3149 -13848
rect -3150 -13928 3149 -13912
rect -3150 -13992 3065 -13928
rect 3129 -13992 3149 -13928
rect -3150 -14008 3149 -13992
rect -3150 -14072 3065 -14008
rect 3129 -14072 3149 -14008
rect -3150 -14088 3149 -14072
rect -3150 -14152 3065 -14088
rect 3129 -14152 3149 -14088
rect -3150 -14168 3149 -14152
rect -3150 -14232 3065 -14168
rect 3129 -14232 3149 -14168
rect -3150 -14248 3149 -14232
rect -3150 -14312 3065 -14248
rect 3129 -14312 3149 -14248
rect -3150 -14328 3149 -14312
rect -3150 -14392 3065 -14328
rect 3129 -14392 3149 -14328
rect -3150 -14408 3149 -14392
rect -3150 -14472 3065 -14408
rect 3129 -14472 3149 -14408
rect -3150 -14488 3149 -14472
rect -3150 -14552 3065 -14488
rect 3129 -14552 3149 -14488
rect -3150 -14568 3149 -14552
rect -3150 -14632 3065 -14568
rect 3129 -14632 3149 -14568
rect -3150 -14648 3149 -14632
rect -3150 -14712 3065 -14648
rect 3129 -14712 3149 -14648
rect -3150 -14728 3149 -14712
rect -3150 -14792 3065 -14728
rect 3129 -14792 3149 -14728
rect -3150 -14808 3149 -14792
rect -3150 -14872 3065 -14808
rect 3129 -14872 3149 -14808
rect -3150 -14888 3149 -14872
rect -3150 -14952 3065 -14888
rect 3129 -14952 3149 -14888
rect -3150 -14968 3149 -14952
rect -3150 -15032 3065 -14968
rect 3129 -15032 3149 -14968
rect -3150 -15048 3149 -15032
rect -3150 -15112 3065 -15048
rect 3129 -15112 3149 -15048
rect -3150 -15128 3149 -15112
rect -3150 -15192 3065 -15128
rect 3129 -15192 3149 -15128
rect -3150 -15208 3149 -15192
rect -3150 -15272 3065 -15208
rect 3129 -15272 3149 -15208
rect -3150 -15288 3149 -15272
rect -3150 -15352 3065 -15288
rect 3129 -15352 3149 -15288
rect -3150 -15368 3149 -15352
rect -3150 -15432 3065 -15368
rect 3129 -15432 3149 -15368
rect -3150 -15448 3149 -15432
rect -3150 -15512 3065 -15448
rect 3129 -15512 3149 -15448
rect -3150 -15528 3149 -15512
rect -3150 -15592 3065 -15528
rect 3129 -15592 3149 -15528
rect -3150 -15608 3149 -15592
rect -3150 -15672 3065 -15608
rect 3129 -15672 3149 -15608
rect -3150 -15700 3149 -15672
rect 3169 -9528 9468 -9500
rect 3169 -9592 9384 -9528
rect 9448 -9592 9468 -9528
rect 3169 -9608 9468 -9592
rect 3169 -9672 9384 -9608
rect 9448 -9672 9468 -9608
rect 3169 -9688 9468 -9672
rect 3169 -9752 9384 -9688
rect 9448 -9752 9468 -9688
rect 3169 -9768 9468 -9752
rect 3169 -9832 9384 -9768
rect 9448 -9832 9468 -9768
rect 3169 -9848 9468 -9832
rect 3169 -9912 9384 -9848
rect 9448 -9912 9468 -9848
rect 3169 -9928 9468 -9912
rect 3169 -9992 9384 -9928
rect 9448 -9992 9468 -9928
rect 3169 -10008 9468 -9992
rect 3169 -10072 9384 -10008
rect 9448 -10072 9468 -10008
rect 3169 -10088 9468 -10072
rect 3169 -10152 9384 -10088
rect 9448 -10152 9468 -10088
rect 3169 -10168 9468 -10152
rect 3169 -10232 9384 -10168
rect 9448 -10232 9468 -10168
rect 3169 -10248 9468 -10232
rect 3169 -10312 9384 -10248
rect 9448 -10312 9468 -10248
rect 3169 -10328 9468 -10312
rect 3169 -10392 9384 -10328
rect 9448 -10392 9468 -10328
rect 3169 -10408 9468 -10392
rect 3169 -10472 9384 -10408
rect 9448 -10472 9468 -10408
rect 3169 -10488 9468 -10472
rect 3169 -10552 9384 -10488
rect 9448 -10552 9468 -10488
rect 3169 -10568 9468 -10552
rect 3169 -10632 9384 -10568
rect 9448 -10632 9468 -10568
rect 3169 -10648 9468 -10632
rect 3169 -10712 9384 -10648
rect 9448 -10712 9468 -10648
rect 3169 -10728 9468 -10712
rect 3169 -10792 9384 -10728
rect 9448 -10792 9468 -10728
rect 3169 -10808 9468 -10792
rect 3169 -10872 9384 -10808
rect 9448 -10872 9468 -10808
rect 3169 -10888 9468 -10872
rect 3169 -10952 9384 -10888
rect 9448 -10952 9468 -10888
rect 3169 -10968 9468 -10952
rect 3169 -11032 9384 -10968
rect 9448 -11032 9468 -10968
rect 3169 -11048 9468 -11032
rect 3169 -11112 9384 -11048
rect 9448 -11112 9468 -11048
rect 3169 -11128 9468 -11112
rect 3169 -11192 9384 -11128
rect 9448 -11192 9468 -11128
rect 3169 -11208 9468 -11192
rect 3169 -11272 9384 -11208
rect 9448 -11272 9468 -11208
rect 3169 -11288 9468 -11272
rect 3169 -11352 9384 -11288
rect 9448 -11352 9468 -11288
rect 3169 -11368 9468 -11352
rect 3169 -11432 9384 -11368
rect 9448 -11432 9468 -11368
rect 3169 -11448 9468 -11432
rect 3169 -11512 9384 -11448
rect 9448 -11512 9468 -11448
rect 3169 -11528 9468 -11512
rect 3169 -11592 9384 -11528
rect 9448 -11592 9468 -11528
rect 3169 -11608 9468 -11592
rect 3169 -11672 9384 -11608
rect 9448 -11672 9468 -11608
rect 3169 -11688 9468 -11672
rect 3169 -11752 9384 -11688
rect 9448 -11752 9468 -11688
rect 3169 -11768 9468 -11752
rect 3169 -11832 9384 -11768
rect 9448 -11832 9468 -11768
rect 3169 -11848 9468 -11832
rect 3169 -11912 9384 -11848
rect 9448 -11912 9468 -11848
rect 3169 -11928 9468 -11912
rect 3169 -11992 9384 -11928
rect 9448 -11992 9468 -11928
rect 3169 -12008 9468 -11992
rect 3169 -12072 9384 -12008
rect 9448 -12072 9468 -12008
rect 3169 -12088 9468 -12072
rect 3169 -12152 9384 -12088
rect 9448 -12152 9468 -12088
rect 3169 -12168 9468 -12152
rect 3169 -12232 9384 -12168
rect 9448 -12232 9468 -12168
rect 3169 -12248 9468 -12232
rect 3169 -12312 9384 -12248
rect 9448 -12312 9468 -12248
rect 3169 -12328 9468 -12312
rect 3169 -12392 9384 -12328
rect 9448 -12392 9468 -12328
rect 3169 -12408 9468 -12392
rect 3169 -12472 9384 -12408
rect 9448 -12472 9468 -12408
rect 3169 -12488 9468 -12472
rect 3169 -12552 9384 -12488
rect 9448 -12552 9468 -12488
rect 3169 -12568 9468 -12552
rect 3169 -12632 9384 -12568
rect 9448 -12632 9468 -12568
rect 3169 -12648 9468 -12632
rect 3169 -12712 9384 -12648
rect 9448 -12712 9468 -12648
rect 3169 -12728 9468 -12712
rect 3169 -12792 9384 -12728
rect 9448 -12792 9468 -12728
rect 3169 -12808 9468 -12792
rect 3169 -12872 9384 -12808
rect 9448 -12872 9468 -12808
rect 3169 -12888 9468 -12872
rect 3169 -12952 9384 -12888
rect 9448 -12952 9468 -12888
rect 3169 -12968 9468 -12952
rect 3169 -13032 9384 -12968
rect 9448 -13032 9468 -12968
rect 3169 -13048 9468 -13032
rect 3169 -13112 9384 -13048
rect 9448 -13112 9468 -13048
rect 3169 -13128 9468 -13112
rect 3169 -13192 9384 -13128
rect 9448 -13192 9468 -13128
rect 3169 -13208 9468 -13192
rect 3169 -13272 9384 -13208
rect 9448 -13272 9468 -13208
rect 3169 -13288 9468 -13272
rect 3169 -13352 9384 -13288
rect 9448 -13352 9468 -13288
rect 3169 -13368 9468 -13352
rect 3169 -13432 9384 -13368
rect 9448 -13432 9468 -13368
rect 3169 -13448 9468 -13432
rect 3169 -13512 9384 -13448
rect 9448 -13512 9468 -13448
rect 3169 -13528 9468 -13512
rect 3169 -13592 9384 -13528
rect 9448 -13592 9468 -13528
rect 3169 -13608 9468 -13592
rect 3169 -13672 9384 -13608
rect 9448 -13672 9468 -13608
rect 3169 -13688 9468 -13672
rect 3169 -13752 9384 -13688
rect 9448 -13752 9468 -13688
rect 3169 -13768 9468 -13752
rect 3169 -13832 9384 -13768
rect 9448 -13832 9468 -13768
rect 3169 -13848 9468 -13832
rect 3169 -13912 9384 -13848
rect 9448 -13912 9468 -13848
rect 3169 -13928 9468 -13912
rect 3169 -13992 9384 -13928
rect 9448 -13992 9468 -13928
rect 3169 -14008 9468 -13992
rect 3169 -14072 9384 -14008
rect 9448 -14072 9468 -14008
rect 3169 -14088 9468 -14072
rect 3169 -14152 9384 -14088
rect 9448 -14152 9468 -14088
rect 3169 -14168 9468 -14152
rect 3169 -14232 9384 -14168
rect 9448 -14232 9468 -14168
rect 3169 -14248 9468 -14232
rect 3169 -14312 9384 -14248
rect 9448 -14312 9468 -14248
rect 3169 -14328 9468 -14312
rect 3169 -14392 9384 -14328
rect 9448 -14392 9468 -14328
rect 3169 -14408 9468 -14392
rect 3169 -14472 9384 -14408
rect 9448 -14472 9468 -14408
rect 3169 -14488 9468 -14472
rect 3169 -14552 9384 -14488
rect 9448 -14552 9468 -14488
rect 3169 -14568 9468 -14552
rect 3169 -14632 9384 -14568
rect 9448 -14632 9468 -14568
rect 3169 -14648 9468 -14632
rect 3169 -14712 9384 -14648
rect 9448 -14712 9468 -14648
rect 3169 -14728 9468 -14712
rect 3169 -14792 9384 -14728
rect 9448 -14792 9468 -14728
rect 3169 -14808 9468 -14792
rect 3169 -14872 9384 -14808
rect 9448 -14872 9468 -14808
rect 3169 -14888 9468 -14872
rect 3169 -14952 9384 -14888
rect 9448 -14952 9468 -14888
rect 3169 -14968 9468 -14952
rect 3169 -15032 9384 -14968
rect 9448 -15032 9468 -14968
rect 3169 -15048 9468 -15032
rect 3169 -15112 9384 -15048
rect 9448 -15112 9468 -15048
rect 3169 -15128 9468 -15112
rect 3169 -15192 9384 -15128
rect 9448 -15192 9468 -15128
rect 3169 -15208 9468 -15192
rect 3169 -15272 9384 -15208
rect 9448 -15272 9468 -15208
rect 3169 -15288 9468 -15272
rect 3169 -15352 9384 -15288
rect 9448 -15352 9468 -15288
rect 3169 -15368 9468 -15352
rect 3169 -15432 9384 -15368
rect 9448 -15432 9468 -15368
rect 3169 -15448 9468 -15432
rect 3169 -15512 9384 -15448
rect 9448 -15512 9468 -15448
rect 3169 -15528 9468 -15512
rect 3169 -15592 9384 -15528
rect 9448 -15592 9468 -15528
rect 3169 -15608 9468 -15592
rect 3169 -15672 9384 -15608
rect 9448 -15672 9468 -15608
rect 3169 -15700 9468 -15672
rect 9488 -9528 15787 -9500
rect 9488 -9592 15703 -9528
rect 15767 -9592 15787 -9528
rect 9488 -9608 15787 -9592
rect 9488 -9672 15703 -9608
rect 15767 -9672 15787 -9608
rect 9488 -9688 15787 -9672
rect 9488 -9752 15703 -9688
rect 15767 -9752 15787 -9688
rect 9488 -9768 15787 -9752
rect 9488 -9832 15703 -9768
rect 15767 -9832 15787 -9768
rect 9488 -9848 15787 -9832
rect 9488 -9912 15703 -9848
rect 15767 -9912 15787 -9848
rect 9488 -9928 15787 -9912
rect 9488 -9992 15703 -9928
rect 15767 -9992 15787 -9928
rect 9488 -10008 15787 -9992
rect 9488 -10072 15703 -10008
rect 15767 -10072 15787 -10008
rect 9488 -10088 15787 -10072
rect 9488 -10152 15703 -10088
rect 15767 -10152 15787 -10088
rect 9488 -10168 15787 -10152
rect 9488 -10232 15703 -10168
rect 15767 -10232 15787 -10168
rect 9488 -10248 15787 -10232
rect 9488 -10312 15703 -10248
rect 15767 -10312 15787 -10248
rect 9488 -10328 15787 -10312
rect 9488 -10392 15703 -10328
rect 15767 -10392 15787 -10328
rect 9488 -10408 15787 -10392
rect 9488 -10472 15703 -10408
rect 15767 -10472 15787 -10408
rect 9488 -10488 15787 -10472
rect 9488 -10552 15703 -10488
rect 15767 -10552 15787 -10488
rect 9488 -10568 15787 -10552
rect 9488 -10632 15703 -10568
rect 15767 -10632 15787 -10568
rect 9488 -10648 15787 -10632
rect 9488 -10712 15703 -10648
rect 15767 -10712 15787 -10648
rect 9488 -10728 15787 -10712
rect 9488 -10792 15703 -10728
rect 15767 -10792 15787 -10728
rect 9488 -10808 15787 -10792
rect 9488 -10872 15703 -10808
rect 15767 -10872 15787 -10808
rect 9488 -10888 15787 -10872
rect 9488 -10952 15703 -10888
rect 15767 -10952 15787 -10888
rect 9488 -10968 15787 -10952
rect 9488 -11032 15703 -10968
rect 15767 -11032 15787 -10968
rect 9488 -11048 15787 -11032
rect 9488 -11112 15703 -11048
rect 15767 -11112 15787 -11048
rect 9488 -11128 15787 -11112
rect 9488 -11192 15703 -11128
rect 15767 -11192 15787 -11128
rect 9488 -11208 15787 -11192
rect 9488 -11272 15703 -11208
rect 15767 -11272 15787 -11208
rect 9488 -11288 15787 -11272
rect 9488 -11352 15703 -11288
rect 15767 -11352 15787 -11288
rect 9488 -11368 15787 -11352
rect 9488 -11432 15703 -11368
rect 15767 -11432 15787 -11368
rect 9488 -11448 15787 -11432
rect 9488 -11512 15703 -11448
rect 15767 -11512 15787 -11448
rect 9488 -11528 15787 -11512
rect 9488 -11592 15703 -11528
rect 15767 -11592 15787 -11528
rect 9488 -11608 15787 -11592
rect 9488 -11672 15703 -11608
rect 15767 -11672 15787 -11608
rect 9488 -11688 15787 -11672
rect 9488 -11752 15703 -11688
rect 15767 -11752 15787 -11688
rect 9488 -11768 15787 -11752
rect 9488 -11832 15703 -11768
rect 15767 -11832 15787 -11768
rect 9488 -11848 15787 -11832
rect 9488 -11912 15703 -11848
rect 15767 -11912 15787 -11848
rect 9488 -11928 15787 -11912
rect 9488 -11992 15703 -11928
rect 15767 -11992 15787 -11928
rect 9488 -12008 15787 -11992
rect 9488 -12072 15703 -12008
rect 15767 -12072 15787 -12008
rect 9488 -12088 15787 -12072
rect 9488 -12152 15703 -12088
rect 15767 -12152 15787 -12088
rect 9488 -12168 15787 -12152
rect 9488 -12232 15703 -12168
rect 15767 -12232 15787 -12168
rect 9488 -12248 15787 -12232
rect 9488 -12312 15703 -12248
rect 15767 -12312 15787 -12248
rect 9488 -12328 15787 -12312
rect 9488 -12392 15703 -12328
rect 15767 -12392 15787 -12328
rect 9488 -12408 15787 -12392
rect 9488 -12472 15703 -12408
rect 15767 -12472 15787 -12408
rect 9488 -12488 15787 -12472
rect 9488 -12552 15703 -12488
rect 15767 -12552 15787 -12488
rect 9488 -12568 15787 -12552
rect 9488 -12632 15703 -12568
rect 15767 -12632 15787 -12568
rect 9488 -12648 15787 -12632
rect 9488 -12712 15703 -12648
rect 15767 -12712 15787 -12648
rect 9488 -12728 15787 -12712
rect 9488 -12792 15703 -12728
rect 15767 -12792 15787 -12728
rect 9488 -12808 15787 -12792
rect 9488 -12872 15703 -12808
rect 15767 -12872 15787 -12808
rect 9488 -12888 15787 -12872
rect 9488 -12952 15703 -12888
rect 15767 -12952 15787 -12888
rect 9488 -12968 15787 -12952
rect 9488 -13032 15703 -12968
rect 15767 -13032 15787 -12968
rect 9488 -13048 15787 -13032
rect 9488 -13112 15703 -13048
rect 15767 -13112 15787 -13048
rect 9488 -13128 15787 -13112
rect 9488 -13192 15703 -13128
rect 15767 -13192 15787 -13128
rect 9488 -13208 15787 -13192
rect 9488 -13272 15703 -13208
rect 15767 -13272 15787 -13208
rect 9488 -13288 15787 -13272
rect 9488 -13352 15703 -13288
rect 15767 -13352 15787 -13288
rect 9488 -13368 15787 -13352
rect 9488 -13432 15703 -13368
rect 15767 -13432 15787 -13368
rect 9488 -13448 15787 -13432
rect 9488 -13512 15703 -13448
rect 15767 -13512 15787 -13448
rect 9488 -13528 15787 -13512
rect 9488 -13592 15703 -13528
rect 15767 -13592 15787 -13528
rect 9488 -13608 15787 -13592
rect 9488 -13672 15703 -13608
rect 15767 -13672 15787 -13608
rect 9488 -13688 15787 -13672
rect 9488 -13752 15703 -13688
rect 15767 -13752 15787 -13688
rect 9488 -13768 15787 -13752
rect 9488 -13832 15703 -13768
rect 15767 -13832 15787 -13768
rect 9488 -13848 15787 -13832
rect 9488 -13912 15703 -13848
rect 15767 -13912 15787 -13848
rect 9488 -13928 15787 -13912
rect 9488 -13992 15703 -13928
rect 15767 -13992 15787 -13928
rect 9488 -14008 15787 -13992
rect 9488 -14072 15703 -14008
rect 15767 -14072 15787 -14008
rect 9488 -14088 15787 -14072
rect 9488 -14152 15703 -14088
rect 15767 -14152 15787 -14088
rect 9488 -14168 15787 -14152
rect 9488 -14232 15703 -14168
rect 15767 -14232 15787 -14168
rect 9488 -14248 15787 -14232
rect 9488 -14312 15703 -14248
rect 15767 -14312 15787 -14248
rect 9488 -14328 15787 -14312
rect 9488 -14392 15703 -14328
rect 15767 -14392 15787 -14328
rect 9488 -14408 15787 -14392
rect 9488 -14472 15703 -14408
rect 15767 -14472 15787 -14408
rect 9488 -14488 15787 -14472
rect 9488 -14552 15703 -14488
rect 15767 -14552 15787 -14488
rect 9488 -14568 15787 -14552
rect 9488 -14632 15703 -14568
rect 15767 -14632 15787 -14568
rect 9488 -14648 15787 -14632
rect 9488 -14712 15703 -14648
rect 15767 -14712 15787 -14648
rect 9488 -14728 15787 -14712
rect 9488 -14792 15703 -14728
rect 15767 -14792 15787 -14728
rect 9488 -14808 15787 -14792
rect 9488 -14872 15703 -14808
rect 15767 -14872 15787 -14808
rect 9488 -14888 15787 -14872
rect 9488 -14952 15703 -14888
rect 15767 -14952 15787 -14888
rect 9488 -14968 15787 -14952
rect 9488 -15032 15703 -14968
rect 15767 -15032 15787 -14968
rect 9488 -15048 15787 -15032
rect 9488 -15112 15703 -15048
rect 15767 -15112 15787 -15048
rect 9488 -15128 15787 -15112
rect 9488 -15192 15703 -15128
rect 15767 -15192 15787 -15128
rect 9488 -15208 15787 -15192
rect 9488 -15272 15703 -15208
rect 15767 -15272 15787 -15208
rect 9488 -15288 15787 -15272
rect 9488 -15352 15703 -15288
rect 15767 -15352 15787 -15288
rect 9488 -15368 15787 -15352
rect 9488 -15432 15703 -15368
rect 15767 -15432 15787 -15368
rect 9488 -15448 15787 -15432
rect 9488 -15512 15703 -15448
rect 15767 -15512 15787 -15448
rect 9488 -15528 15787 -15512
rect 9488 -15592 15703 -15528
rect 15767 -15592 15787 -15528
rect 9488 -15608 15787 -15592
rect 9488 -15672 15703 -15608
rect 15767 -15672 15787 -15608
rect 9488 -15700 15787 -15672
rect 15807 -9528 22106 -9500
rect 15807 -9592 22022 -9528
rect 22086 -9592 22106 -9528
rect 15807 -9608 22106 -9592
rect 15807 -9672 22022 -9608
rect 22086 -9672 22106 -9608
rect 15807 -9688 22106 -9672
rect 15807 -9752 22022 -9688
rect 22086 -9752 22106 -9688
rect 15807 -9768 22106 -9752
rect 15807 -9832 22022 -9768
rect 22086 -9832 22106 -9768
rect 15807 -9848 22106 -9832
rect 15807 -9912 22022 -9848
rect 22086 -9912 22106 -9848
rect 15807 -9928 22106 -9912
rect 15807 -9992 22022 -9928
rect 22086 -9992 22106 -9928
rect 15807 -10008 22106 -9992
rect 15807 -10072 22022 -10008
rect 22086 -10072 22106 -10008
rect 15807 -10088 22106 -10072
rect 15807 -10152 22022 -10088
rect 22086 -10152 22106 -10088
rect 15807 -10168 22106 -10152
rect 15807 -10232 22022 -10168
rect 22086 -10232 22106 -10168
rect 15807 -10248 22106 -10232
rect 15807 -10312 22022 -10248
rect 22086 -10312 22106 -10248
rect 15807 -10328 22106 -10312
rect 15807 -10392 22022 -10328
rect 22086 -10392 22106 -10328
rect 15807 -10408 22106 -10392
rect 15807 -10472 22022 -10408
rect 22086 -10472 22106 -10408
rect 15807 -10488 22106 -10472
rect 15807 -10552 22022 -10488
rect 22086 -10552 22106 -10488
rect 15807 -10568 22106 -10552
rect 15807 -10632 22022 -10568
rect 22086 -10632 22106 -10568
rect 15807 -10648 22106 -10632
rect 15807 -10712 22022 -10648
rect 22086 -10712 22106 -10648
rect 15807 -10728 22106 -10712
rect 15807 -10792 22022 -10728
rect 22086 -10792 22106 -10728
rect 15807 -10808 22106 -10792
rect 15807 -10872 22022 -10808
rect 22086 -10872 22106 -10808
rect 15807 -10888 22106 -10872
rect 15807 -10952 22022 -10888
rect 22086 -10952 22106 -10888
rect 15807 -10968 22106 -10952
rect 15807 -11032 22022 -10968
rect 22086 -11032 22106 -10968
rect 15807 -11048 22106 -11032
rect 15807 -11112 22022 -11048
rect 22086 -11112 22106 -11048
rect 15807 -11128 22106 -11112
rect 15807 -11192 22022 -11128
rect 22086 -11192 22106 -11128
rect 15807 -11208 22106 -11192
rect 15807 -11272 22022 -11208
rect 22086 -11272 22106 -11208
rect 15807 -11288 22106 -11272
rect 15807 -11352 22022 -11288
rect 22086 -11352 22106 -11288
rect 15807 -11368 22106 -11352
rect 15807 -11432 22022 -11368
rect 22086 -11432 22106 -11368
rect 15807 -11448 22106 -11432
rect 15807 -11512 22022 -11448
rect 22086 -11512 22106 -11448
rect 15807 -11528 22106 -11512
rect 15807 -11592 22022 -11528
rect 22086 -11592 22106 -11528
rect 15807 -11608 22106 -11592
rect 15807 -11672 22022 -11608
rect 22086 -11672 22106 -11608
rect 15807 -11688 22106 -11672
rect 15807 -11752 22022 -11688
rect 22086 -11752 22106 -11688
rect 15807 -11768 22106 -11752
rect 15807 -11832 22022 -11768
rect 22086 -11832 22106 -11768
rect 15807 -11848 22106 -11832
rect 15807 -11912 22022 -11848
rect 22086 -11912 22106 -11848
rect 15807 -11928 22106 -11912
rect 15807 -11992 22022 -11928
rect 22086 -11992 22106 -11928
rect 15807 -12008 22106 -11992
rect 15807 -12072 22022 -12008
rect 22086 -12072 22106 -12008
rect 15807 -12088 22106 -12072
rect 15807 -12152 22022 -12088
rect 22086 -12152 22106 -12088
rect 15807 -12168 22106 -12152
rect 15807 -12232 22022 -12168
rect 22086 -12232 22106 -12168
rect 15807 -12248 22106 -12232
rect 15807 -12312 22022 -12248
rect 22086 -12312 22106 -12248
rect 15807 -12328 22106 -12312
rect 15807 -12392 22022 -12328
rect 22086 -12392 22106 -12328
rect 15807 -12408 22106 -12392
rect 15807 -12472 22022 -12408
rect 22086 -12472 22106 -12408
rect 15807 -12488 22106 -12472
rect 15807 -12552 22022 -12488
rect 22086 -12552 22106 -12488
rect 15807 -12568 22106 -12552
rect 15807 -12632 22022 -12568
rect 22086 -12632 22106 -12568
rect 15807 -12648 22106 -12632
rect 15807 -12712 22022 -12648
rect 22086 -12712 22106 -12648
rect 15807 -12728 22106 -12712
rect 15807 -12792 22022 -12728
rect 22086 -12792 22106 -12728
rect 15807 -12808 22106 -12792
rect 15807 -12872 22022 -12808
rect 22086 -12872 22106 -12808
rect 15807 -12888 22106 -12872
rect 15807 -12952 22022 -12888
rect 22086 -12952 22106 -12888
rect 15807 -12968 22106 -12952
rect 15807 -13032 22022 -12968
rect 22086 -13032 22106 -12968
rect 15807 -13048 22106 -13032
rect 15807 -13112 22022 -13048
rect 22086 -13112 22106 -13048
rect 15807 -13128 22106 -13112
rect 15807 -13192 22022 -13128
rect 22086 -13192 22106 -13128
rect 15807 -13208 22106 -13192
rect 15807 -13272 22022 -13208
rect 22086 -13272 22106 -13208
rect 15807 -13288 22106 -13272
rect 15807 -13352 22022 -13288
rect 22086 -13352 22106 -13288
rect 15807 -13368 22106 -13352
rect 15807 -13432 22022 -13368
rect 22086 -13432 22106 -13368
rect 15807 -13448 22106 -13432
rect 15807 -13512 22022 -13448
rect 22086 -13512 22106 -13448
rect 15807 -13528 22106 -13512
rect 15807 -13592 22022 -13528
rect 22086 -13592 22106 -13528
rect 15807 -13608 22106 -13592
rect 15807 -13672 22022 -13608
rect 22086 -13672 22106 -13608
rect 15807 -13688 22106 -13672
rect 15807 -13752 22022 -13688
rect 22086 -13752 22106 -13688
rect 15807 -13768 22106 -13752
rect 15807 -13832 22022 -13768
rect 22086 -13832 22106 -13768
rect 15807 -13848 22106 -13832
rect 15807 -13912 22022 -13848
rect 22086 -13912 22106 -13848
rect 15807 -13928 22106 -13912
rect 15807 -13992 22022 -13928
rect 22086 -13992 22106 -13928
rect 15807 -14008 22106 -13992
rect 15807 -14072 22022 -14008
rect 22086 -14072 22106 -14008
rect 15807 -14088 22106 -14072
rect 15807 -14152 22022 -14088
rect 22086 -14152 22106 -14088
rect 15807 -14168 22106 -14152
rect 15807 -14232 22022 -14168
rect 22086 -14232 22106 -14168
rect 15807 -14248 22106 -14232
rect 15807 -14312 22022 -14248
rect 22086 -14312 22106 -14248
rect 15807 -14328 22106 -14312
rect 15807 -14392 22022 -14328
rect 22086 -14392 22106 -14328
rect 15807 -14408 22106 -14392
rect 15807 -14472 22022 -14408
rect 22086 -14472 22106 -14408
rect 15807 -14488 22106 -14472
rect 15807 -14552 22022 -14488
rect 22086 -14552 22106 -14488
rect 15807 -14568 22106 -14552
rect 15807 -14632 22022 -14568
rect 22086 -14632 22106 -14568
rect 15807 -14648 22106 -14632
rect 15807 -14712 22022 -14648
rect 22086 -14712 22106 -14648
rect 15807 -14728 22106 -14712
rect 15807 -14792 22022 -14728
rect 22086 -14792 22106 -14728
rect 15807 -14808 22106 -14792
rect 15807 -14872 22022 -14808
rect 22086 -14872 22106 -14808
rect 15807 -14888 22106 -14872
rect 15807 -14952 22022 -14888
rect 22086 -14952 22106 -14888
rect 15807 -14968 22106 -14952
rect 15807 -15032 22022 -14968
rect 22086 -15032 22106 -14968
rect 15807 -15048 22106 -15032
rect 15807 -15112 22022 -15048
rect 22086 -15112 22106 -15048
rect 15807 -15128 22106 -15112
rect 15807 -15192 22022 -15128
rect 22086 -15192 22106 -15128
rect 15807 -15208 22106 -15192
rect 15807 -15272 22022 -15208
rect 22086 -15272 22106 -15208
rect 15807 -15288 22106 -15272
rect 15807 -15352 22022 -15288
rect 22086 -15352 22106 -15288
rect 15807 -15368 22106 -15352
rect 15807 -15432 22022 -15368
rect 22086 -15432 22106 -15368
rect 15807 -15448 22106 -15432
rect 15807 -15512 22022 -15448
rect 22086 -15512 22106 -15448
rect 15807 -15528 22106 -15512
rect 15807 -15592 22022 -15528
rect 22086 -15592 22106 -15528
rect 15807 -15608 22106 -15592
rect 15807 -15672 22022 -15608
rect 22086 -15672 22106 -15608
rect 15807 -15700 22106 -15672
rect 22126 -9528 28425 -9500
rect 22126 -9592 28341 -9528
rect 28405 -9592 28425 -9528
rect 22126 -9608 28425 -9592
rect 22126 -9672 28341 -9608
rect 28405 -9672 28425 -9608
rect 22126 -9688 28425 -9672
rect 22126 -9752 28341 -9688
rect 28405 -9752 28425 -9688
rect 22126 -9768 28425 -9752
rect 22126 -9832 28341 -9768
rect 28405 -9832 28425 -9768
rect 22126 -9848 28425 -9832
rect 22126 -9912 28341 -9848
rect 28405 -9912 28425 -9848
rect 22126 -9928 28425 -9912
rect 22126 -9992 28341 -9928
rect 28405 -9992 28425 -9928
rect 22126 -10008 28425 -9992
rect 22126 -10072 28341 -10008
rect 28405 -10072 28425 -10008
rect 22126 -10088 28425 -10072
rect 22126 -10152 28341 -10088
rect 28405 -10152 28425 -10088
rect 22126 -10168 28425 -10152
rect 22126 -10232 28341 -10168
rect 28405 -10232 28425 -10168
rect 22126 -10248 28425 -10232
rect 22126 -10312 28341 -10248
rect 28405 -10312 28425 -10248
rect 22126 -10328 28425 -10312
rect 22126 -10392 28341 -10328
rect 28405 -10392 28425 -10328
rect 22126 -10408 28425 -10392
rect 22126 -10472 28341 -10408
rect 28405 -10472 28425 -10408
rect 22126 -10488 28425 -10472
rect 22126 -10552 28341 -10488
rect 28405 -10552 28425 -10488
rect 22126 -10568 28425 -10552
rect 22126 -10632 28341 -10568
rect 28405 -10632 28425 -10568
rect 22126 -10648 28425 -10632
rect 22126 -10712 28341 -10648
rect 28405 -10712 28425 -10648
rect 22126 -10728 28425 -10712
rect 22126 -10792 28341 -10728
rect 28405 -10792 28425 -10728
rect 22126 -10808 28425 -10792
rect 22126 -10872 28341 -10808
rect 28405 -10872 28425 -10808
rect 22126 -10888 28425 -10872
rect 22126 -10952 28341 -10888
rect 28405 -10952 28425 -10888
rect 22126 -10968 28425 -10952
rect 22126 -11032 28341 -10968
rect 28405 -11032 28425 -10968
rect 22126 -11048 28425 -11032
rect 22126 -11112 28341 -11048
rect 28405 -11112 28425 -11048
rect 22126 -11128 28425 -11112
rect 22126 -11192 28341 -11128
rect 28405 -11192 28425 -11128
rect 22126 -11208 28425 -11192
rect 22126 -11272 28341 -11208
rect 28405 -11272 28425 -11208
rect 22126 -11288 28425 -11272
rect 22126 -11352 28341 -11288
rect 28405 -11352 28425 -11288
rect 22126 -11368 28425 -11352
rect 22126 -11432 28341 -11368
rect 28405 -11432 28425 -11368
rect 22126 -11448 28425 -11432
rect 22126 -11512 28341 -11448
rect 28405 -11512 28425 -11448
rect 22126 -11528 28425 -11512
rect 22126 -11592 28341 -11528
rect 28405 -11592 28425 -11528
rect 22126 -11608 28425 -11592
rect 22126 -11672 28341 -11608
rect 28405 -11672 28425 -11608
rect 22126 -11688 28425 -11672
rect 22126 -11752 28341 -11688
rect 28405 -11752 28425 -11688
rect 22126 -11768 28425 -11752
rect 22126 -11832 28341 -11768
rect 28405 -11832 28425 -11768
rect 22126 -11848 28425 -11832
rect 22126 -11912 28341 -11848
rect 28405 -11912 28425 -11848
rect 22126 -11928 28425 -11912
rect 22126 -11992 28341 -11928
rect 28405 -11992 28425 -11928
rect 22126 -12008 28425 -11992
rect 22126 -12072 28341 -12008
rect 28405 -12072 28425 -12008
rect 22126 -12088 28425 -12072
rect 22126 -12152 28341 -12088
rect 28405 -12152 28425 -12088
rect 22126 -12168 28425 -12152
rect 22126 -12232 28341 -12168
rect 28405 -12232 28425 -12168
rect 22126 -12248 28425 -12232
rect 22126 -12312 28341 -12248
rect 28405 -12312 28425 -12248
rect 22126 -12328 28425 -12312
rect 22126 -12392 28341 -12328
rect 28405 -12392 28425 -12328
rect 22126 -12408 28425 -12392
rect 22126 -12472 28341 -12408
rect 28405 -12472 28425 -12408
rect 22126 -12488 28425 -12472
rect 22126 -12552 28341 -12488
rect 28405 -12552 28425 -12488
rect 22126 -12568 28425 -12552
rect 22126 -12632 28341 -12568
rect 28405 -12632 28425 -12568
rect 22126 -12648 28425 -12632
rect 22126 -12712 28341 -12648
rect 28405 -12712 28425 -12648
rect 22126 -12728 28425 -12712
rect 22126 -12792 28341 -12728
rect 28405 -12792 28425 -12728
rect 22126 -12808 28425 -12792
rect 22126 -12872 28341 -12808
rect 28405 -12872 28425 -12808
rect 22126 -12888 28425 -12872
rect 22126 -12952 28341 -12888
rect 28405 -12952 28425 -12888
rect 22126 -12968 28425 -12952
rect 22126 -13032 28341 -12968
rect 28405 -13032 28425 -12968
rect 22126 -13048 28425 -13032
rect 22126 -13112 28341 -13048
rect 28405 -13112 28425 -13048
rect 22126 -13128 28425 -13112
rect 22126 -13192 28341 -13128
rect 28405 -13192 28425 -13128
rect 22126 -13208 28425 -13192
rect 22126 -13272 28341 -13208
rect 28405 -13272 28425 -13208
rect 22126 -13288 28425 -13272
rect 22126 -13352 28341 -13288
rect 28405 -13352 28425 -13288
rect 22126 -13368 28425 -13352
rect 22126 -13432 28341 -13368
rect 28405 -13432 28425 -13368
rect 22126 -13448 28425 -13432
rect 22126 -13512 28341 -13448
rect 28405 -13512 28425 -13448
rect 22126 -13528 28425 -13512
rect 22126 -13592 28341 -13528
rect 28405 -13592 28425 -13528
rect 22126 -13608 28425 -13592
rect 22126 -13672 28341 -13608
rect 28405 -13672 28425 -13608
rect 22126 -13688 28425 -13672
rect 22126 -13752 28341 -13688
rect 28405 -13752 28425 -13688
rect 22126 -13768 28425 -13752
rect 22126 -13832 28341 -13768
rect 28405 -13832 28425 -13768
rect 22126 -13848 28425 -13832
rect 22126 -13912 28341 -13848
rect 28405 -13912 28425 -13848
rect 22126 -13928 28425 -13912
rect 22126 -13992 28341 -13928
rect 28405 -13992 28425 -13928
rect 22126 -14008 28425 -13992
rect 22126 -14072 28341 -14008
rect 28405 -14072 28425 -14008
rect 22126 -14088 28425 -14072
rect 22126 -14152 28341 -14088
rect 28405 -14152 28425 -14088
rect 22126 -14168 28425 -14152
rect 22126 -14232 28341 -14168
rect 28405 -14232 28425 -14168
rect 22126 -14248 28425 -14232
rect 22126 -14312 28341 -14248
rect 28405 -14312 28425 -14248
rect 22126 -14328 28425 -14312
rect 22126 -14392 28341 -14328
rect 28405 -14392 28425 -14328
rect 22126 -14408 28425 -14392
rect 22126 -14472 28341 -14408
rect 28405 -14472 28425 -14408
rect 22126 -14488 28425 -14472
rect 22126 -14552 28341 -14488
rect 28405 -14552 28425 -14488
rect 22126 -14568 28425 -14552
rect 22126 -14632 28341 -14568
rect 28405 -14632 28425 -14568
rect 22126 -14648 28425 -14632
rect 22126 -14712 28341 -14648
rect 28405 -14712 28425 -14648
rect 22126 -14728 28425 -14712
rect 22126 -14792 28341 -14728
rect 28405 -14792 28425 -14728
rect 22126 -14808 28425 -14792
rect 22126 -14872 28341 -14808
rect 28405 -14872 28425 -14808
rect 22126 -14888 28425 -14872
rect 22126 -14952 28341 -14888
rect 28405 -14952 28425 -14888
rect 22126 -14968 28425 -14952
rect 22126 -15032 28341 -14968
rect 28405 -15032 28425 -14968
rect 22126 -15048 28425 -15032
rect 22126 -15112 28341 -15048
rect 28405 -15112 28425 -15048
rect 22126 -15128 28425 -15112
rect 22126 -15192 28341 -15128
rect 28405 -15192 28425 -15128
rect 22126 -15208 28425 -15192
rect 22126 -15272 28341 -15208
rect 28405 -15272 28425 -15208
rect 22126 -15288 28425 -15272
rect 22126 -15352 28341 -15288
rect 28405 -15352 28425 -15288
rect 22126 -15368 28425 -15352
rect 22126 -15432 28341 -15368
rect 28405 -15432 28425 -15368
rect 22126 -15448 28425 -15432
rect 22126 -15512 28341 -15448
rect 28405 -15512 28425 -15448
rect 22126 -15528 28425 -15512
rect 22126 -15592 28341 -15528
rect 28405 -15592 28425 -15528
rect 22126 -15608 28425 -15592
rect 22126 -15672 28341 -15608
rect 28405 -15672 28425 -15608
rect 22126 -15700 28425 -15672
rect 28445 -9528 34744 -9500
rect 28445 -9592 34660 -9528
rect 34724 -9592 34744 -9528
rect 28445 -9608 34744 -9592
rect 28445 -9672 34660 -9608
rect 34724 -9672 34744 -9608
rect 28445 -9688 34744 -9672
rect 28445 -9752 34660 -9688
rect 34724 -9752 34744 -9688
rect 28445 -9768 34744 -9752
rect 28445 -9832 34660 -9768
rect 34724 -9832 34744 -9768
rect 28445 -9848 34744 -9832
rect 28445 -9912 34660 -9848
rect 34724 -9912 34744 -9848
rect 28445 -9928 34744 -9912
rect 28445 -9992 34660 -9928
rect 34724 -9992 34744 -9928
rect 28445 -10008 34744 -9992
rect 28445 -10072 34660 -10008
rect 34724 -10072 34744 -10008
rect 28445 -10088 34744 -10072
rect 28445 -10152 34660 -10088
rect 34724 -10152 34744 -10088
rect 28445 -10168 34744 -10152
rect 28445 -10232 34660 -10168
rect 34724 -10232 34744 -10168
rect 28445 -10248 34744 -10232
rect 28445 -10312 34660 -10248
rect 34724 -10312 34744 -10248
rect 28445 -10328 34744 -10312
rect 28445 -10392 34660 -10328
rect 34724 -10392 34744 -10328
rect 28445 -10408 34744 -10392
rect 28445 -10472 34660 -10408
rect 34724 -10472 34744 -10408
rect 28445 -10488 34744 -10472
rect 28445 -10552 34660 -10488
rect 34724 -10552 34744 -10488
rect 28445 -10568 34744 -10552
rect 28445 -10632 34660 -10568
rect 34724 -10632 34744 -10568
rect 28445 -10648 34744 -10632
rect 28445 -10712 34660 -10648
rect 34724 -10712 34744 -10648
rect 28445 -10728 34744 -10712
rect 28445 -10792 34660 -10728
rect 34724 -10792 34744 -10728
rect 28445 -10808 34744 -10792
rect 28445 -10872 34660 -10808
rect 34724 -10872 34744 -10808
rect 28445 -10888 34744 -10872
rect 28445 -10952 34660 -10888
rect 34724 -10952 34744 -10888
rect 28445 -10968 34744 -10952
rect 28445 -11032 34660 -10968
rect 34724 -11032 34744 -10968
rect 28445 -11048 34744 -11032
rect 28445 -11112 34660 -11048
rect 34724 -11112 34744 -11048
rect 28445 -11128 34744 -11112
rect 28445 -11192 34660 -11128
rect 34724 -11192 34744 -11128
rect 28445 -11208 34744 -11192
rect 28445 -11272 34660 -11208
rect 34724 -11272 34744 -11208
rect 28445 -11288 34744 -11272
rect 28445 -11352 34660 -11288
rect 34724 -11352 34744 -11288
rect 28445 -11368 34744 -11352
rect 28445 -11432 34660 -11368
rect 34724 -11432 34744 -11368
rect 28445 -11448 34744 -11432
rect 28445 -11512 34660 -11448
rect 34724 -11512 34744 -11448
rect 28445 -11528 34744 -11512
rect 28445 -11592 34660 -11528
rect 34724 -11592 34744 -11528
rect 28445 -11608 34744 -11592
rect 28445 -11672 34660 -11608
rect 34724 -11672 34744 -11608
rect 28445 -11688 34744 -11672
rect 28445 -11752 34660 -11688
rect 34724 -11752 34744 -11688
rect 28445 -11768 34744 -11752
rect 28445 -11832 34660 -11768
rect 34724 -11832 34744 -11768
rect 28445 -11848 34744 -11832
rect 28445 -11912 34660 -11848
rect 34724 -11912 34744 -11848
rect 28445 -11928 34744 -11912
rect 28445 -11992 34660 -11928
rect 34724 -11992 34744 -11928
rect 28445 -12008 34744 -11992
rect 28445 -12072 34660 -12008
rect 34724 -12072 34744 -12008
rect 28445 -12088 34744 -12072
rect 28445 -12152 34660 -12088
rect 34724 -12152 34744 -12088
rect 28445 -12168 34744 -12152
rect 28445 -12232 34660 -12168
rect 34724 -12232 34744 -12168
rect 28445 -12248 34744 -12232
rect 28445 -12312 34660 -12248
rect 34724 -12312 34744 -12248
rect 28445 -12328 34744 -12312
rect 28445 -12392 34660 -12328
rect 34724 -12392 34744 -12328
rect 28445 -12408 34744 -12392
rect 28445 -12472 34660 -12408
rect 34724 -12472 34744 -12408
rect 28445 -12488 34744 -12472
rect 28445 -12552 34660 -12488
rect 34724 -12552 34744 -12488
rect 28445 -12568 34744 -12552
rect 28445 -12632 34660 -12568
rect 34724 -12632 34744 -12568
rect 28445 -12648 34744 -12632
rect 28445 -12712 34660 -12648
rect 34724 -12712 34744 -12648
rect 28445 -12728 34744 -12712
rect 28445 -12792 34660 -12728
rect 34724 -12792 34744 -12728
rect 28445 -12808 34744 -12792
rect 28445 -12872 34660 -12808
rect 34724 -12872 34744 -12808
rect 28445 -12888 34744 -12872
rect 28445 -12952 34660 -12888
rect 34724 -12952 34744 -12888
rect 28445 -12968 34744 -12952
rect 28445 -13032 34660 -12968
rect 34724 -13032 34744 -12968
rect 28445 -13048 34744 -13032
rect 28445 -13112 34660 -13048
rect 34724 -13112 34744 -13048
rect 28445 -13128 34744 -13112
rect 28445 -13192 34660 -13128
rect 34724 -13192 34744 -13128
rect 28445 -13208 34744 -13192
rect 28445 -13272 34660 -13208
rect 34724 -13272 34744 -13208
rect 28445 -13288 34744 -13272
rect 28445 -13352 34660 -13288
rect 34724 -13352 34744 -13288
rect 28445 -13368 34744 -13352
rect 28445 -13432 34660 -13368
rect 34724 -13432 34744 -13368
rect 28445 -13448 34744 -13432
rect 28445 -13512 34660 -13448
rect 34724 -13512 34744 -13448
rect 28445 -13528 34744 -13512
rect 28445 -13592 34660 -13528
rect 34724 -13592 34744 -13528
rect 28445 -13608 34744 -13592
rect 28445 -13672 34660 -13608
rect 34724 -13672 34744 -13608
rect 28445 -13688 34744 -13672
rect 28445 -13752 34660 -13688
rect 34724 -13752 34744 -13688
rect 28445 -13768 34744 -13752
rect 28445 -13832 34660 -13768
rect 34724 -13832 34744 -13768
rect 28445 -13848 34744 -13832
rect 28445 -13912 34660 -13848
rect 34724 -13912 34744 -13848
rect 28445 -13928 34744 -13912
rect 28445 -13992 34660 -13928
rect 34724 -13992 34744 -13928
rect 28445 -14008 34744 -13992
rect 28445 -14072 34660 -14008
rect 34724 -14072 34744 -14008
rect 28445 -14088 34744 -14072
rect 28445 -14152 34660 -14088
rect 34724 -14152 34744 -14088
rect 28445 -14168 34744 -14152
rect 28445 -14232 34660 -14168
rect 34724 -14232 34744 -14168
rect 28445 -14248 34744 -14232
rect 28445 -14312 34660 -14248
rect 34724 -14312 34744 -14248
rect 28445 -14328 34744 -14312
rect 28445 -14392 34660 -14328
rect 34724 -14392 34744 -14328
rect 28445 -14408 34744 -14392
rect 28445 -14472 34660 -14408
rect 34724 -14472 34744 -14408
rect 28445 -14488 34744 -14472
rect 28445 -14552 34660 -14488
rect 34724 -14552 34744 -14488
rect 28445 -14568 34744 -14552
rect 28445 -14632 34660 -14568
rect 34724 -14632 34744 -14568
rect 28445 -14648 34744 -14632
rect 28445 -14712 34660 -14648
rect 34724 -14712 34744 -14648
rect 28445 -14728 34744 -14712
rect 28445 -14792 34660 -14728
rect 34724 -14792 34744 -14728
rect 28445 -14808 34744 -14792
rect 28445 -14872 34660 -14808
rect 34724 -14872 34744 -14808
rect 28445 -14888 34744 -14872
rect 28445 -14952 34660 -14888
rect 34724 -14952 34744 -14888
rect 28445 -14968 34744 -14952
rect 28445 -15032 34660 -14968
rect 34724 -15032 34744 -14968
rect 28445 -15048 34744 -15032
rect 28445 -15112 34660 -15048
rect 34724 -15112 34744 -15048
rect 28445 -15128 34744 -15112
rect 28445 -15192 34660 -15128
rect 34724 -15192 34744 -15128
rect 28445 -15208 34744 -15192
rect 28445 -15272 34660 -15208
rect 34724 -15272 34744 -15208
rect 28445 -15288 34744 -15272
rect 28445 -15352 34660 -15288
rect 34724 -15352 34744 -15288
rect 28445 -15368 34744 -15352
rect 28445 -15432 34660 -15368
rect 34724 -15432 34744 -15368
rect 28445 -15448 34744 -15432
rect 28445 -15512 34660 -15448
rect 34724 -15512 34744 -15448
rect 28445 -15528 34744 -15512
rect 28445 -15592 34660 -15528
rect 34724 -15592 34744 -15528
rect 28445 -15608 34744 -15592
rect 28445 -15672 34660 -15608
rect 34724 -15672 34744 -15608
rect 28445 -15700 34744 -15672
rect 34764 -9528 41063 -9500
rect 34764 -9592 40979 -9528
rect 41043 -9592 41063 -9528
rect 34764 -9608 41063 -9592
rect 34764 -9672 40979 -9608
rect 41043 -9672 41063 -9608
rect 34764 -9688 41063 -9672
rect 34764 -9752 40979 -9688
rect 41043 -9752 41063 -9688
rect 34764 -9768 41063 -9752
rect 34764 -9832 40979 -9768
rect 41043 -9832 41063 -9768
rect 34764 -9848 41063 -9832
rect 34764 -9912 40979 -9848
rect 41043 -9912 41063 -9848
rect 34764 -9928 41063 -9912
rect 34764 -9992 40979 -9928
rect 41043 -9992 41063 -9928
rect 34764 -10008 41063 -9992
rect 34764 -10072 40979 -10008
rect 41043 -10072 41063 -10008
rect 34764 -10088 41063 -10072
rect 34764 -10152 40979 -10088
rect 41043 -10152 41063 -10088
rect 34764 -10168 41063 -10152
rect 34764 -10232 40979 -10168
rect 41043 -10232 41063 -10168
rect 34764 -10248 41063 -10232
rect 34764 -10312 40979 -10248
rect 41043 -10312 41063 -10248
rect 34764 -10328 41063 -10312
rect 34764 -10392 40979 -10328
rect 41043 -10392 41063 -10328
rect 34764 -10408 41063 -10392
rect 34764 -10472 40979 -10408
rect 41043 -10472 41063 -10408
rect 34764 -10488 41063 -10472
rect 34764 -10552 40979 -10488
rect 41043 -10552 41063 -10488
rect 34764 -10568 41063 -10552
rect 34764 -10632 40979 -10568
rect 41043 -10632 41063 -10568
rect 34764 -10648 41063 -10632
rect 34764 -10712 40979 -10648
rect 41043 -10712 41063 -10648
rect 34764 -10728 41063 -10712
rect 34764 -10792 40979 -10728
rect 41043 -10792 41063 -10728
rect 34764 -10808 41063 -10792
rect 34764 -10872 40979 -10808
rect 41043 -10872 41063 -10808
rect 34764 -10888 41063 -10872
rect 34764 -10952 40979 -10888
rect 41043 -10952 41063 -10888
rect 34764 -10968 41063 -10952
rect 34764 -11032 40979 -10968
rect 41043 -11032 41063 -10968
rect 34764 -11048 41063 -11032
rect 34764 -11112 40979 -11048
rect 41043 -11112 41063 -11048
rect 34764 -11128 41063 -11112
rect 34764 -11192 40979 -11128
rect 41043 -11192 41063 -11128
rect 34764 -11208 41063 -11192
rect 34764 -11272 40979 -11208
rect 41043 -11272 41063 -11208
rect 34764 -11288 41063 -11272
rect 34764 -11352 40979 -11288
rect 41043 -11352 41063 -11288
rect 34764 -11368 41063 -11352
rect 34764 -11432 40979 -11368
rect 41043 -11432 41063 -11368
rect 34764 -11448 41063 -11432
rect 34764 -11512 40979 -11448
rect 41043 -11512 41063 -11448
rect 34764 -11528 41063 -11512
rect 34764 -11592 40979 -11528
rect 41043 -11592 41063 -11528
rect 34764 -11608 41063 -11592
rect 34764 -11672 40979 -11608
rect 41043 -11672 41063 -11608
rect 34764 -11688 41063 -11672
rect 34764 -11752 40979 -11688
rect 41043 -11752 41063 -11688
rect 34764 -11768 41063 -11752
rect 34764 -11832 40979 -11768
rect 41043 -11832 41063 -11768
rect 34764 -11848 41063 -11832
rect 34764 -11912 40979 -11848
rect 41043 -11912 41063 -11848
rect 34764 -11928 41063 -11912
rect 34764 -11992 40979 -11928
rect 41043 -11992 41063 -11928
rect 34764 -12008 41063 -11992
rect 34764 -12072 40979 -12008
rect 41043 -12072 41063 -12008
rect 34764 -12088 41063 -12072
rect 34764 -12152 40979 -12088
rect 41043 -12152 41063 -12088
rect 34764 -12168 41063 -12152
rect 34764 -12232 40979 -12168
rect 41043 -12232 41063 -12168
rect 34764 -12248 41063 -12232
rect 34764 -12312 40979 -12248
rect 41043 -12312 41063 -12248
rect 34764 -12328 41063 -12312
rect 34764 -12392 40979 -12328
rect 41043 -12392 41063 -12328
rect 34764 -12408 41063 -12392
rect 34764 -12472 40979 -12408
rect 41043 -12472 41063 -12408
rect 34764 -12488 41063 -12472
rect 34764 -12552 40979 -12488
rect 41043 -12552 41063 -12488
rect 34764 -12568 41063 -12552
rect 34764 -12632 40979 -12568
rect 41043 -12632 41063 -12568
rect 34764 -12648 41063 -12632
rect 34764 -12712 40979 -12648
rect 41043 -12712 41063 -12648
rect 34764 -12728 41063 -12712
rect 34764 -12792 40979 -12728
rect 41043 -12792 41063 -12728
rect 34764 -12808 41063 -12792
rect 34764 -12872 40979 -12808
rect 41043 -12872 41063 -12808
rect 34764 -12888 41063 -12872
rect 34764 -12952 40979 -12888
rect 41043 -12952 41063 -12888
rect 34764 -12968 41063 -12952
rect 34764 -13032 40979 -12968
rect 41043 -13032 41063 -12968
rect 34764 -13048 41063 -13032
rect 34764 -13112 40979 -13048
rect 41043 -13112 41063 -13048
rect 34764 -13128 41063 -13112
rect 34764 -13192 40979 -13128
rect 41043 -13192 41063 -13128
rect 34764 -13208 41063 -13192
rect 34764 -13272 40979 -13208
rect 41043 -13272 41063 -13208
rect 34764 -13288 41063 -13272
rect 34764 -13352 40979 -13288
rect 41043 -13352 41063 -13288
rect 34764 -13368 41063 -13352
rect 34764 -13432 40979 -13368
rect 41043 -13432 41063 -13368
rect 34764 -13448 41063 -13432
rect 34764 -13512 40979 -13448
rect 41043 -13512 41063 -13448
rect 34764 -13528 41063 -13512
rect 34764 -13592 40979 -13528
rect 41043 -13592 41063 -13528
rect 34764 -13608 41063 -13592
rect 34764 -13672 40979 -13608
rect 41043 -13672 41063 -13608
rect 34764 -13688 41063 -13672
rect 34764 -13752 40979 -13688
rect 41043 -13752 41063 -13688
rect 34764 -13768 41063 -13752
rect 34764 -13832 40979 -13768
rect 41043 -13832 41063 -13768
rect 34764 -13848 41063 -13832
rect 34764 -13912 40979 -13848
rect 41043 -13912 41063 -13848
rect 34764 -13928 41063 -13912
rect 34764 -13992 40979 -13928
rect 41043 -13992 41063 -13928
rect 34764 -14008 41063 -13992
rect 34764 -14072 40979 -14008
rect 41043 -14072 41063 -14008
rect 34764 -14088 41063 -14072
rect 34764 -14152 40979 -14088
rect 41043 -14152 41063 -14088
rect 34764 -14168 41063 -14152
rect 34764 -14232 40979 -14168
rect 41043 -14232 41063 -14168
rect 34764 -14248 41063 -14232
rect 34764 -14312 40979 -14248
rect 41043 -14312 41063 -14248
rect 34764 -14328 41063 -14312
rect 34764 -14392 40979 -14328
rect 41043 -14392 41063 -14328
rect 34764 -14408 41063 -14392
rect 34764 -14472 40979 -14408
rect 41043 -14472 41063 -14408
rect 34764 -14488 41063 -14472
rect 34764 -14552 40979 -14488
rect 41043 -14552 41063 -14488
rect 34764 -14568 41063 -14552
rect 34764 -14632 40979 -14568
rect 41043 -14632 41063 -14568
rect 34764 -14648 41063 -14632
rect 34764 -14712 40979 -14648
rect 41043 -14712 41063 -14648
rect 34764 -14728 41063 -14712
rect 34764 -14792 40979 -14728
rect 41043 -14792 41063 -14728
rect 34764 -14808 41063 -14792
rect 34764 -14872 40979 -14808
rect 41043 -14872 41063 -14808
rect 34764 -14888 41063 -14872
rect 34764 -14952 40979 -14888
rect 41043 -14952 41063 -14888
rect 34764 -14968 41063 -14952
rect 34764 -15032 40979 -14968
rect 41043 -15032 41063 -14968
rect 34764 -15048 41063 -15032
rect 34764 -15112 40979 -15048
rect 41043 -15112 41063 -15048
rect 34764 -15128 41063 -15112
rect 34764 -15192 40979 -15128
rect 41043 -15192 41063 -15128
rect 34764 -15208 41063 -15192
rect 34764 -15272 40979 -15208
rect 41043 -15272 41063 -15208
rect 34764 -15288 41063 -15272
rect 34764 -15352 40979 -15288
rect 41043 -15352 41063 -15288
rect 34764 -15368 41063 -15352
rect 34764 -15432 40979 -15368
rect 41043 -15432 41063 -15368
rect 34764 -15448 41063 -15432
rect 34764 -15512 40979 -15448
rect 41043 -15512 41063 -15448
rect 34764 -15528 41063 -15512
rect 34764 -15592 40979 -15528
rect 41043 -15592 41063 -15528
rect 34764 -15608 41063 -15592
rect 34764 -15672 40979 -15608
rect 41043 -15672 41063 -15608
rect 34764 -15700 41063 -15672
rect 41083 -9528 47382 -9500
rect 41083 -9592 47298 -9528
rect 47362 -9592 47382 -9528
rect 41083 -9608 47382 -9592
rect 41083 -9672 47298 -9608
rect 47362 -9672 47382 -9608
rect 41083 -9688 47382 -9672
rect 41083 -9752 47298 -9688
rect 47362 -9752 47382 -9688
rect 41083 -9768 47382 -9752
rect 41083 -9832 47298 -9768
rect 47362 -9832 47382 -9768
rect 41083 -9848 47382 -9832
rect 41083 -9912 47298 -9848
rect 47362 -9912 47382 -9848
rect 41083 -9928 47382 -9912
rect 41083 -9992 47298 -9928
rect 47362 -9992 47382 -9928
rect 41083 -10008 47382 -9992
rect 41083 -10072 47298 -10008
rect 47362 -10072 47382 -10008
rect 41083 -10088 47382 -10072
rect 41083 -10152 47298 -10088
rect 47362 -10152 47382 -10088
rect 41083 -10168 47382 -10152
rect 41083 -10232 47298 -10168
rect 47362 -10232 47382 -10168
rect 41083 -10248 47382 -10232
rect 41083 -10312 47298 -10248
rect 47362 -10312 47382 -10248
rect 41083 -10328 47382 -10312
rect 41083 -10392 47298 -10328
rect 47362 -10392 47382 -10328
rect 41083 -10408 47382 -10392
rect 41083 -10472 47298 -10408
rect 47362 -10472 47382 -10408
rect 41083 -10488 47382 -10472
rect 41083 -10552 47298 -10488
rect 47362 -10552 47382 -10488
rect 41083 -10568 47382 -10552
rect 41083 -10632 47298 -10568
rect 47362 -10632 47382 -10568
rect 41083 -10648 47382 -10632
rect 41083 -10712 47298 -10648
rect 47362 -10712 47382 -10648
rect 41083 -10728 47382 -10712
rect 41083 -10792 47298 -10728
rect 47362 -10792 47382 -10728
rect 41083 -10808 47382 -10792
rect 41083 -10872 47298 -10808
rect 47362 -10872 47382 -10808
rect 41083 -10888 47382 -10872
rect 41083 -10952 47298 -10888
rect 47362 -10952 47382 -10888
rect 41083 -10968 47382 -10952
rect 41083 -11032 47298 -10968
rect 47362 -11032 47382 -10968
rect 41083 -11048 47382 -11032
rect 41083 -11112 47298 -11048
rect 47362 -11112 47382 -11048
rect 41083 -11128 47382 -11112
rect 41083 -11192 47298 -11128
rect 47362 -11192 47382 -11128
rect 41083 -11208 47382 -11192
rect 41083 -11272 47298 -11208
rect 47362 -11272 47382 -11208
rect 41083 -11288 47382 -11272
rect 41083 -11352 47298 -11288
rect 47362 -11352 47382 -11288
rect 41083 -11368 47382 -11352
rect 41083 -11432 47298 -11368
rect 47362 -11432 47382 -11368
rect 41083 -11448 47382 -11432
rect 41083 -11512 47298 -11448
rect 47362 -11512 47382 -11448
rect 41083 -11528 47382 -11512
rect 41083 -11592 47298 -11528
rect 47362 -11592 47382 -11528
rect 41083 -11608 47382 -11592
rect 41083 -11672 47298 -11608
rect 47362 -11672 47382 -11608
rect 41083 -11688 47382 -11672
rect 41083 -11752 47298 -11688
rect 47362 -11752 47382 -11688
rect 41083 -11768 47382 -11752
rect 41083 -11832 47298 -11768
rect 47362 -11832 47382 -11768
rect 41083 -11848 47382 -11832
rect 41083 -11912 47298 -11848
rect 47362 -11912 47382 -11848
rect 41083 -11928 47382 -11912
rect 41083 -11992 47298 -11928
rect 47362 -11992 47382 -11928
rect 41083 -12008 47382 -11992
rect 41083 -12072 47298 -12008
rect 47362 -12072 47382 -12008
rect 41083 -12088 47382 -12072
rect 41083 -12152 47298 -12088
rect 47362 -12152 47382 -12088
rect 41083 -12168 47382 -12152
rect 41083 -12232 47298 -12168
rect 47362 -12232 47382 -12168
rect 41083 -12248 47382 -12232
rect 41083 -12312 47298 -12248
rect 47362 -12312 47382 -12248
rect 41083 -12328 47382 -12312
rect 41083 -12392 47298 -12328
rect 47362 -12392 47382 -12328
rect 41083 -12408 47382 -12392
rect 41083 -12472 47298 -12408
rect 47362 -12472 47382 -12408
rect 41083 -12488 47382 -12472
rect 41083 -12552 47298 -12488
rect 47362 -12552 47382 -12488
rect 41083 -12568 47382 -12552
rect 41083 -12632 47298 -12568
rect 47362 -12632 47382 -12568
rect 41083 -12648 47382 -12632
rect 41083 -12712 47298 -12648
rect 47362 -12712 47382 -12648
rect 41083 -12728 47382 -12712
rect 41083 -12792 47298 -12728
rect 47362 -12792 47382 -12728
rect 41083 -12808 47382 -12792
rect 41083 -12872 47298 -12808
rect 47362 -12872 47382 -12808
rect 41083 -12888 47382 -12872
rect 41083 -12952 47298 -12888
rect 47362 -12952 47382 -12888
rect 41083 -12968 47382 -12952
rect 41083 -13032 47298 -12968
rect 47362 -13032 47382 -12968
rect 41083 -13048 47382 -13032
rect 41083 -13112 47298 -13048
rect 47362 -13112 47382 -13048
rect 41083 -13128 47382 -13112
rect 41083 -13192 47298 -13128
rect 47362 -13192 47382 -13128
rect 41083 -13208 47382 -13192
rect 41083 -13272 47298 -13208
rect 47362 -13272 47382 -13208
rect 41083 -13288 47382 -13272
rect 41083 -13352 47298 -13288
rect 47362 -13352 47382 -13288
rect 41083 -13368 47382 -13352
rect 41083 -13432 47298 -13368
rect 47362 -13432 47382 -13368
rect 41083 -13448 47382 -13432
rect 41083 -13512 47298 -13448
rect 47362 -13512 47382 -13448
rect 41083 -13528 47382 -13512
rect 41083 -13592 47298 -13528
rect 47362 -13592 47382 -13528
rect 41083 -13608 47382 -13592
rect 41083 -13672 47298 -13608
rect 47362 -13672 47382 -13608
rect 41083 -13688 47382 -13672
rect 41083 -13752 47298 -13688
rect 47362 -13752 47382 -13688
rect 41083 -13768 47382 -13752
rect 41083 -13832 47298 -13768
rect 47362 -13832 47382 -13768
rect 41083 -13848 47382 -13832
rect 41083 -13912 47298 -13848
rect 47362 -13912 47382 -13848
rect 41083 -13928 47382 -13912
rect 41083 -13992 47298 -13928
rect 47362 -13992 47382 -13928
rect 41083 -14008 47382 -13992
rect 41083 -14072 47298 -14008
rect 47362 -14072 47382 -14008
rect 41083 -14088 47382 -14072
rect 41083 -14152 47298 -14088
rect 47362 -14152 47382 -14088
rect 41083 -14168 47382 -14152
rect 41083 -14232 47298 -14168
rect 47362 -14232 47382 -14168
rect 41083 -14248 47382 -14232
rect 41083 -14312 47298 -14248
rect 47362 -14312 47382 -14248
rect 41083 -14328 47382 -14312
rect 41083 -14392 47298 -14328
rect 47362 -14392 47382 -14328
rect 41083 -14408 47382 -14392
rect 41083 -14472 47298 -14408
rect 47362 -14472 47382 -14408
rect 41083 -14488 47382 -14472
rect 41083 -14552 47298 -14488
rect 47362 -14552 47382 -14488
rect 41083 -14568 47382 -14552
rect 41083 -14632 47298 -14568
rect 47362 -14632 47382 -14568
rect 41083 -14648 47382 -14632
rect 41083 -14712 47298 -14648
rect 47362 -14712 47382 -14648
rect 41083 -14728 47382 -14712
rect 41083 -14792 47298 -14728
rect 47362 -14792 47382 -14728
rect 41083 -14808 47382 -14792
rect 41083 -14872 47298 -14808
rect 47362 -14872 47382 -14808
rect 41083 -14888 47382 -14872
rect 41083 -14952 47298 -14888
rect 47362 -14952 47382 -14888
rect 41083 -14968 47382 -14952
rect 41083 -15032 47298 -14968
rect 47362 -15032 47382 -14968
rect 41083 -15048 47382 -15032
rect 41083 -15112 47298 -15048
rect 47362 -15112 47382 -15048
rect 41083 -15128 47382 -15112
rect 41083 -15192 47298 -15128
rect 47362 -15192 47382 -15128
rect 41083 -15208 47382 -15192
rect 41083 -15272 47298 -15208
rect 47362 -15272 47382 -15208
rect 41083 -15288 47382 -15272
rect 41083 -15352 47298 -15288
rect 47362 -15352 47382 -15288
rect 41083 -15368 47382 -15352
rect 41083 -15432 47298 -15368
rect 47362 -15432 47382 -15368
rect 41083 -15448 47382 -15432
rect 41083 -15512 47298 -15448
rect 47362 -15512 47382 -15448
rect 41083 -15528 47382 -15512
rect 41083 -15592 47298 -15528
rect 47362 -15592 47382 -15528
rect 41083 -15608 47382 -15592
rect 41083 -15672 47298 -15608
rect 47362 -15672 47382 -15608
rect 41083 -15700 47382 -15672
rect -47383 -15828 -41084 -15800
rect -47383 -15892 -41168 -15828
rect -41104 -15892 -41084 -15828
rect -47383 -15908 -41084 -15892
rect -47383 -15972 -41168 -15908
rect -41104 -15972 -41084 -15908
rect -47383 -15988 -41084 -15972
rect -47383 -16052 -41168 -15988
rect -41104 -16052 -41084 -15988
rect -47383 -16068 -41084 -16052
rect -47383 -16132 -41168 -16068
rect -41104 -16132 -41084 -16068
rect -47383 -16148 -41084 -16132
rect -47383 -16212 -41168 -16148
rect -41104 -16212 -41084 -16148
rect -47383 -16228 -41084 -16212
rect -47383 -16292 -41168 -16228
rect -41104 -16292 -41084 -16228
rect -47383 -16308 -41084 -16292
rect -47383 -16372 -41168 -16308
rect -41104 -16372 -41084 -16308
rect -47383 -16388 -41084 -16372
rect -47383 -16452 -41168 -16388
rect -41104 -16452 -41084 -16388
rect -47383 -16468 -41084 -16452
rect -47383 -16532 -41168 -16468
rect -41104 -16532 -41084 -16468
rect -47383 -16548 -41084 -16532
rect -47383 -16612 -41168 -16548
rect -41104 -16612 -41084 -16548
rect -47383 -16628 -41084 -16612
rect -47383 -16692 -41168 -16628
rect -41104 -16692 -41084 -16628
rect -47383 -16708 -41084 -16692
rect -47383 -16772 -41168 -16708
rect -41104 -16772 -41084 -16708
rect -47383 -16788 -41084 -16772
rect -47383 -16852 -41168 -16788
rect -41104 -16852 -41084 -16788
rect -47383 -16868 -41084 -16852
rect -47383 -16932 -41168 -16868
rect -41104 -16932 -41084 -16868
rect -47383 -16948 -41084 -16932
rect -47383 -17012 -41168 -16948
rect -41104 -17012 -41084 -16948
rect -47383 -17028 -41084 -17012
rect -47383 -17092 -41168 -17028
rect -41104 -17092 -41084 -17028
rect -47383 -17108 -41084 -17092
rect -47383 -17172 -41168 -17108
rect -41104 -17172 -41084 -17108
rect -47383 -17188 -41084 -17172
rect -47383 -17252 -41168 -17188
rect -41104 -17252 -41084 -17188
rect -47383 -17268 -41084 -17252
rect -47383 -17332 -41168 -17268
rect -41104 -17332 -41084 -17268
rect -47383 -17348 -41084 -17332
rect -47383 -17412 -41168 -17348
rect -41104 -17412 -41084 -17348
rect -47383 -17428 -41084 -17412
rect -47383 -17492 -41168 -17428
rect -41104 -17492 -41084 -17428
rect -47383 -17508 -41084 -17492
rect -47383 -17572 -41168 -17508
rect -41104 -17572 -41084 -17508
rect -47383 -17588 -41084 -17572
rect -47383 -17652 -41168 -17588
rect -41104 -17652 -41084 -17588
rect -47383 -17668 -41084 -17652
rect -47383 -17732 -41168 -17668
rect -41104 -17732 -41084 -17668
rect -47383 -17748 -41084 -17732
rect -47383 -17812 -41168 -17748
rect -41104 -17812 -41084 -17748
rect -47383 -17828 -41084 -17812
rect -47383 -17892 -41168 -17828
rect -41104 -17892 -41084 -17828
rect -47383 -17908 -41084 -17892
rect -47383 -17972 -41168 -17908
rect -41104 -17972 -41084 -17908
rect -47383 -17988 -41084 -17972
rect -47383 -18052 -41168 -17988
rect -41104 -18052 -41084 -17988
rect -47383 -18068 -41084 -18052
rect -47383 -18132 -41168 -18068
rect -41104 -18132 -41084 -18068
rect -47383 -18148 -41084 -18132
rect -47383 -18212 -41168 -18148
rect -41104 -18212 -41084 -18148
rect -47383 -18228 -41084 -18212
rect -47383 -18292 -41168 -18228
rect -41104 -18292 -41084 -18228
rect -47383 -18308 -41084 -18292
rect -47383 -18372 -41168 -18308
rect -41104 -18372 -41084 -18308
rect -47383 -18388 -41084 -18372
rect -47383 -18452 -41168 -18388
rect -41104 -18452 -41084 -18388
rect -47383 -18468 -41084 -18452
rect -47383 -18532 -41168 -18468
rect -41104 -18532 -41084 -18468
rect -47383 -18548 -41084 -18532
rect -47383 -18612 -41168 -18548
rect -41104 -18612 -41084 -18548
rect -47383 -18628 -41084 -18612
rect -47383 -18692 -41168 -18628
rect -41104 -18692 -41084 -18628
rect -47383 -18708 -41084 -18692
rect -47383 -18772 -41168 -18708
rect -41104 -18772 -41084 -18708
rect -47383 -18788 -41084 -18772
rect -47383 -18852 -41168 -18788
rect -41104 -18852 -41084 -18788
rect -47383 -18868 -41084 -18852
rect -47383 -18932 -41168 -18868
rect -41104 -18932 -41084 -18868
rect -47383 -18948 -41084 -18932
rect -47383 -19012 -41168 -18948
rect -41104 -19012 -41084 -18948
rect -47383 -19028 -41084 -19012
rect -47383 -19092 -41168 -19028
rect -41104 -19092 -41084 -19028
rect -47383 -19108 -41084 -19092
rect -47383 -19172 -41168 -19108
rect -41104 -19172 -41084 -19108
rect -47383 -19188 -41084 -19172
rect -47383 -19252 -41168 -19188
rect -41104 -19252 -41084 -19188
rect -47383 -19268 -41084 -19252
rect -47383 -19332 -41168 -19268
rect -41104 -19332 -41084 -19268
rect -47383 -19348 -41084 -19332
rect -47383 -19412 -41168 -19348
rect -41104 -19412 -41084 -19348
rect -47383 -19428 -41084 -19412
rect -47383 -19492 -41168 -19428
rect -41104 -19492 -41084 -19428
rect -47383 -19508 -41084 -19492
rect -47383 -19572 -41168 -19508
rect -41104 -19572 -41084 -19508
rect -47383 -19588 -41084 -19572
rect -47383 -19652 -41168 -19588
rect -41104 -19652 -41084 -19588
rect -47383 -19668 -41084 -19652
rect -47383 -19732 -41168 -19668
rect -41104 -19732 -41084 -19668
rect -47383 -19748 -41084 -19732
rect -47383 -19812 -41168 -19748
rect -41104 -19812 -41084 -19748
rect -47383 -19828 -41084 -19812
rect -47383 -19892 -41168 -19828
rect -41104 -19892 -41084 -19828
rect -47383 -19908 -41084 -19892
rect -47383 -19972 -41168 -19908
rect -41104 -19972 -41084 -19908
rect -47383 -19988 -41084 -19972
rect -47383 -20052 -41168 -19988
rect -41104 -20052 -41084 -19988
rect -47383 -20068 -41084 -20052
rect -47383 -20132 -41168 -20068
rect -41104 -20132 -41084 -20068
rect -47383 -20148 -41084 -20132
rect -47383 -20212 -41168 -20148
rect -41104 -20212 -41084 -20148
rect -47383 -20228 -41084 -20212
rect -47383 -20292 -41168 -20228
rect -41104 -20292 -41084 -20228
rect -47383 -20308 -41084 -20292
rect -47383 -20372 -41168 -20308
rect -41104 -20372 -41084 -20308
rect -47383 -20388 -41084 -20372
rect -47383 -20452 -41168 -20388
rect -41104 -20452 -41084 -20388
rect -47383 -20468 -41084 -20452
rect -47383 -20532 -41168 -20468
rect -41104 -20532 -41084 -20468
rect -47383 -20548 -41084 -20532
rect -47383 -20612 -41168 -20548
rect -41104 -20612 -41084 -20548
rect -47383 -20628 -41084 -20612
rect -47383 -20692 -41168 -20628
rect -41104 -20692 -41084 -20628
rect -47383 -20708 -41084 -20692
rect -47383 -20772 -41168 -20708
rect -41104 -20772 -41084 -20708
rect -47383 -20788 -41084 -20772
rect -47383 -20852 -41168 -20788
rect -41104 -20852 -41084 -20788
rect -47383 -20868 -41084 -20852
rect -47383 -20932 -41168 -20868
rect -41104 -20932 -41084 -20868
rect -47383 -20948 -41084 -20932
rect -47383 -21012 -41168 -20948
rect -41104 -21012 -41084 -20948
rect -47383 -21028 -41084 -21012
rect -47383 -21092 -41168 -21028
rect -41104 -21092 -41084 -21028
rect -47383 -21108 -41084 -21092
rect -47383 -21172 -41168 -21108
rect -41104 -21172 -41084 -21108
rect -47383 -21188 -41084 -21172
rect -47383 -21252 -41168 -21188
rect -41104 -21252 -41084 -21188
rect -47383 -21268 -41084 -21252
rect -47383 -21332 -41168 -21268
rect -41104 -21332 -41084 -21268
rect -47383 -21348 -41084 -21332
rect -47383 -21412 -41168 -21348
rect -41104 -21412 -41084 -21348
rect -47383 -21428 -41084 -21412
rect -47383 -21492 -41168 -21428
rect -41104 -21492 -41084 -21428
rect -47383 -21508 -41084 -21492
rect -47383 -21572 -41168 -21508
rect -41104 -21572 -41084 -21508
rect -47383 -21588 -41084 -21572
rect -47383 -21652 -41168 -21588
rect -41104 -21652 -41084 -21588
rect -47383 -21668 -41084 -21652
rect -47383 -21732 -41168 -21668
rect -41104 -21732 -41084 -21668
rect -47383 -21748 -41084 -21732
rect -47383 -21812 -41168 -21748
rect -41104 -21812 -41084 -21748
rect -47383 -21828 -41084 -21812
rect -47383 -21892 -41168 -21828
rect -41104 -21892 -41084 -21828
rect -47383 -21908 -41084 -21892
rect -47383 -21972 -41168 -21908
rect -41104 -21972 -41084 -21908
rect -47383 -22000 -41084 -21972
rect -41064 -15828 -34765 -15800
rect -41064 -15892 -34849 -15828
rect -34785 -15892 -34765 -15828
rect -41064 -15908 -34765 -15892
rect -41064 -15972 -34849 -15908
rect -34785 -15972 -34765 -15908
rect -41064 -15988 -34765 -15972
rect -41064 -16052 -34849 -15988
rect -34785 -16052 -34765 -15988
rect -41064 -16068 -34765 -16052
rect -41064 -16132 -34849 -16068
rect -34785 -16132 -34765 -16068
rect -41064 -16148 -34765 -16132
rect -41064 -16212 -34849 -16148
rect -34785 -16212 -34765 -16148
rect -41064 -16228 -34765 -16212
rect -41064 -16292 -34849 -16228
rect -34785 -16292 -34765 -16228
rect -41064 -16308 -34765 -16292
rect -41064 -16372 -34849 -16308
rect -34785 -16372 -34765 -16308
rect -41064 -16388 -34765 -16372
rect -41064 -16452 -34849 -16388
rect -34785 -16452 -34765 -16388
rect -41064 -16468 -34765 -16452
rect -41064 -16532 -34849 -16468
rect -34785 -16532 -34765 -16468
rect -41064 -16548 -34765 -16532
rect -41064 -16612 -34849 -16548
rect -34785 -16612 -34765 -16548
rect -41064 -16628 -34765 -16612
rect -41064 -16692 -34849 -16628
rect -34785 -16692 -34765 -16628
rect -41064 -16708 -34765 -16692
rect -41064 -16772 -34849 -16708
rect -34785 -16772 -34765 -16708
rect -41064 -16788 -34765 -16772
rect -41064 -16852 -34849 -16788
rect -34785 -16852 -34765 -16788
rect -41064 -16868 -34765 -16852
rect -41064 -16932 -34849 -16868
rect -34785 -16932 -34765 -16868
rect -41064 -16948 -34765 -16932
rect -41064 -17012 -34849 -16948
rect -34785 -17012 -34765 -16948
rect -41064 -17028 -34765 -17012
rect -41064 -17092 -34849 -17028
rect -34785 -17092 -34765 -17028
rect -41064 -17108 -34765 -17092
rect -41064 -17172 -34849 -17108
rect -34785 -17172 -34765 -17108
rect -41064 -17188 -34765 -17172
rect -41064 -17252 -34849 -17188
rect -34785 -17252 -34765 -17188
rect -41064 -17268 -34765 -17252
rect -41064 -17332 -34849 -17268
rect -34785 -17332 -34765 -17268
rect -41064 -17348 -34765 -17332
rect -41064 -17412 -34849 -17348
rect -34785 -17412 -34765 -17348
rect -41064 -17428 -34765 -17412
rect -41064 -17492 -34849 -17428
rect -34785 -17492 -34765 -17428
rect -41064 -17508 -34765 -17492
rect -41064 -17572 -34849 -17508
rect -34785 -17572 -34765 -17508
rect -41064 -17588 -34765 -17572
rect -41064 -17652 -34849 -17588
rect -34785 -17652 -34765 -17588
rect -41064 -17668 -34765 -17652
rect -41064 -17732 -34849 -17668
rect -34785 -17732 -34765 -17668
rect -41064 -17748 -34765 -17732
rect -41064 -17812 -34849 -17748
rect -34785 -17812 -34765 -17748
rect -41064 -17828 -34765 -17812
rect -41064 -17892 -34849 -17828
rect -34785 -17892 -34765 -17828
rect -41064 -17908 -34765 -17892
rect -41064 -17972 -34849 -17908
rect -34785 -17972 -34765 -17908
rect -41064 -17988 -34765 -17972
rect -41064 -18052 -34849 -17988
rect -34785 -18052 -34765 -17988
rect -41064 -18068 -34765 -18052
rect -41064 -18132 -34849 -18068
rect -34785 -18132 -34765 -18068
rect -41064 -18148 -34765 -18132
rect -41064 -18212 -34849 -18148
rect -34785 -18212 -34765 -18148
rect -41064 -18228 -34765 -18212
rect -41064 -18292 -34849 -18228
rect -34785 -18292 -34765 -18228
rect -41064 -18308 -34765 -18292
rect -41064 -18372 -34849 -18308
rect -34785 -18372 -34765 -18308
rect -41064 -18388 -34765 -18372
rect -41064 -18452 -34849 -18388
rect -34785 -18452 -34765 -18388
rect -41064 -18468 -34765 -18452
rect -41064 -18532 -34849 -18468
rect -34785 -18532 -34765 -18468
rect -41064 -18548 -34765 -18532
rect -41064 -18612 -34849 -18548
rect -34785 -18612 -34765 -18548
rect -41064 -18628 -34765 -18612
rect -41064 -18692 -34849 -18628
rect -34785 -18692 -34765 -18628
rect -41064 -18708 -34765 -18692
rect -41064 -18772 -34849 -18708
rect -34785 -18772 -34765 -18708
rect -41064 -18788 -34765 -18772
rect -41064 -18852 -34849 -18788
rect -34785 -18852 -34765 -18788
rect -41064 -18868 -34765 -18852
rect -41064 -18932 -34849 -18868
rect -34785 -18932 -34765 -18868
rect -41064 -18948 -34765 -18932
rect -41064 -19012 -34849 -18948
rect -34785 -19012 -34765 -18948
rect -41064 -19028 -34765 -19012
rect -41064 -19092 -34849 -19028
rect -34785 -19092 -34765 -19028
rect -41064 -19108 -34765 -19092
rect -41064 -19172 -34849 -19108
rect -34785 -19172 -34765 -19108
rect -41064 -19188 -34765 -19172
rect -41064 -19252 -34849 -19188
rect -34785 -19252 -34765 -19188
rect -41064 -19268 -34765 -19252
rect -41064 -19332 -34849 -19268
rect -34785 -19332 -34765 -19268
rect -41064 -19348 -34765 -19332
rect -41064 -19412 -34849 -19348
rect -34785 -19412 -34765 -19348
rect -41064 -19428 -34765 -19412
rect -41064 -19492 -34849 -19428
rect -34785 -19492 -34765 -19428
rect -41064 -19508 -34765 -19492
rect -41064 -19572 -34849 -19508
rect -34785 -19572 -34765 -19508
rect -41064 -19588 -34765 -19572
rect -41064 -19652 -34849 -19588
rect -34785 -19652 -34765 -19588
rect -41064 -19668 -34765 -19652
rect -41064 -19732 -34849 -19668
rect -34785 -19732 -34765 -19668
rect -41064 -19748 -34765 -19732
rect -41064 -19812 -34849 -19748
rect -34785 -19812 -34765 -19748
rect -41064 -19828 -34765 -19812
rect -41064 -19892 -34849 -19828
rect -34785 -19892 -34765 -19828
rect -41064 -19908 -34765 -19892
rect -41064 -19972 -34849 -19908
rect -34785 -19972 -34765 -19908
rect -41064 -19988 -34765 -19972
rect -41064 -20052 -34849 -19988
rect -34785 -20052 -34765 -19988
rect -41064 -20068 -34765 -20052
rect -41064 -20132 -34849 -20068
rect -34785 -20132 -34765 -20068
rect -41064 -20148 -34765 -20132
rect -41064 -20212 -34849 -20148
rect -34785 -20212 -34765 -20148
rect -41064 -20228 -34765 -20212
rect -41064 -20292 -34849 -20228
rect -34785 -20292 -34765 -20228
rect -41064 -20308 -34765 -20292
rect -41064 -20372 -34849 -20308
rect -34785 -20372 -34765 -20308
rect -41064 -20388 -34765 -20372
rect -41064 -20452 -34849 -20388
rect -34785 -20452 -34765 -20388
rect -41064 -20468 -34765 -20452
rect -41064 -20532 -34849 -20468
rect -34785 -20532 -34765 -20468
rect -41064 -20548 -34765 -20532
rect -41064 -20612 -34849 -20548
rect -34785 -20612 -34765 -20548
rect -41064 -20628 -34765 -20612
rect -41064 -20692 -34849 -20628
rect -34785 -20692 -34765 -20628
rect -41064 -20708 -34765 -20692
rect -41064 -20772 -34849 -20708
rect -34785 -20772 -34765 -20708
rect -41064 -20788 -34765 -20772
rect -41064 -20852 -34849 -20788
rect -34785 -20852 -34765 -20788
rect -41064 -20868 -34765 -20852
rect -41064 -20932 -34849 -20868
rect -34785 -20932 -34765 -20868
rect -41064 -20948 -34765 -20932
rect -41064 -21012 -34849 -20948
rect -34785 -21012 -34765 -20948
rect -41064 -21028 -34765 -21012
rect -41064 -21092 -34849 -21028
rect -34785 -21092 -34765 -21028
rect -41064 -21108 -34765 -21092
rect -41064 -21172 -34849 -21108
rect -34785 -21172 -34765 -21108
rect -41064 -21188 -34765 -21172
rect -41064 -21252 -34849 -21188
rect -34785 -21252 -34765 -21188
rect -41064 -21268 -34765 -21252
rect -41064 -21332 -34849 -21268
rect -34785 -21332 -34765 -21268
rect -41064 -21348 -34765 -21332
rect -41064 -21412 -34849 -21348
rect -34785 -21412 -34765 -21348
rect -41064 -21428 -34765 -21412
rect -41064 -21492 -34849 -21428
rect -34785 -21492 -34765 -21428
rect -41064 -21508 -34765 -21492
rect -41064 -21572 -34849 -21508
rect -34785 -21572 -34765 -21508
rect -41064 -21588 -34765 -21572
rect -41064 -21652 -34849 -21588
rect -34785 -21652 -34765 -21588
rect -41064 -21668 -34765 -21652
rect -41064 -21732 -34849 -21668
rect -34785 -21732 -34765 -21668
rect -41064 -21748 -34765 -21732
rect -41064 -21812 -34849 -21748
rect -34785 -21812 -34765 -21748
rect -41064 -21828 -34765 -21812
rect -41064 -21892 -34849 -21828
rect -34785 -21892 -34765 -21828
rect -41064 -21908 -34765 -21892
rect -41064 -21972 -34849 -21908
rect -34785 -21972 -34765 -21908
rect -41064 -22000 -34765 -21972
rect -34745 -15828 -28446 -15800
rect -34745 -15892 -28530 -15828
rect -28466 -15892 -28446 -15828
rect -34745 -15908 -28446 -15892
rect -34745 -15972 -28530 -15908
rect -28466 -15972 -28446 -15908
rect -34745 -15988 -28446 -15972
rect -34745 -16052 -28530 -15988
rect -28466 -16052 -28446 -15988
rect -34745 -16068 -28446 -16052
rect -34745 -16132 -28530 -16068
rect -28466 -16132 -28446 -16068
rect -34745 -16148 -28446 -16132
rect -34745 -16212 -28530 -16148
rect -28466 -16212 -28446 -16148
rect -34745 -16228 -28446 -16212
rect -34745 -16292 -28530 -16228
rect -28466 -16292 -28446 -16228
rect -34745 -16308 -28446 -16292
rect -34745 -16372 -28530 -16308
rect -28466 -16372 -28446 -16308
rect -34745 -16388 -28446 -16372
rect -34745 -16452 -28530 -16388
rect -28466 -16452 -28446 -16388
rect -34745 -16468 -28446 -16452
rect -34745 -16532 -28530 -16468
rect -28466 -16532 -28446 -16468
rect -34745 -16548 -28446 -16532
rect -34745 -16612 -28530 -16548
rect -28466 -16612 -28446 -16548
rect -34745 -16628 -28446 -16612
rect -34745 -16692 -28530 -16628
rect -28466 -16692 -28446 -16628
rect -34745 -16708 -28446 -16692
rect -34745 -16772 -28530 -16708
rect -28466 -16772 -28446 -16708
rect -34745 -16788 -28446 -16772
rect -34745 -16852 -28530 -16788
rect -28466 -16852 -28446 -16788
rect -34745 -16868 -28446 -16852
rect -34745 -16932 -28530 -16868
rect -28466 -16932 -28446 -16868
rect -34745 -16948 -28446 -16932
rect -34745 -17012 -28530 -16948
rect -28466 -17012 -28446 -16948
rect -34745 -17028 -28446 -17012
rect -34745 -17092 -28530 -17028
rect -28466 -17092 -28446 -17028
rect -34745 -17108 -28446 -17092
rect -34745 -17172 -28530 -17108
rect -28466 -17172 -28446 -17108
rect -34745 -17188 -28446 -17172
rect -34745 -17252 -28530 -17188
rect -28466 -17252 -28446 -17188
rect -34745 -17268 -28446 -17252
rect -34745 -17332 -28530 -17268
rect -28466 -17332 -28446 -17268
rect -34745 -17348 -28446 -17332
rect -34745 -17412 -28530 -17348
rect -28466 -17412 -28446 -17348
rect -34745 -17428 -28446 -17412
rect -34745 -17492 -28530 -17428
rect -28466 -17492 -28446 -17428
rect -34745 -17508 -28446 -17492
rect -34745 -17572 -28530 -17508
rect -28466 -17572 -28446 -17508
rect -34745 -17588 -28446 -17572
rect -34745 -17652 -28530 -17588
rect -28466 -17652 -28446 -17588
rect -34745 -17668 -28446 -17652
rect -34745 -17732 -28530 -17668
rect -28466 -17732 -28446 -17668
rect -34745 -17748 -28446 -17732
rect -34745 -17812 -28530 -17748
rect -28466 -17812 -28446 -17748
rect -34745 -17828 -28446 -17812
rect -34745 -17892 -28530 -17828
rect -28466 -17892 -28446 -17828
rect -34745 -17908 -28446 -17892
rect -34745 -17972 -28530 -17908
rect -28466 -17972 -28446 -17908
rect -34745 -17988 -28446 -17972
rect -34745 -18052 -28530 -17988
rect -28466 -18052 -28446 -17988
rect -34745 -18068 -28446 -18052
rect -34745 -18132 -28530 -18068
rect -28466 -18132 -28446 -18068
rect -34745 -18148 -28446 -18132
rect -34745 -18212 -28530 -18148
rect -28466 -18212 -28446 -18148
rect -34745 -18228 -28446 -18212
rect -34745 -18292 -28530 -18228
rect -28466 -18292 -28446 -18228
rect -34745 -18308 -28446 -18292
rect -34745 -18372 -28530 -18308
rect -28466 -18372 -28446 -18308
rect -34745 -18388 -28446 -18372
rect -34745 -18452 -28530 -18388
rect -28466 -18452 -28446 -18388
rect -34745 -18468 -28446 -18452
rect -34745 -18532 -28530 -18468
rect -28466 -18532 -28446 -18468
rect -34745 -18548 -28446 -18532
rect -34745 -18612 -28530 -18548
rect -28466 -18612 -28446 -18548
rect -34745 -18628 -28446 -18612
rect -34745 -18692 -28530 -18628
rect -28466 -18692 -28446 -18628
rect -34745 -18708 -28446 -18692
rect -34745 -18772 -28530 -18708
rect -28466 -18772 -28446 -18708
rect -34745 -18788 -28446 -18772
rect -34745 -18852 -28530 -18788
rect -28466 -18852 -28446 -18788
rect -34745 -18868 -28446 -18852
rect -34745 -18932 -28530 -18868
rect -28466 -18932 -28446 -18868
rect -34745 -18948 -28446 -18932
rect -34745 -19012 -28530 -18948
rect -28466 -19012 -28446 -18948
rect -34745 -19028 -28446 -19012
rect -34745 -19092 -28530 -19028
rect -28466 -19092 -28446 -19028
rect -34745 -19108 -28446 -19092
rect -34745 -19172 -28530 -19108
rect -28466 -19172 -28446 -19108
rect -34745 -19188 -28446 -19172
rect -34745 -19252 -28530 -19188
rect -28466 -19252 -28446 -19188
rect -34745 -19268 -28446 -19252
rect -34745 -19332 -28530 -19268
rect -28466 -19332 -28446 -19268
rect -34745 -19348 -28446 -19332
rect -34745 -19412 -28530 -19348
rect -28466 -19412 -28446 -19348
rect -34745 -19428 -28446 -19412
rect -34745 -19492 -28530 -19428
rect -28466 -19492 -28446 -19428
rect -34745 -19508 -28446 -19492
rect -34745 -19572 -28530 -19508
rect -28466 -19572 -28446 -19508
rect -34745 -19588 -28446 -19572
rect -34745 -19652 -28530 -19588
rect -28466 -19652 -28446 -19588
rect -34745 -19668 -28446 -19652
rect -34745 -19732 -28530 -19668
rect -28466 -19732 -28446 -19668
rect -34745 -19748 -28446 -19732
rect -34745 -19812 -28530 -19748
rect -28466 -19812 -28446 -19748
rect -34745 -19828 -28446 -19812
rect -34745 -19892 -28530 -19828
rect -28466 -19892 -28446 -19828
rect -34745 -19908 -28446 -19892
rect -34745 -19972 -28530 -19908
rect -28466 -19972 -28446 -19908
rect -34745 -19988 -28446 -19972
rect -34745 -20052 -28530 -19988
rect -28466 -20052 -28446 -19988
rect -34745 -20068 -28446 -20052
rect -34745 -20132 -28530 -20068
rect -28466 -20132 -28446 -20068
rect -34745 -20148 -28446 -20132
rect -34745 -20212 -28530 -20148
rect -28466 -20212 -28446 -20148
rect -34745 -20228 -28446 -20212
rect -34745 -20292 -28530 -20228
rect -28466 -20292 -28446 -20228
rect -34745 -20308 -28446 -20292
rect -34745 -20372 -28530 -20308
rect -28466 -20372 -28446 -20308
rect -34745 -20388 -28446 -20372
rect -34745 -20452 -28530 -20388
rect -28466 -20452 -28446 -20388
rect -34745 -20468 -28446 -20452
rect -34745 -20532 -28530 -20468
rect -28466 -20532 -28446 -20468
rect -34745 -20548 -28446 -20532
rect -34745 -20612 -28530 -20548
rect -28466 -20612 -28446 -20548
rect -34745 -20628 -28446 -20612
rect -34745 -20692 -28530 -20628
rect -28466 -20692 -28446 -20628
rect -34745 -20708 -28446 -20692
rect -34745 -20772 -28530 -20708
rect -28466 -20772 -28446 -20708
rect -34745 -20788 -28446 -20772
rect -34745 -20852 -28530 -20788
rect -28466 -20852 -28446 -20788
rect -34745 -20868 -28446 -20852
rect -34745 -20932 -28530 -20868
rect -28466 -20932 -28446 -20868
rect -34745 -20948 -28446 -20932
rect -34745 -21012 -28530 -20948
rect -28466 -21012 -28446 -20948
rect -34745 -21028 -28446 -21012
rect -34745 -21092 -28530 -21028
rect -28466 -21092 -28446 -21028
rect -34745 -21108 -28446 -21092
rect -34745 -21172 -28530 -21108
rect -28466 -21172 -28446 -21108
rect -34745 -21188 -28446 -21172
rect -34745 -21252 -28530 -21188
rect -28466 -21252 -28446 -21188
rect -34745 -21268 -28446 -21252
rect -34745 -21332 -28530 -21268
rect -28466 -21332 -28446 -21268
rect -34745 -21348 -28446 -21332
rect -34745 -21412 -28530 -21348
rect -28466 -21412 -28446 -21348
rect -34745 -21428 -28446 -21412
rect -34745 -21492 -28530 -21428
rect -28466 -21492 -28446 -21428
rect -34745 -21508 -28446 -21492
rect -34745 -21572 -28530 -21508
rect -28466 -21572 -28446 -21508
rect -34745 -21588 -28446 -21572
rect -34745 -21652 -28530 -21588
rect -28466 -21652 -28446 -21588
rect -34745 -21668 -28446 -21652
rect -34745 -21732 -28530 -21668
rect -28466 -21732 -28446 -21668
rect -34745 -21748 -28446 -21732
rect -34745 -21812 -28530 -21748
rect -28466 -21812 -28446 -21748
rect -34745 -21828 -28446 -21812
rect -34745 -21892 -28530 -21828
rect -28466 -21892 -28446 -21828
rect -34745 -21908 -28446 -21892
rect -34745 -21972 -28530 -21908
rect -28466 -21972 -28446 -21908
rect -34745 -22000 -28446 -21972
rect -28426 -15828 -22127 -15800
rect -28426 -15892 -22211 -15828
rect -22147 -15892 -22127 -15828
rect -28426 -15908 -22127 -15892
rect -28426 -15972 -22211 -15908
rect -22147 -15972 -22127 -15908
rect -28426 -15988 -22127 -15972
rect -28426 -16052 -22211 -15988
rect -22147 -16052 -22127 -15988
rect -28426 -16068 -22127 -16052
rect -28426 -16132 -22211 -16068
rect -22147 -16132 -22127 -16068
rect -28426 -16148 -22127 -16132
rect -28426 -16212 -22211 -16148
rect -22147 -16212 -22127 -16148
rect -28426 -16228 -22127 -16212
rect -28426 -16292 -22211 -16228
rect -22147 -16292 -22127 -16228
rect -28426 -16308 -22127 -16292
rect -28426 -16372 -22211 -16308
rect -22147 -16372 -22127 -16308
rect -28426 -16388 -22127 -16372
rect -28426 -16452 -22211 -16388
rect -22147 -16452 -22127 -16388
rect -28426 -16468 -22127 -16452
rect -28426 -16532 -22211 -16468
rect -22147 -16532 -22127 -16468
rect -28426 -16548 -22127 -16532
rect -28426 -16612 -22211 -16548
rect -22147 -16612 -22127 -16548
rect -28426 -16628 -22127 -16612
rect -28426 -16692 -22211 -16628
rect -22147 -16692 -22127 -16628
rect -28426 -16708 -22127 -16692
rect -28426 -16772 -22211 -16708
rect -22147 -16772 -22127 -16708
rect -28426 -16788 -22127 -16772
rect -28426 -16852 -22211 -16788
rect -22147 -16852 -22127 -16788
rect -28426 -16868 -22127 -16852
rect -28426 -16932 -22211 -16868
rect -22147 -16932 -22127 -16868
rect -28426 -16948 -22127 -16932
rect -28426 -17012 -22211 -16948
rect -22147 -17012 -22127 -16948
rect -28426 -17028 -22127 -17012
rect -28426 -17092 -22211 -17028
rect -22147 -17092 -22127 -17028
rect -28426 -17108 -22127 -17092
rect -28426 -17172 -22211 -17108
rect -22147 -17172 -22127 -17108
rect -28426 -17188 -22127 -17172
rect -28426 -17252 -22211 -17188
rect -22147 -17252 -22127 -17188
rect -28426 -17268 -22127 -17252
rect -28426 -17332 -22211 -17268
rect -22147 -17332 -22127 -17268
rect -28426 -17348 -22127 -17332
rect -28426 -17412 -22211 -17348
rect -22147 -17412 -22127 -17348
rect -28426 -17428 -22127 -17412
rect -28426 -17492 -22211 -17428
rect -22147 -17492 -22127 -17428
rect -28426 -17508 -22127 -17492
rect -28426 -17572 -22211 -17508
rect -22147 -17572 -22127 -17508
rect -28426 -17588 -22127 -17572
rect -28426 -17652 -22211 -17588
rect -22147 -17652 -22127 -17588
rect -28426 -17668 -22127 -17652
rect -28426 -17732 -22211 -17668
rect -22147 -17732 -22127 -17668
rect -28426 -17748 -22127 -17732
rect -28426 -17812 -22211 -17748
rect -22147 -17812 -22127 -17748
rect -28426 -17828 -22127 -17812
rect -28426 -17892 -22211 -17828
rect -22147 -17892 -22127 -17828
rect -28426 -17908 -22127 -17892
rect -28426 -17972 -22211 -17908
rect -22147 -17972 -22127 -17908
rect -28426 -17988 -22127 -17972
rect -28426 -18052 -22211 -17988
rect -22147 -18052 -22127 -17988
rect -28426 -18068 -22127 -18052
rect -28426 -18132 -22211 -18068
rect -22147 -18132 -22127 -18068
rect -28426 -18148 -22127 -18132
rect -28426 -18212 -22211 -18148
rect -22147 -18212 -22127 -18148
rect -28426 -18228 -22127 -18212
rect -28426 -18292 -22211 -18228
rect -22147 -18292 -22127 -18228
rect -28426 -18308 -22127 -18292
rect -28426 -18372 -22211 -18308
rect -22147 -18372 -22127 -18308
rect -28426 -18388 -22127 -18372
rect -28426 -18452 -22211 -18388
rect -22147 -18452 -22127 -18388
rect -28426 -18468 -22127 -18452
rect -28426 -18532 -22211 -18468
rect -22147 -18532 -22127 -18468
rect -28426 -18548 -22127 -18532
rect -28426 -18612 -22211 -18548
rect -22147 -18612 -22127 -18548
rect -28426 -18628 -22127 -18612
rect -28426 -18692 -22211 -18628
rect -22147 -18692 -22127 -18628
rect -28426 -18708 -22127 -18692
rect -28426 -18772 -22211 -18708
rect -22147 -18772 -22127 -18708
rect -28426 -18788 -22127 -18772
rect -28426 -18852 -22211 -18788
rect -22147 -18852 -22127 -18788
rect -28426 -18868 -22127 -18852
rect -28426 -18932 -22211 -18868
rect -22147 -18932 -22127 -18868
rect -28426 -18948 -22127 -18932
rect -28426 -19012 -22211 -18948
rect -22147 -19012 -22127 -18948
rect -28426 -19028 -22127 -19012
rect -28426 -19092 -22211 -19028
rect -22147 -19092 -22127 -19028
rect -28426 -19108 -22127 -19092
rect -28426 -19172 -22211 -19108
rect -22147 -19172 -22127 -19108
rect -28426 -19188 -22127 -19172
rect -28426 -19252 -22211 -19188
rect -22147 -19252 -22127 -19188
rect -28426 -19268 -22127 -19252
rect -28426 -19332 -22211 -19268
rect -22147 -19332 -22127 -19268
rect -28426 -19348 -22127 -19332
rect -28426 -19412 -22211 -19348
rect -22147 -19412 -22127 -19348
rect -28426 -19428 -22127 -19412
rect -28426 -19492 -22211 -19428
rect -22147 -19492 -22127 -19428
rect -28426 -19508 -22127 -19492
rect -28426 -19572 -22211 -19508
rect -22147 -19572 -22127 -19508
rect -28426 -19588 -22127 -19572
rect -28426 -19652 -22211 -19588
rect -22147 -19652 -22127 -19588
rect -28426 -19668 -22127 -19652
rect -28426 -19732 -22211 -19668
rect -22147 -19732 -22127 -19668
rect -28426 -19748 -22127 -19732
rect -28426 -19812 -22211 -19748
rect -22147 -19812 -22127 -19748
rect -28426 -19828 -22127 -19812
rect -28426 -19892 -22211 -19828
rect -22147 -19892 -22127 -19828
rect -28426 -19908 -22127 -19892
rect -28426 -19972 -22211 -19908
rect -22147 -19972 -22127 -19908
rect -28426 -19988 -22127 -19972
rect -28426 -20052 -22211 -19988
rect -22147 -20052 -22127 -19988
rect -28426 -20068 -22127 -20052
rect -28426 -20132 -22211 -20068
rect -22147 -20132 -22127 -20068
rect -28426 -20148 -22127 -20132
rect -28426 -20212 -22211 -20148
rect -22147 -20212 -22127 -20148
rect -28426 -20228 -22127 -20212
rect -28426 -20292 -22211 -20228
rect -22147 -20292 -22127 -20228
rect -28426 -20308 -22127 -20292
rect -28426 -20372 -22211 -20308
rect -22147 -20372 -22127 -20308
rect -28426 -20388 -22127 -20372
rect -28426 -20452 -22211 -20388
rect -22147 -20452 -22127 -20388
rect -28426 -20468 -22127 -20452
rect -28426 -20532 -22211 -20468
rect -22147 -20532 -22127 -20468
rect -28426 -20548 -22127 -20532
rect -28426 -20612 -22211 -20548
rect -22147 -20612 -22127 -20548
rect -28426 -20628 -22127 -20612
rect -28426 -20692 -22211 -20628
rect -22147 -20692 -22127 -20628
rect -28426 -20708 -22127 -20692
rect -28426 -20772 -22211 -20708
rect -22147 -20772 -22127 -20708
rect -28426 -20788 -22127 -20772
rect -28426 -20852 -22211 -20788
rect -22147 -20852 -22127 -20788
rect -28426 -20868 -22127 -20852
rect -28426 -20932 -22211 -20868
rect -22147 -20932 -22127 -20868
rect -28426 -20948 -22127 -20932
rect -28426 -21012 -22211 -20948
rect -22147 -21012 -22127 -20948
rect -28426 -21028 -22127 -21012
rect -28426 -21092 -22211 -21028
rect -22147 -21092 -22127 -21028
rect -28426 -21108 -22127 -21092
rect -28426 -21172 -22211 -21108
rect -22147 -21172 -22127 -21108
rect -28426 -21188 -22127 -21172
rect -28426 -21252 -22211 -21188
rect -22147 -21252 -22127 -21188
rect -28426 -21268 -22127 -21252
rect -28426 -21332 -22211 -21268
rect -22147 -21332 -22127 -21268
rect -28426 -21348 -22127 -21332
rect -28426 -21412 -22211 -21348
rect -22147 -21412 -22127 -21348
rect -28426 -21428 -22127 -21412
rect -28426 -21492 -22211 -21428
rect -22147 -21492 -22127 -21428
rect -28426 -21508 -22127 -21492
rect -28426 -21572 -22211 -21508
rect -22147 -21572 -22127 -21508
rect -28426 -21588 -22127 -21572
rect -28426 -21652 -22211 -21588
rect -22147 -21652 -22127 -21588
rect -28426 -21668 -22127 -21652
rect -28426 -21732 -22211 -21668
rect -22147 -21732 -22127 -21668
rect -28426 -21748 -22127 -21732
rect -28426 -21812 -22211 -21748
rect -22147 -21812 -22127 -21748
rect -28426 -21828 -22127 -21812
rect -28426 -21892 -22211 -21828
rect -22147 -21892 -22127 -21828
rect -28426 -21908 -22127 -21892
rect -28426 -21972 -22211 -21908
rect -22147 -21972 -22127 -21908
rect -28426 -22000 -22127 -21972
rect -22107 -15828 -15808 -15800
rect -22107 -15892 -15892 -15828
rect -15828 -15892 -15808 -15828
rect -22107 -15908 -15808 -15892
rect -22107 -15972 -15892 -15908
rect -15828 -15972 -15808 -15908
rect -22107 -15988 -15808 -15972
rect -22107 -16052 -15892 -15988
rect -15828 -16052 -15808 -15988
rect -22107 -16068 -15808 -16052
rect -22107 -16132 -15892 -16068
rect -15828 -16132 -15808 -16068
rect -22107 -16148 -15808 -16132
rect -22107 -16212 -15892 -16148
rect -15828 -16212 -15808 -16148
rect -22107 -16228 -15808 -16212
rect -22107 -16292 -15892 -16228
rect -15828 -16292 -15808 -16228
rect -22107 -16308 -15808 -16292
rect -22107 -16372 -15892 -16308
rect -15828 -16372 -15808 -16308
rect -22107 -16388 -15808 -16372
rect -22107 -16452 -15892 -16388
rect -15828 -16452 -15808 -16388
rect -22107 -16468 -15808 -16452
rect -22107 -16532 -15892 -16468
rect -15828 -16532 -15808 -16468
rect -22107 -16548 -15808 -16532
rect -22107 -16612 -15892 -16548
rect -15828 -16612 -15808 -16548
rect -22107 -16628 -15808 -16612
rect -22107 -16692 -15892 -16628
rect -15828 -16692 -15808 -16628
rect -22107 -16708 -15808 -16692
rect -22107 -16772 -15892 -16708
rect -15828 -16772 -15808 -16708
rect -22107 -16788 -15808 -16772
rect -22107 -16852 -15892 -16788
rect -15828 -16852 -15808 -16788
rect -22107 -16868 -15808 -16852
rect -22107 -16932 -15892 -16868
rect -15828 -16932 -15808 -16868
rect -22107 -16948 -15808 -16932
rect -22107 -17012 -15892 -16948
rect -15828 -17012 -15808 -16948
rect -22107 -17028 -15808 -17012
rect -22107 -17092 -15892 -17028
rect -15828 -17092 -15808 -17028
rect -22107 -17108 -15808 -17092
rect -22107 -17172 -15892 -17108
rect -15828 -17172 -15808 -17108
rect -22107 -17188 -15808 -17172
rect -22107 -17252 -15892 -17188
rect -15828 -17252 -15808 -17188
rect -22107 -17268 -15808 -17252
rect -22107 -17332 -15892 -17268
rect -15828 -17332 -15808 -17268
rect -22107 -17348 -15808 -17332
rect -22107 -17412 -15892 -17348
rect -15828 -17412 -15808 -17348
rect -22107 -17428 -15808 -17412
rect -22107 -17492 -15892 -17428
rect -15828 -17492 -15808 -17428
rect -22107 -17508 -15808 -17492
rect -22107 -17572 -15892 -17508
rect -15828 -17572 -15808 -17508
rect -22107 -17588 -15808 -17572
rect -22107 -17652 -15892 -17588
rect -15828 -17652 -15808 -17588
rect -22107 -17668 -15808 -17652
rect -22107 -17732 -15892 -17668
rect -15828 -17732 -15808 -17668
rect -22107 -17748 -15808 -17732
rect -22107 -17812 -15892 -17748
rect -15828 -17812 -15808 -17748
rect -22107 -17828 -15808 -17812
rect -22107 -17892 -15892 -17828
rect -15828 -17892 -15808 -17828
rect -22107 -17908 -15808 -17892
rect -22107 -17972 -15892 -17908
rect -15828 -17972 -15808 -17908
rect -22107 -17988 -15808 -17972
rect -22107 -18052 -15892 -17988
rect -15828 -18052 -15808 -17988
rect -22107 -18068 -15808 -18052
rect -22107 -18132 -15892 -18068
rect -15828 -18132 -15808 -18068
rect -22107 -18148 -15808 -18132
rect -22107 -18212 -15892 -18148
rect -15828 -18212 -15808 -18148
rect -22107 -18228 -15808 -18212
rect -22107 -18292 -15892 -18228
rect -15828 -18292 -15808 -18228
rect -22107 -18308 -15808 -18292
rect -22107 -18372 -15892 -18308
rect -15828 -18372 -15808 -18308
rect -22107 -18388 -15808 -18372
rect -22107 -18452 -15892 -18388
rect -15828 -18452 -15808 -18388
rect -22107 -18468 -15808 -18452
rect -22107 -18532 -15892 -18468
rect -15828 -18532 -15808 -18468
rect -22107 -18548 -15808 -18532
rect -22107 -18612 -15892 -18548
rect -15828 -18612 -15808 -18548
rect -22107 -18628 -15808 -18612
rect -22107 -18692 -15892 -18628
rect -15828 -18692 -15808 -18628
rect -22107 -18708 -15808 -18692
rect -22107 -18772 -15892 -18708
rect -15828 -18772 -15808 -18708
rect -22107 -18788 -15808 -18772
rect -22107 -18852 -15892 -18788
rect -15828 -18852 -15808 -18788
rect -22107 -18868 -15808 -18852
rect -22107 -18932 -15892 -18868
rect -15828 -18932 -15808 -18868
rect -22107 -18948 -15808 -18932
rect -22107 -19012 -15892 -18948
rect -15828 -19012 -15808 -18948
rect -22107 -19028 -15808 -19012
rect -22107 -19092 -15892 -19028
rect -15828 -19092 -15808 -19028
rect -22107 -19108 -15808 -19092
rect -22107 -19172 -15892 -19108
rect -15828 -19172 -15808 -19108
rect -22107 -19188 -15808 -19172
rect -22107 -19252 -15892 -19188
rect -15828 -19252 -15808 -19188
rect -22107 -19268 -15808 -19252
rect -22107 -19332 -15892 -19268
rect -15828 -19332 -15808 -19268
rect -22107 -19348 -15808 -19332
rect -22107 -19412 -15892 -19348
rect -15828 -19412 -15808 -19348
rect -22107 -19428 -15808 -19412
rect -22107 -19492 -15892 -19428
rect -15828 -19492 -15808 -19428
rect -22107 -19508 -15808 -19492
rect -22107 -19572 -15892 -19508
rect -15828 -19572 -15808 -19508
rect -22107 -19588 -15808 -19572
rect -22107 -19652 -15892 -19588
rect -15828 -19652 -15808 -19588
rect -22107 -19668 -15808 -19652
rect -22107 -19732 -15892 -19668
rect -15828 -19732 -15808 -19668
rect -22107 -19748 -15808 -19732
rect -22107 -19812 -15892 -19748
rect -15828 -19812 -15808 -19748
rect -22107 -19828 -15808 -19812
rect -22107 -19892 -15892 -19828
rect -15828 -19892 -15808 -19828
rect -22107 -19908 -15808 -19892
rect -22107 -19972 -15892 -19908
rect -15828 -19972 -15808 -19908
rect -22107 -19988 -15808 -19972
rect -22107 -20052 -15892 -19988
rect -15828 -20052 -15808 -19988
rect -22107 -20068 -15808 -20052
rect -22107 -20132 -15892 -20068
rect -15828 -20132 -15808 -20068
rect -22107 -20148 -15808 -20132
rect -22107 -20212 -15892 -20148
rect -15828 -20212 -15808 -20148
rect -22107 -20228 -15808 -20212
rect -22107 -20292 -15892 -20228
rect -15828 -20292 -15808 -20228
rect -22107 -20308 -15808 -20292
rect -22107 -20372 -15892 -20308
rect -15828 -20372 -15808 -20308
rect -22107 -20388 -15808 -20372
rect -22107 -20452 -15892 -20388
rect -15828 -20452 -15808 -20388
rect -22107 -20468 -15808 -20452
rect -22107 -20532 -15892 -20468
rect -15828 -20532 -15808 -20468
rect -22107 -20548 -15808 -20532
rect -22107 -20612 -15892 -20548
rect -15828 -20612 -15808 -20548
rect -22107 -20628 -15808 -20612
rect -22107 -20692 -15892 -20628
rect -15828 -20692 -15808 -20628
rect -22107 -20708 -15808 -20692
rect -22107 -20772 -15892 -20708
rect -15828 -20772 -15808 -20708
rect -22107 -20788 -15808 -20772
rect -22107 -20852 -15892 -20788
rect -15828 -20852 -15808 -20788
rect -22107 -20868 -15808 -20852
rect -22107 -20932 -15892 -20868
rect -15828 -20932 -15808 -20868
rect -22107 -20948 -15808 -20932
rect -22107 -21012 -15892 -20948
rect -15828 -21012 -15808 -20948
rect -22107 -21028 -15808 -21012
rect -22107 -21092 -15892 -21028
rect -15828 -21092 -15808 -21028
rect -22107 -21108 -15808 -21092
rect -22107 -21172 -15892 -21108
rect -15828 -21172 -15808 -21108
rect -22107 -21188 -15808 -21172
rect -22107 -21252 -15892 -21188
rect -15828 -21252 -15808 -21188
rect -22107 -21268 -15808 -21252
rect -22107 -21332 -15892 -21268
rect -15828 -21332 -15808 -21268
rect -22107 -21348 -15808 -21332
rect -22107 -21412 -15892 -21348
rect -15828 -21412 -15808 -21348
rect -22107 -21428 -15808 -21412
rect -22107 -21492 -15892 -21428
rect -15828 -21492 -15808 -21428
rect -22107 -21508 -15808 -21492
rect -22107 -21572 -15892 -21508
rect -15828 -21572 -15808 -21508
rect -22107 -21588 -15808 -21572
rect -22107 -21652 -15892 -21588
rect -15828 -21652 -15808 -21588
rect -22107 -21668 -15808 -21652
rect -22107 -21732 -15892 -21668
rect -15828 -21732 -15808 -21668
rect -22107 -21748 -15808 -21732
rect -22107 -21812 -15892 -21748
rect -15828 -21812 -15808 -21748
rect -22107 -21828 -15808 -21812
rect -22107 -21892 -15892 -21828
rect -15828 -21892 -15808 -21828
rect -22107 -21908 -15808 -21892
rect -22107 -21972 -15892 -21908
rect -15828 -21972 -15808 -21908
rect -22107 -22000 -15808 -21972
rect -15788 -15828 -9489 -15800
rect -15788 -15892 -9573 -15828
rect -9509 -15892 -9489 -15828
rect -15788 -15908 -9489 -15892
rect -15788 -15972 -9573 -15908
rect -9509 -15972 -9489 -15908
rect -15788 -15988 -9489 -15972
rect -15788 -16052 -9573 -15988
rect -9509 -16052 -9489 -15988
rect -15788 -16068 -9489 -16052
rect -15788 -16132 -9573 -16068
rect -9509 -16132 -9489 -16068
rect -15788 -16148 -9489 -16132
rect -15788 -16212 -9573 -16148
rect -9509 -16212 -9489 -16148
rect -15788 -16228 -9489 -16212
rect -15788 -16292 -9573 -16228
rect -9509 -16292 -9489 -16228
rect -15788 -16308 -9489 -16292
rect -15788 -16372 -9573 -16308
rect -9509 -16372 -9489 -16308
rect -15788 -16388 -9489 -16372
rect -15788 -16452 -9573 -16388
rect -9509 -16452 -9489 -16388
rect -15788 -16468 -9489 -16452
rect -15788 -16532 -9573 -16468
rect -9509 -16532 -9489 -16468
rect -15788 -16548 -9489 -16532
rect -15788 -16612 -9573 -16548
rect -9509 -16612 -9489 -16548
rect -15788 -16628 -9489 -16612
rect -15788 -16692 -9573 -16628
rect -9509 -16692 -9489 -16628
rect -15788 -16708 -9489 -16692
rect -15788 -16772 -9573 -16708
rect -9509 -16772 -9489 -16708
rect -15788 -16788 -9489 -16772
rect -15788 -16852 -9573 -16788
rect -9509 -16852 -9489 -16788
rect -15788 -16868 -9489 -16852
rect -15788 -16932 -9573 -16868
rect -9509 -16932 -9489 -16868
rect -15788 -16948 -9489 -16932
rect -15788 -17012 -9573 -16948
rect -9509 -17012 -9489 -16948
rect -15788 -17028 -9489 -17012
rect -15788 -17092 -9573 -17028
rect -9509 -17092 -9489 -17028
rect -15788 -17108 -9489 -17092
rect -15788 -17172 -9573 -17108
rect -9509 -17172 -9489 -17108
rect -15788 -17188 -9489 -17172
rect -15788 -17252 -9573 -17188
rect -9509 -17252 -9489 -17188
rect -15788 -17268 -9489 -17252
rect -15788 -17332 -9573 -17268
rect -9509 -17332 -9489 -17268
rect -15788 -17348 -9489 -17332
rect -15788 -17412 -9573 -17348
rect -9509 -17412 -9489 -17348
rect -15788 -17428 -9489 -17412
rect -15788 -17492 -9573 -17428
rect -9509 -17492 -9489 -17428
rect -15788 -17508 -9489 -17492
rect -15788 -17572 -9573 -17508
rect -9509 -17572 -9489 -17508
rect -15788 -17588 -9489 -17572
rect -15788 -17652 -9573 -17588
rect -9509 -17652 -9489 -17588
rect -15788 -17668 -9489 -17652
rect -15788 -17732 -9573 -17668
rect -9509 -17732 -9489 -17668
rect -15788 -17748 -9489 -17732
rect -15788 -17812 -9573 -17748
rect -9509 -17812 -9489 -17748
rect -15788 -17828 -9489 -17812
rect -15788 -17892 -9573 -17828
rect -9509 -17892 -9489 -17828
rect -15788 -17908 -9489 -17892
rect -15788 -17972 -9573 -17908
rect -9509 -17972 -9489 -17908
rect -15788 -17988 -9489 -17972
rect -15788 -18052 -9573 -17988
rect -9509 -18052 -9489 -17988
rect -15788 -18068 -9489 -18052
rect -15788 -18132 -9573 -18068
rect -9509 -18132 -9489 -18068
rect -15788 -18148 -9489 -18132
rect -15788 -18212 -9573 -18148
rect -9509 -18212 -9489 -18148
rect -15788 -18228 -9489 -18212
rect -15788 -18292 -9573 -18228
rect -9509 -18292 -9489 -18228
rect -15788 -18308 -9489 -18292
rect -15788 -18372 -9573 -18308
rect -9509 -18372 -9489 -18308
rect -15788 -18388 -9489 -18372
rect -15788 -18452 -9573 -18388
rect -9509 -18452 -9489 -18388
rect -15788 -18468 -9489 -18452
rect -15788 -18532 -9573 -18468
rect -9509 -18532 -9489 -18468
rect -15788 -18548 -9489 -18532
rect -15788 -18612 -9573 -18548
rect -9509 -18612 -9489 -18548
rect -15788 -18628 -9489 -18612
rect -15788 -18692 -9573 -18628
rect -9509 -18692 -9489 -18628
rect -15788 -18708 -9489 -18692
rect -15788 -18772 -9573 -18708
rect -9509 -18772 -9489 -18708
rect -15788 -18788 -9489 -18772
rect -15788 -18852 -9573 -18788
rect -9509 -18852 -9489 -18788
rect -15788 -18868 -9489 -18852
rect -15788 -18932 -9573 -18868
rect -9509 -18932 -9489 -18868
rect -15788 -18948 -9489 -18932
rect -15788 -19012 -9573 -18948
rect -9509 -19012 -9489 -18948
rect -15788 -19028 -9489 -19012
rect -15788 -19092 -9573 -19028
rect -9509 -19092 -9489 -19028
rect -15788 -19108 -9489 -19092
rect -15788 -19172 -9573 -19108
rect -9509 -19172 -9489 -19108
rect -15788 -19188 -9489 -19172
rect -15788 -19252 -9573 -19188
rect -9509 -19252 -9489 -19188
rect -15788 -19268 -9489 -19252
rect -15788 -19332 -9573 -19268
rect -9509 -19332 -9489 -19268
rect -15788 -19348 -9489 -19332
rect -15788 -19412 -9573 -19348
rect -9509 -19412 -9489 -19348
rect -15788 -19428 -9489 -19412
rect -15788 -19492 -9573 -19428
rect -9509 -19492 -9489 -19428
rect -15788 -19508 -9489 -19492
rect -15788 -19572 -9573 -19508
rect -9509 -19572 -9489 -19508
rect -15788 -19588 -9489 -19572
rect -15788 -19652 -9573 -19588
rect -9509 -19652 -9489 -19588
rect -15788 -19668 -9489 -19652
rect -15788 -19732 -9573 -19668
rect -9509 -19732 -9489 -19668
rect -15788 -19748 -9489 -19732
rect -15788 -19812 -9573 -19748
rect -9509 -19812 -9489 -19748
rect -15788 -19828 -9489 -19812
rect -15788 -19892 -9573 -19828
rect -9509 -19892 -9489 -19828
rect -15788 -19908 -9489 -19892
rect -15788 -19972 -9573 -19908
rect -9509 -19972 -9489 -19908
rect -15788 -19988 -9489 -19972
rect -15788 -20052 -9573 -19988
rect -9509 -20052 -9489 -19988
rect -15788 -20068 -9489 -20052
rect -15788 -20132 -9573 -20068
rect -9509 -20132 -9489 -20068
rect -15788 -20148 -9489 -20132
rect -15788 -20212 -9573 -20148
rect -9509 -20212 -9489 -20148
rect -15788 -20228 -9489 -20212
rect -15788 -20292 -9573 -20228
rect -9509 -20292 -9489 -20228
rect -15788 -20308 -9489 -20292
rect -15788 -20372 -9573 -20308
rect -9509 -20372 -9489 -20308
rect -15788 -20388 -9489 -20372
rect -15788 -20452 -9573 -20388
rect -9509 -20452 -9489 -20388
rect -15788 -20468 -9489 -20452
rect -15788 -20532 -9573 -20468
rect -9509 -20532 -9489 -20468
rect -15788 -20548 -9489 -20532
rect -15788 -20612 -9573 -20548
rect -9509 -20612 -9489 -20548
rect -15788 -20628 -9489 -20612
rect -15788 -20692 -9573 -20628
rect -9509 -20692 -9489 -20628
rect -15788 -20708 -9489 -20692
rect -15788 -20772 -9573 -20708
rect -9509 -20772 -9489 -20708
rect -15788 -20788 -9489 -20772
rect -15788 -20852 -9573 -20788
rect -9509 -20852 -9489 -20788
rect -15788 -20868 -9489 -20852
rect -15788 -20932 -9573 -20868
rect -9509 -20932 -9489 -20868
rect -15788 -20948 -9489 -20932
rect -15788 -21012 -9573 -20948
rect -9509 -21012 -9489 -20948
rect -15788 -21028 -9489 -21012
rect -15788 -21092 -9573 -21028
rect -9509 -21092 -9489 -21028
rect -15788 -21108 -9489 -21092
rect -15788 -21172 -9573 -21108
rect -9509 -21172 -9489 -21108
rect -15788 -21188 -9489 -21172
rect -15788 -21252 -9573 -21188
rect -9509 -21252 -9489 -21188
rect -15788 -21268 -9489 -21252
rect -15788 -21332 -9573 -21268
rect -9509 -21332 -9489 -21268
rect -15788 -21348 -9489 -21332
rect -15788 -21412 -9573 -21348
rect -9509 -21412 -9489 -21348
rect -15788 -21428 -9489 -21412
rect -15788 -21492 -9573 -21428
rect -9509 -21492 -9489 -21428
rect -15788 -21508 -9489 -21492
rect -15788 -21572 -9573 -21508
rect -9509 -21572 -9489 -21508
rect -15788 -21588 -9489 -21572
rect -15788 -21652 -9573 -21588
rect -9509 -21652 -9489 -21588
rect -15788 -21668 -9489 -21652
rect -15788 -21732 -9573 -21668
rect -9509 -21732 -9489 -21668
rect -15788 -21748 -9489 -21732
rect -15788 -21812 -9573 -21748
rect -9509 -21812 -9489 -21748
rect -15788 -21828 -9489 -21812
rect -15788 -21892 -9573 -21828
rect -9509 -21892 -9489 -21828
rect -15788 -21908 -9489 -21892
rect -15788 -21972 -9573 -21908
rect -9509 -21972 -9489 -21908
rect -15788 -22000 -9489 -21972
rect -9469 -15828 -3170 -15800
rect -9469 -15892 -3254 -15828
rect -3190 -15892 -3170 -15828
rect -9469 -15908 -3170 -15892
rect -9469 -15972 -3254 -15908
rect -3190 -15972 -3170 -15908
rect -9469 -15988 -3170 -15972
rect -9469 -16052 -3254 -15988
rect -3190 -16052 -3170 -15988
rect -9469 -16068 -3170 -16052
rect -9469 -16132 -3254 -16068
rect -3190 -16132 -3170 -16068
rect -9469 -16148 -3170 -16132
rect -9469 -16212 -3254 -16148
rect -3190 -16212 -3170 -16148
rect -9469 -16228 -3170 -16212
rect -9469 -16292 -3254 -16228
rect -3190 -16292 -3170 -16228
rect -9469 -16308 -3170 -16292
rect -9469 -16372 -3254 -16308
rect -3190 -16372 -3170 -16308
rect -9469 -16388 -3170 -16372
rect -9469 -16452 -3254 -16388
rect -3190 -16452 -3170 -16388
rect -9469 -16468 -3170 -16452
rect -9469 -16532 -3254 -16468
rect -3190 -16532 -3170 -16468
rect -9469 -16548 -3170 -16532
rect -9469 -16612 -3254 -16548
rect -3190 -16612 -3170 -16548
rect -9469 -16628 -3170 -16612
rect -9469 -16692 -3254 -16628
rect -3190 -16692 -3170 -16628
rect -9469 -16708 -3170 -16692
rect -9469 -16772 -3254 -16708
rect -3190 -16772 -3170 -16708
rect -9469 -16788 -3170 -16772
rect -9469 -16852 -3254 -16788
rect -3190 -16852 -3170 -16788
rect -9469 -16868 -3170 -16852
rect -9469 -16932 -3254 -16868
rect -3190 -16932 -3170 -16868
rect -9469 -16948 -3170 -16932
rect -9469 -17012 -3254 -16948
rect -3190 -17012 -3170 -16948
rect -9469 -17028 -3170 -17012
rect -9469 -17092 -3254 -17028
rect -3190 -17092 -3170 -17028
rect -9469 -17108 -3170 -17092
rect -9469 -17172 -3254 -17108
rect -3190 -17172 -3170 -17108
rect -9469 -17188 -3170 -17172
rect -9469 -17252 -3254 -17188
rect -3190 -17252 -3170 -17188
rect -9469 -17268 -3170 -17252
rect -9469 -17332 -3254 -17268
rect -3190 -17332 -3170 -17268
rect -9469 -17348 -3170 -17332
rect -9469 -17412 -3254 -17348
rect -3190 -17412 -3170 -17348
rect -9469 -17428 -3170 -17412
rect -9469 -17492 -3254 -17428
rect -3190 -17492 -3170 -17428
rect -9469 -17508 -3170 -17492
rect -9469 -17572 -3254 -17508
rect -3190 -17572 -3170 -17508
rect -9469 -17588 -3170 -17572
rect -9469 -17652 -3254 -17588
rect -3190 -17652 -3170 -17588
rect -9469 -17668 -3170 -17652
rect -9469 -17732 -3254 -17668
rect -3190 -17732 -3170 -17668
rect -9469 -17748 -3170 -17732
rect -9469 -17812 -3254 -17748
rect -3190 -17812 -3170 -17748
rect -9469 -17828 -3170 -17812
rect -9469 -17892 -3254 -17828
rect -3190 -17892 -3170 -17828
rect -9469 -17908 -3170 -17892
rect -9469 -17972 -3254 -17908
rect -3190 -17972 -3170 -17908
rect -9469 -17988 -3170 -17972
rect -9469 -18052 -3254 -17988
rect -3190 -18052 -3170 -17988
rect -9469 -18068 -3170 -18052
rect -9469 -18132 -3254 -18068
rect -3190 -18132 -3170 -18068
rect -9469 -18148 -3170 -18132
rect -9469 -18212 -3254 -18148
rect -3190 -18212 -3170 -18148
rect -9469 -18228 -3170 -18212
rect -9469 -18292 -3254 -18228
rect -3190 -18292 -3170 -18228
rect -9469 -18308 -3170 -18292
rect -9469 -18372 -3254 -18308
rect -3190 -18372 -3170 -18308
rect -9469 -18388 -3170 -18372
rect -9469 -18452 -3254 -18388
rect -3190 -18452 -3170 -18388
rect -9469 -18468 -3170 -18452
rect -9469 -18532 -3254 -18468
rect -3190 -18532 -3170 -18468
rect -9469 -18548 -3170 -18532
rect -9469 -18612 -3254 -18548
rect -3190 -18612 -3170 -18548
rect -9469 -18628 -3170 -18612
rect -9469 -18692 -3254 -18628
rect -3190 -18692 -3170 -18628
rect -9469 -18708 -3170 -18692
rect -9469 -18772 -3254 -18708
rect -3190 -18772 -3170 -18708
rect -9469 -18788 -3170 -18772
rect -9469 -18852 -3254 -18788
rect -3190 -18852 -3170 -18788
rect -9469 -18868 -3170 -18852
rect -9469 -18932 -3254 -18868
rect -3190 -18932 -3170 -18868
rect -9469 -18948 -3170 -18932
rect -9469 -19012 -3254 -18948
rect -3190 -19012 -3170 -18948
rect -9469 -19028 -3170 -19012
rect -9469 -19092 -3254 -19028
rect -3190 -19092 -3170 -19028
rect -9469 -19108 -3170 -19092
rect -9469 -19172 -3254 -19108
rect -3190 -19172 -3170 -19108
rect -9469 -19188 -3170 -19172
rect -9469 -19252 -3254 -19188
rect -3190 -19252 -3170 -19188
rect -9469 -19268 -3170 -19252
rect -9469 -19332 -3254 -19268
rect -3190 -19332 -3170 -19268
rect -9469 -19348 -3170 -19332
rect -9469 -19412 -3254 -19348
rect -3190 -19412 -3170 -19348
rect -9469 -19428 -3170 -19412
rect -9469 -19492 -3254 -19428
rect -3190 -19492 -3170 -19428
rect -9469 -19508 -3170 -19492
rect -9469 -19572 -3254 -19508
rect -3190 -19572 -3170 -19508
rect -9469 -19588 -3170 -19572
rect -9469 -19652 -3254 -19588
rect -3190 -19652 -3170 -19588
rect -9469 -19668 -3170 -19652
rect -9469 -19732 -3254 -19668
rect -3190 -19732 -3170 -19668
rect -9469 -19748 -3170 -19732
rect -9469 -19812 -3254 -19748
rect -3190 -19812 -3170 -19748
rect -9469 -19828 -3170 -19812
rect -9469 -19892 -3254 -19828
rect -3190 -19892 -3170 -19828
rect -9469 -19908 -3170 -19892
rect -9469 -19972 -3254 -19908
rect -3190 -19972 -3170 -19908
rect -9469 -19988 -3170 -19972
rect -9469 -20052 -3254 -19988
rect -3190 -20052 -3170 -19988
rect -9469 -20068 -3170 -20052
rect -9469 -20132 -3254 -20068
rect -3190 -20132 -3170 -20068
rect -9469 -20148 -3170 -20132
rect -9469 -20212 -3254 -20148
rect -3190 -20212 -3170 -20148
rect -9469 -20228 -3170 -20212
rect -9469 -20292 -3254 -20228
rect -3190 -20292 -3170 -20228
rect -9469 -20308 -3170 -20292
rect -9469 -20372 -3254 -20308
rect -3190 -20372 -3170 -20308
rect -9469 -20388 -3170 -20372
rect -9469 -20452 -3254 -20388
rect -3190 -20452 -3170 -20388
rect -9469 -20468 -3170 -20452
rect -9469 -20532 -3254 -20468
rect -3190 -20532 -3170 -20468
rect -9469 -20548 -3170 -20532
rect -9469 -20612 -3254 -20548
rect -3190 -20612 -3170 -20548
rect -9469 -20628 -3170 -20612
rect -9469 -20692 -3254 -20628
rect -3190 -20692 -3170 -20628
rect -9469 -20708 -3170 -20692
rect -9469 -20772 -3254 -20708
rect -3190 -20772 -3170 -20708
rect -9469 -20788 -3170 -20772
rect -9469 -20852 -3254 -20788
rect -3190 -20852 -3170 -20788
rect -9469 -20868 -3170 -20852
rect -9469 -20932 -3254 -20868
rect -3190 -20932 -3170 -20868
rect -9469 -20948 -3170 -20932
rect -9469 -21012 -3254 -20948
rect -3190 -21012 -3170 -20948
rect -9469 -21028 -3170 -21012
rect -9469 -21092 -3254 -21028
rect -3190 -21092 -3170 -21028
rect -9469 -21108 -3170 -21092
rect -9469 -21172 -3254 -21108
rect -3190 -21172 -3170 -21108
rect -9469 -21188 -3170 -21172
rect -9469 -21252 -3254 -21188
rect -3190 -21252 -3170 -21188
rect -9469 -21268 -3170 -21252
rect -9469 -21332 -3254 -21268
rect -3190 -21332 -3170 -21268
rect -9469 -21348 -3170 -21332
rect -9469 -21412 -3254 -21348
rect -3190 -21412 -3170 -21348
rect -9469 -21428 -3170 -21412
rect -9469 -21492 -3254 -21428
rect -3190 -21492 -3170 -21428
rect -9469 -21508 -3170 -21492
rect -9469 -21572 -3254 -21508
rect -3190 -21572 -3170 -21508
rect -9469 -21588 -3170 -21572
rect -9469 -21652 -3254 -21588
rect -3190 -21652 -3170 -21588
rect -9469 -21668 -3170 -21652
rect -9469 -21732 -3254 -21668
rect -3190 -21732 -3170 -21668
rect -9469 -21748 -3170 -21732
rect -9469 -21812 -3254 -21748
rect -3190 -21812 -3170 -21748
rect -9469 -21828 -3170 -21812
rect -9469 -21892 -3254 -21828
rect -3190 -21892 -3170 -21828
rect -9469 -21908 -3170 -21892
rect -9469 -21972 -3254 -21908
rect -3190 -21972 -3170 -21908
rect -9469 -22000 -3170 -21972
rect -3150 -15828 3149 -15800
rect -3150 -15892 3065 -15828
rect 3129 -15892 3149 -15828
rect -3150 -15908 3149 -15892
rect -3150 -15972 3065 -15908
rect 3129 -15972 3149 -15908
rect -3150 -15988 3149 -15972
rect -3150 -16052 3065 -15988
rect 3129 -16052 3149 -15988
rect -3150 -16068 3149 -16052
rect -3150 -16132 3065 -16068
rect 3129 -16132 3149 -16068
rect -3150 -16148 3149 -16132
rect -3150 -16212 3065 -16148
rect 3129 -16212 3149 -16148
rect -3150 -16228 3149 -16212
rect -3150 -16292 3065 -16228
rect 3129 -16292 3149 -16228
rect -3150 -16308 3149 -16292
rect -3150 -16372 3065 -16308
rect 3129 -16372 3149 -16308
rect -3150 -16388 3149 -16372
rect -3150 -16452 3065 -16388
rect 3129 -16452 3149 -16388
rect -3150 -16468 3149 -16452
rect -3150 -16532 3065 -16468
rect 3129 -16532 3149 -16468
rect -3150 -16548 3149 -16532
rect -3150 -16612 3065 -16548
rect 3129 -16612 3149 -16548
rect -3150 -16628 3149 -16612
rect -3150 -16692 3065 -16628
rect 3129 -16692 3149 -16628
rect -3150 -16708 3149 -16692
rect -3150 -16772 3065 -16708
rect 3129 -16772 3149 -16708
rect -3150 -16788 3149 -16772
rect -3150 -16852 3065 -16788
rect 3129 -16852 3149 -16788
rect -3150 -16868 3149 -16852
rect -3150 -16932 3065 -16868
rect 3129 -16932 3149 -16868
rect -3150 -16948 3149 -16932
rect -3150 -17012 3065 -16948
rect 3129 -17012 3149 -16948
rect -3150 -17028 3149 -17012
rect -3150 -17092 3065 -17028
rect 3129 -17092 3149 -17028
rect -3150 -17108 3149 -17092
rect -3150 -17172 3065 -17108
rect 3129 -17172 3149 -17108
rect -3150 -17188 3149 -17172
rect -3150 -17252 3065 -17188
rect 3129 -17252 3149 -17188
rect -3150 -17268 3149 -17252
rect -3150 -17332 3065 -17268
rect 3129 -17332 3149 -17268
rect -3150 -17348 3149 -17332
rect -3150 -17412 3065 -17348
rect 3129 -17412 3149 -17348
rect -3150 -17428 3149 -17412
rect -3150 -17492 3065 -17428
rect 3129 -17492 3149 -17428
rect -3150 -17508 3149 -17492
rect -3150 -17572 3065 -17508
rect 3129 -17572 3149 -17508
rect -3150 -17588 3149 -17572
rect -3150 -17652 3065 -17588
rect 3129 -17652 3149 -17588
rect -3150 -17668 3149 -17652
rect -3150 -17732 3065 -17668
rect 3129 -17732 3149 -17668
rect -3150 -17748 3149 -17732
rect -3150 -17812 3065 -17748
rect 3129 -17812 3149 -17748
rect -3150 -17828 3149 -17812
rect -3150 -17892 3065 -17828
rect 3129 -17892 3149 -17828
rect -3150 -17908 3149 -17892
rect -3150 -17972 3065 -17908
rect 3129 -17972 3149 -17908
rect -3150 -17988 3149 -17972
rect -3150 -18052 3065 -17988
rect 3129 -18052 3149 -17988
rect -3150 -18068 3149 -18052
rect -3150 -18132 3065 -18068
rect 3129 -18132 3149 -18068
rect -3150 -18148 3149 -18132
rect -3150 -18212 3065 -18148
rect 3129 -18212 3149 -18148
rect -3150 -18228 3149 -18212
rect -3150 -18292 3065 -18228
rect 3129 -18292 3149 -18228
rect -3150 -18308 3149 -18292
rect -3150 -18372 3065 -18308
rect 3129 -18372 3149 -18308
rect -3150 -18388 3149 -18372
rect -3150 -18452 3065 -18388
rect 3129 -18452 3149 -18388
rect -3150 -18468 3149 -18452
rect -3150 -18532 3065 -18468
rect 3129 -18532 3149 -18468
rect -3150 -18548 3149 -18532
rect -3150 -18612 3065 -18548
rect 3129 -18612 3149 -18548
rect -3150 -18628 3149 -18612
rect -3150 -18692 3065 -18628
rect 3129 -18692 3149 -18628
rect -3150 -18708 3149 -18692
rect -3150 -18772 3065 -18708
rect 3129 -18772 3149 -18708
rect -3150 -18788 3149 -18772
rect -3150 -18852 3065 -18788
rect 3129 -18852 3149 -18788
rect -3150 -18868 3149 -18852
rect -3150 -18932 3065 -18868
rect 3129 -18932 3149 -18868
rect -3150 -18948 3149 -18932
rect -3150 -19012 3065 -18948
rect 3129 -19012 3149 -18948
rect -3150 -19028 3149 -19012
rect -3150 -19092 3065 -19028
rect 3129 -19092 3149 -19028
rect -3150 -19108 3149 -19092
rect -3150 -19172 3065 -19108
rect 3129 -19172 3149 -19108
rect -3150 -19188 3149 -19172
rect -3150 -19252 3065 -19188
rect 3129 -19252 3149 -19188
rect -3150 -19268 3149 -19252
rect -3150 -19332 3065 -19268
rect 3129 -19332 3149 -19268
rect -3150 -19348 3149 -19332
rect -3150 -19412 3065 -19348
rect 3129 -19412 3149 -19348
rect -3150 -19428 3149 -19412
rect -3150 -19492 3065 -19428
rect 3129 -19492 3149 -19428
rect -3150 -19508 3149 -19492
rect -3150 -19572 3065 -19508
rect 3129 -19572 3149 -19508
rect -3150 -19588 3149 -19572
rect -3150 -19652 3065 -19588
rect 3129 -19652 3149 -19588
rect -3150 -19668 3149 -19652
rect -3150 -19732 3065 -19668
rect 3129 -19732 3149 -19668
rect -3150 -19748 3149 -19732
rect -3150 -19812 3065 -19748
rect 3129 -19812 3149 -19748
rect -3150 -19828 3149 -19812
rect -3150 -19892 3065 -19828
rect 3129 -19892 3149 -19828
rect -3150 -19908 3149 -19892
rect -3150 -19972 3065 -19908
rect 3129 -19972 3149 -19908
rect -3150 -19988 3149 -19972
rect -3150 -20052 3065 -19988
rect 3129 -20052 3149 -19988
rect -3150 -20068 3149 -20052
rect -3150 -20132 3065 -20068
rect 3129 -20132 3149 -20068
rect -3150 -20148 3149 -20132
rect -3150 -20212 3065 -20148
rect 3129 -20212 3149 -20148
rect -3150 -20228 3149 -20212
rect -3150 -20292 3065 -20228
rect 3129 -20292 3149 -20228
rect -3150 -20308 3149 -20292
rect -3150 -20372 3065 -20308
rect 3129 -20372 3149 -20308
rect -3150 -20388 3149 -20372
rect -3150 -20452 3065 -20388
rect 3129 -20452 3149 -20388
rect -3150 -20468 3149 -20452
rect -3150 -20532 3065 -20468
rect 3129 -20532 3149 -20468
rect -3150 -20548 3149 -20532
rect -3150 -20612 3065 -20548
rect 3129 -20612 3149 -20548
rect -3150 -20628 3149 -20612
rect -3150 -20692 3065 -20628
rect 3129 -20692 3149 -20628
rect -3150 -20708 3149 -20692
rect -3150 -20772 3065 -20708
rect 3129 -20772 3149 -20708
rect -3150 -20788 3149 -20772
rect -3150 -20852 3065 -20788
rect 3129 -20852 3149 -20788
rect -3150 -20868 3149 -20852
rect -3150 -20932 3065 -20868
rect 3129 -20932 3149 -20868
rect -3150 -20948 3149 -20932
rect -3150 -21012 3065 -20948
rect 3129 -21012 3149 -20948
rect -3150 -21028 3149 -21012
rect -3150 -21092 3065 -21028
rect 3129 -21092 3149 -21028
rect -3150 -21108 3149 -21092
rect -3150 -21172 3065 -21108
rect 3129 -21172 3149 -21108
rect -3150 -21188 3149 -21172
rect -3150 -21252 3065 -21188
rect 3129 -21252 3149 -21188
rect -3150 -21268 3149 -21252
rect -3150 -21332 3065 -21268
rect 3129 -21332 3149 -21268
rect -3150 -21348 3149 -21332
rect -3150 -21412 3065 -21348
rect 3129 -21412 3149 -21348
rect -3150 -21428 3149 -21412
rect -3150 -21492 3065 -21428
rect 3129 -21492 3149 -21428
rect -3150 -21508 3149 -21492
rect -3150 -21572 3065 -21508
rect 3129 -21572 3149 -21508
rect -3150 -21588 3149 -21572
rect -3150 -21652 3065 -21588
rect 3129 -21652 3149 -21588
rect -3150 -21668 3149 -21652
rect -3150 -21732 3065 -21668
rect 3129 -21732 3149 -21668
rect -3150 -21748 3149 -21732
rect -3150 -21812 3065 -21748
rect 3129 -21812 3149 -21748
rect -3150 -21828 3149 -21812
rect -3150 -21892 3065 -21828
rect 3129 -21892 3149 -21828
rect -3150 -21908 3149 -21892
rect -3150 -21972 3065 -21908
rect 3129 -21972 3149 -21908
rect -3150 -22000 3149 -21972
rect 3169 -15828 9468 -15800
rect 3169 -15892 9384 -15828
rect 9448 -15892 9468 -15828
rect 3169 -15908 9468 -15892
rect 3169 -15972 9384 -15908
rect 9448 -15972 9468 -15908
rect 3169 -15988 9468 -15972
rect 3169 -16052 9384 -15988
rect 9448 -16052 9468 -15988
rect 3169 -16068 9468 -16052
rect 3169 -16132 9384 -16068
rect 9448 -16132 9468 -16068
rect 3169 -16148 9468 -16132
rect 3169 -16212 9384 -16148
rect 9448 -16212 9468 -16148
rect 3169 -16228 9468 -16212
rect 3169 -16292 9384 -16228
rect 9448 -16292 9468 -16228
rect 3169 -16308 9468 -16292
rect 3169 -16372 9384 -16308
rect 9448 -16372 9468 -16308
rect 3169 -16388 9468 -16372
rect 3169 -16452 9384 -16388
rect 9448 -16452 9468 -16388
rect 3169 -16468 9468 -16452
rect 3169 -16532 9384 -16468
rect 9448 -16532 9468 -16468
rect 3169 -16548 9468 -16532
rect 3169 -16612 9384 -16548
rect 9448 -16612 9468 -16548
rect 3169 -16628 9468 -16612
rect 3169 -16692 9384 -16628
rect 9448 -16692 9468 -16628
rect 3169 -16708 9468 -16692
rect 3169 -16772 9384 -16708
rect 9448 -16772 9468 -16708
rect 3169 -16788 9468 -16772
rect 3169 -16852 9384 -16788
rect 9448 -16852 9468 -16788
rect 3169 -16868 9468 -16852
rect 3169 -16932 9384 -16868
rect 9448 -16932 9468 -16868
rect 3169 -16948 9468 -16932
rect 3169 -17012 9384 -16948
rect 9448 -17012 9468 -16948
rect 3169 -17028 9468 -17012
rect 3169 -17092 9384 -17028
rect 9448 -17092 9468 -17028
rect 3169 -17108 9468 -17092
rect 3169 -17172 9384 -17108
rect 9448 -17172 9468 -17108
rect 3169 -17188 9468 -17172
rect 3169 -17252 9384 -17188
rect 9448 -17252 9468 -17188
rect 3169 -17268 9468 -17252
rect 3169 -17332 9384 -17268
rect 9448 -17332 9468 -17268
rect 3169 -17348 9468 -17332
rect 3169 -17412 9384 -17348
rect 9448 -17412 9468 -17348
rect 3169 -17428 9468 -17412
rect 3169 -17492 9384 -17428
rect 9448 -17492 9468 -17428
rect 3169 -17508 9468 -17492
rect 3169 -17572 9384 -17508
rect 9448 -17572 9468 -17508
rect 3169 -17588 9468 -17572
rect 3169 -17652 9384 -17588
rect 9448 -17652 9468 -17588
rect 3169 -17668 9468 -17652
rect 3169 -17732 9384 -17668
rect 9448 -17732 9468 -17668
rect 3169 -17748 9468 -17732
rect 3169 -17812 9384 -17748
rect 9448 -17812 9468 -17748
rect 3169 -17828 9468 -17812
rect 3169 -17892 9384 -17828
rect 9448 -17892 9468 -17828
rect 3169 -17908 9468 -17892
rect 3169 -17972 9384 -17908
rect 9448 -17972 9468 -17908
rect 3169 -17988 9468 -17972
rect 3169 -18052 9384 -17988
rect 9448 -18052 9468 -17988
rect 3169 -18068 9468 -18052
rect 3169 -18132 9384 -18068
rect 9448 -18132 9468 -18068
rect 3169 -18148 9468 -18132
rect 3169 -18212 9384 -18148
rect 9448 -18212 9468 -18148
rect 3169 -18228 9468 -18212
rect 3169 -18292 9384 -18228
rect 9448 -18292 9468 -18228
rect 3169 -18308 9468 -18292
rect 3169 -18372 9384 -18308
rect 9448 -18372 9468 -18308
rect 3169 -18388 9468 -18372
rect 3169 -18452 9384 -18388
rect 9448 -18452 9468 -18388
rect 3169 -18468 9468 -18452
rect 3169 -18532 9384 -18468
rect 9448 -18532 9468 -18468
rect 3169 -18548 9468 -18532
rect 3169 -18612 9384 -18548
rect 9448 -18612 9468 -18548
rect 3169 -18628 9468 -18612
rect 3169 -18692 9384 -18628
rect 9448 -18692 9468 -18628
rect 3169 -18708 9468 -18692
rect 3169 -18772 9384 -18708
rect 9448 -18772 9468 -18708
rect 3169 -18788 9468 -18772
rect 3169 -18852 9384 -18788
rect 9448 -18852 9468 -18788
rect 3169 -18868 9468 -18852
rect 3169 -18932 9384 -18868
rect 9448 -18932 9468 -18868
rect 3169 -18948 9468 -18932
rect 3169 -19012 9384 -18948
rect 9448 -19012 9468 -18948
rect 3169 -19028 9468 -19012
rect 3169 -19092 9384 -19028
rect 9448 -19092 9468 -19028
rect 3169 -19108 9468 -19092
rect 3169 -19172 9384 -19108
rect 9448 -19172 9468 -19108
rect 3169 -19188 9468 -19172
rect 3169 -19252 9384 -19188
rect 9448 -19252 9468 -19188
rect 3169 -19268 9468 -19252
rect 3169 -19332 9384 -19268
rect 9448 -19332 9468 -19268
rect 3169 -19348 9468 -19332
rect 3169 -19412 9384 -19348
rect 9448 -19412 9468 -19348
rect 3169 -19428 9468 -19412
rect 3169 -19492 9384 -19428
rect 9448 -19492 9468 -19428
rect 3169 -19508 9468 -19492
rect 3169 -19572 9384 -19508
rect 9448 -19572 9468 -19508
rect 3169 -19588 9468 -19572
rect 3169 -19652 9384 -19588
rect 9448 -19652 9468 -19588
rect 3169 -19668 9468 -19652
rect 3169 -19732 9384 -19668
rect 9448 -19732 9468 -19668
rect 3169 -19748 9468 -19732
rect 3169 -19812 9384 -19748
rect 9448 -19812 9468 -19748
rect 3169 -19828 9468 -19812
rect 3169 -19892 9384 -19828
rect 9448 -19892 9468 -19828
rect 3169 -19908 9468 -19892
rect 3169 -19972 9384 -19908
rect 9448 -19972 9468 -19908
rect 3169 -19988 9468 -19972
rect 3169 -20052 9384 -19988
rect 9448 -20052 9468 -19988
rect 3169 -20068 9468 -20052
rect 3169 -20132 9384 -20068
rect 9448 -20132 9468 -20068
rect 3169 -20148 9468 -20132
rect 3169 -20212 9384 -20148
rect 9448 -20212 9468 -20148
rect 3169 -20228 9468 -20212
rect 3169 -20292 9384 -20228
rect 9448 -20292 9468 -20228
rect 3169 -20308 9468 -20292
rect 3169 -20372 9384 -20308
rect 9448 -20372 9468 -20308
rect 3169 -20388 9468 -20372
rect 3169 -20452 9384 -20388
rect 9448 -20452 9468 -20388
rect 3169 -20468 9468 -20452
rect 3169 -20532 9384 -20468
rect 9448 -20532 9468 -20468
rect 3169 -20548 9468 -20532
rect 3169 -20612 9384 -20548
rect 9448 -20612 9468 -20548
rect 3169 -20628 9468 -20612
rect 3169 -20692 9384 -20628
rect 9448 -20692 9468 -20628
rect 3169 -20708 9468 -20692
rect 3169 -20772 9384 -20708
rect 9448 -20772 9468 -20708
rect 3169 -20788 9468 -20772
rect 3169 -20852 9384 -20788
rect 9448 -20852 9468 -20788
rect 3169 -20868 9468 -20852
rect 3169 -20932 9384 -20868
rect 9448 -20932 9468 -20868
rect 3169 -20948 9468 -20932
rect 3169 -21012 9384 -20948
rect 9448 -21012 9468 -20948
rect 3169 -21028 9468 -21012
rect 3169 -21092 9384 -21028
rect 9448 -21092 9468 -21028
rect 3169 -21108 9468 -21092
rect 3169 -21172 9384 -21108
rect 9448 -21172 9468 -21108
rect 3169 -21188 9468 -21172
rect 3169 -21252 9384 -21188
rect 9448 -21252 9468 -21188
rect 3169 -21268 9468 -21252
rect 3169 -21332 9384 -21268
rect 9448 -21332 9468 -21268
rect 3169 -21348 9468 -21332
rect 3169 -21412 9384 -21348
rect 9448 -21412 9468 -21348
rect 3169 -21428 9468 -21412
rect 3169 -21492 9384 -21428
rect 9448 -21492 9468 -21428
rect 3169 -21508 9468 -21492
rect 3169 -21572 9384 -21508
rect 9448 -21572 9468 -21508
rect 3169 -21588 9468 -21572
rect 3169 -21652 9384 -21588
rect 9448 -21652 9468 -21588
rect 3169 -21668 9468 -21652
rect 3169 -21732 9384 -21668
rect 9448 -21732 9468 -21668
rect 3169 -21748 9468 -21732
rect 3169 -21812 9384 -21748
rect 9448 -21812 9468 -21748
rect 3169 -21828 9468 -21812
rect 3169 -21892 9384 -21828
rect 9448 -21892 9468 -21828
rect 3169 -21908 9468 -21892
rect 3169 -21972 9384 -21908
rect 9448 -21972 9468 -21908
rect 3169 -22000 9468 -21972
rect 9488 -15828 15787 -15800
rect 9488 -15892 15703 -15828
rect 15767 -15892 15787 -15828
rect 9488 -15908 15787 -15892
rect 9488 -15972 15703 -15908
rect 15767 -15972 15787 -15908
rect 9488 -15988 15787 -15972
rect 9488 -16052 15703 -15988
rect 15767 -16052 15787 -15988
rect 9488 -16068 15787 -16052
rect 9488 -16132 15703 -16068
rect 15767 -16132 15787 -16068
rect 9488 -16148 15787 -16132
rect 9488 -16212 15703 -16148
rect 15767 -16212 15787 -16148
rect 9488 -16228 15787 -16212
rect 9488 -16292 15703 -16228
rect 15767 -16292 15787 -16228
rect 9488 -16308 15787 -16292
rect 9488 -16372 15703 -16308
rect 15767 -16372 15787 -16308
rect 9488 -16388 15787 -16372
rect 9488 -16452 15703 -16388
rect 15767 -16452 15787 -16388
rect 9488 -16468 15787 -16452
rect 9488 -16532 15703 -16468
rect 15767 -16532 15787 -16468
rect 9488 -16548 15787 -16532
rect 9488 -16612 15703 -16548
rect 15767 -16612 15787 -16548
rect 9488 -16628 15787 -16612
rect 9488 -16692 15703 -16628
rect 15767 -16692 15787 -16628
rect 9488 -16708 15787 -16692
rect 9488 -16772 15703 -16708
rect 15767 -16772 15787 -16708
rect 9488 -16788 15787 -16772
rect 9488 -16852 15703 -16788
rect 15767 -16852 15787 -16788
rect 9488 -16868 15787 -16852
rect 9488 -16932 15703 -16868
rect 15767 -16932 15787 -16868
rect 9488 -16948 15787 -16932
rect 9488 -17012 15703 -16948
rect 15767 -17012 15787 -16948
rect 9488 -17028 15787 -17012
rect 9488 -17092 15703 -17028
rect 15767 -17092 15787 -17028
rect 9488 -17108 15787 -17092
rect 9488 -17172 15703 -17108
rect 15767 -17172 15787 -17108
rect 9488 -17188 15787 -17172
rect 9488 -17252 15703 -17188
rect 15767 -17252 15787 -17188
rect 9488 -17268 15787 -17252
rect 9488 -17332 15703 -17268
rect 15767 -17332 15787 -17268
rect 9488 -17348 15787 -17332
rect 9488 -17412 15703 -17348
rect 15767 -17412 15787 -17348
rect 9488 -17428 15787 -17412
rect 9488 -17492 15703 -17428
rect 15767 -17492 15787 -17428
rect 9488 -17508 15787 -17492
rect 9488 -17572 15703 -17508
rect 15767 -17572 15787 -17508
rect 9488 -17588 15787 -17572
rect 9488 -17652 15703 -17588
rect 15767 -17652 15787 -17588
rect 9488 -17668 15787 -17652
rect 9488 -17732 15703 -17668
rect 15767 -17732 15787 -17668
rect 9488 -17748 15787 -17732
rect 9488 -17812 15703 -17748
rect 15767 -17812 15787 -17748
rect 9488 -17828 15787 -17812
rect 9488 -17892 15703 -17828
rect 15767 -17892 15787 -17828
rect 9488 -17908 15787 -17892
rect 9488 -17972 15703 -17908
rect 15767 -17972 15787 -17908
rect 9488 -17988 15787 -17972
rect 9488 -18052 15703 -17988
rect 15767 -18052 15787 -17988
rect 9488 -18068 15787 -18052
rect 9488 -18132 15703 -18068
rect 15767 -18132 15787 -18068
rect 9488 -18148 15787 -18132
rect 9488 -18212 15703 -18148
rect 15767 -18212 15787 -18148
rect 9488 -18228 15787 -18212
rect 9488 -18292 15703 -18228
rect 15767 -18292 15787 -18228
rect 9488 -18308 15787 -18292
rect 9488 -18372 15703 -18308
rect 15767 -18372 15787 -18308
rect 9488 -18388 15787 -18372
rect 9488 -18452 15703 -18388
rect 15767 -18452 15787 -18388
rect 9488 -18468 15787 -18452
rect 9488 -18532 15703 -18468
rect 15767 -18532 15787 -18468
rect 9488 -18548 15787 -18532
rect 9488 -18612 15703 -18548
rect 15767 -18612 15787 -18548
rect 9488 -18628 15787 -18612
rect 9488 -18692 15703 -18628
rect 15767 -18692 15787 -18628
rect 9488 -18708 15787 -18692
rect 9488 -18772 15703 -18708
rect 15767 -18772 15787 -18708
rect 9488 -18788 15787 -18772
rect 9488 -18852 15703 -18788
rect 15767 -18852 15787 -18788
rect 9488 -18868 15787 -18852
rect 9488 -18932 15703 -18868
rect 15767 -18932 15787 -18868
rect 9488 -18948 15787 -18932
rect 9488 -19012 15703 -18948
rect 15767 -19012 15787 -18948
rect 9488 -19028 15787 -19012
rect 9488 -19092 15703 -19028
rect 15767 -19092 15787 -19028
rect 9488 -19108 15787 -19092
rect 9488 -19172 15703 -19108
rect 15767 -19172 15787 -19108
rect 9488 -19188 15787 -19172
rect 9488 -19252 15703 -19188
rect 15767 -19252 15787 -19188
rect 9488 -19268 15787 -19252
rect 9488 -19332 15703 -19268
rect 15767 -19332 15787 -19268
rect 9488 -19348 15787 -19332
rect 9488 -19412 15703 -19348
rect 15767 -19412 15787 -19348
rect 9488 -19428 15787 -19412
rect 9488 -19492 15703 -19428
rect 15767 -19492 15787 -19428
rect 9488 -19508 15787 -19492
rect 9488 -19572 15703 -19508
rect 15767 -19572 15787 -19508
rect 9488 -19588 15787 -19572
rect 9488 -19652 15703 -19588
rect 15767 -19652 15787 -19588
rect 9488 -19668 15787 -19652
rect 9488 -19732 15703 -19668
rect 15767 -19732 15787 -19668
rect 9488 -19748 15787 -19732
rect 9488 -19812 15703 -19748
rect 15767 -19812 15787 -19748
rect 9488 -19828 15787 -19812
rect 9488 -19892 15703 -19828
rect 15767 -19892 15787 -19828
rect 9488 -19908 15787 -19892
rect 9488 -19972 15703 -19908
rect 15767 -19972 15787 -19908
rect 9488 -19988 15787 -19972
rect 9488 -20052 15703 -19988
rect 15767 -20052 15787 -19988
rect 9488 -20068 15787 -20052
rect 9488 -20132 15703 -20068
rect 15767 -20132 15787 -20068
rect 9488 -20148 15787 -20132
rect 9488 -20212 15703 -20148
rect 15767 -20212 15787 -20148
rect 9488 -20228 15787 -20212
rect 9488 -20292 15703 -20228
rect 15767 -20292 15787 -20228
rect 9488 -20308 15787 -20292
rect 9488 -20372 15703 -20308
rect 15767 -20372 15787 -20308
rect 9488 -20388 15787 -20372
rect 9488 -20452 15703 -20388
rect 15767 -20452 15787 -20388
rect 9488 -20468 15787 -20452
rect 9488 -20532 15703 -20468
rect 15767 -20532 15787 -20468
rect 9488 -20548 15787 -20532
rect 9488 -20612 15703 -20548
rect 15767 -20612 15787 -20548
rect 9488 -20628 15787 -20612
rect 9488 -20692 15703 -20628
rect 15767 -20692 15787 -20628
rect 9488 -20708 15787 -20692
rect 9488 -20772 15703 -20708
rect 15767 -20772 15787 -20708
rect 9488 -20788 15787 -20772
rect 9488 -20852 15703 -20788
rect 15767 -20852 15787 -20788
rect 9488 -20868 15787 -20852
rect 9488 -20932 15703 -20868
rect 15767 -20932 15787 -20868
rect 9488 -20948 15787 -20932
rect 9488 -21012 15703 -20948
rect 15767 -21012 15787 -20948
rect 9488 -21028 15787 -21012
rect 9488 -21092 15703 -21028
rect 15767 -21092 15787 -21028
rect 9488 -21108 15787 -21092
rect 9488 -21172 15703 -21108
rect 15767 -21172 15787 -21108
rect 9488 -21188 15787 -21172
rect 9488 -21252 15703 -21188
rect 15767 -21252 15787 -21188
rect 9488 -21268 15787 -21252
rect 9488 -21332 15703 -21268
rect 15767 -21332 15787 -21268
rect 9488 -21348 15787 -21332
rect 9488 -21412 15703 -21348
rect 15767 -21412 15787 -21348
rect 9488 -21428 15787 -21412
rect 9488 -21492 15703 -21428
rect 15767 -21492 15787 -21428
rect 9488 -21508 15787 -21492
rect 9488 -21572 15703 -21508
rect 15767 -21572 15787 -21508
rect 9488 -21588 15787 -21572
rect 9488 -21652 15703 -21588
rect 15767 -21652 15787 -21588
rect 9488 -21668 15787 -21652
rect 9488 -21732 15703 -21668
rect 15767 -21732 15787 -21668
rect 9488 -21748 15787 -21732
rect 9488 -21812 15703 -21748
rect 15767 -21812 15787 -21748
rect 9488 -21828 15787 -21812
rect 9488 -21892 15703 -21828
rect 15767 -21892 15787 -21828
rect 9488 -21908 15787 -21892
rect 9488 -21972 15703 -21908
rect 15767 -21972 15787 -21908
rect 9488 -22000 15787 -21972
rect 15807 -15828 22106 -15800
rect 15807 -15892 22022 -15828
rect 22086 -15892 22106 -15828
rect 15807 -15908 22106 -15892
rect 15807 -15972 22022 -15908
rect 22086 -15972 22106 -15908
rect 15807 -15988 22106 -15972
rect 15807 -16052 22022 -15988
rect 22086 -16052 22106 -15988
rect 15807 -16068 22106 -16052
rect 15807 -16132 22022 -16068
rect 22086 -16132 22106 -16068
rect 15807 -16148 22106 -16132
rect 15807 -16212 22022 -16148
rect 22086 -16212 22106 -16148
rect 15807 -16228 22106 -16212
rect 15807 -16292 22022 -16228
rect 22086 -16292 22106 -16228
rect 15807 -16308 22106 -16292
rect 15807 -16372 22022 -16308
rect 22086 -16372 22106 -16308
rect 15807 -16388 22106 -16372
rect 15807 -16452 22022 -16388
rect 22086 -16452 22106 -16388
rect 15807 -16468 22106 -16452
rect 15807 -16532 22022 -16468
rect 22086 -16532 22106 -16468
rect 15807 -16548 22106 -16532
rect 15807 -16612 22022 -16548
rect 22086 -16612 22106 -16548
rect 15807 -16628 22106 -16612
rect 15807 -16692 22022 -16628
rect 22086 -16692 22106 -16628
rect 15807 -16708 22106 -16692
rect 15807 -16772 22022 -16708
rect 22086 -16772 22106 -16708
rect 15807 -16788 22106 -16772
rect 15807 -16852 22022 -16788
rect 22086 -16852 22106 -16788
rect 15807 -16868 22106 -16852
rect 15807 -16932 22022 -16868
rect 22086 -16932 22106 -16868
rect 15807 -16948 22106 -16932
rect 15807 -17012 22022 -16948
rect 22086 -17012 22106 -16948
rect 15807 -17028 22106 -17012
rect 15807 -17092 22022 -17028
rect 22086 -17092 22106 -17028
rect 15807 -17108 22106 -17092
rect 15807 -17172 22022 -17108
rect 22086 -17172 22106 -17108
rect 15807 -17188 22106 -17172
rect 15807 -17252 22022 -17188
rect 22086 -17252 22106 -17188
rect 15807 -17268 22106 -17252
rect 15807 -17332 22022 -17268
rect 22086 -17332 22106 -17268
rect 15807 -17348 22106 -17332
rect 15807 -17412 22022 -17348
rect 22086 -17412 22106 -17348
rect 15807 -17428 22106 -17412
rect 15807 -17492 22022 -17428
rect 22086 -17492 22106 -17428
rect 15807 -17508 22106 -17492
rect 15807 -17572 22022 -17508
rect 22086 -17572 22106 -17508
rect 15807 -17588 22106 -17572
rect 15807 -17652 22022 -17588
rect 22086 -17652 22106 -17588
rect 15807 -17668 22106 -17652
rect 15807 -17732 22022 -17668
rect 22086 -17732 22106 -17668
rect 15807 -17748 22106 -17732
rect 15807 -17812 22022 -17748
rect 22086 -17812 22106 -17748
rect 15807 -17828 22106 -17812
rect 15807 -17892 22022 -17828
rect 22086 -17892 22106 -17828
rect 15807 -17908 22106 -17892
rect 15807 -17972 22022 -17908
rect 22086 -17972 22106 -17908
rect 15807 -17988 22106 -17972
rect 15807 -18052 22022 -17988
rect 22086 -18052 22106 -17988
rect 15807 -18068 22106 -18052
rect 15807 -18132 22022 -18068
rect 22086 -18132 22106 -18068
rect 15807 -18148 22106 -18132
rect 15807 -18212 22022 -18148
rect 22086 -18212 22106 -18148
rect 15807 -18228 22106 -18212
rect 15807 -18292 22022 -18228
rect 22086 -18292 22106 -18228
rect 15807 -18308 22106 -18292
rect 15807 -18372 22022 -18308
rect 22086 -18372 22106 -18308
rect 15807 -18388 22106 -18372
rect 15807 -18452 22022 -18388
rect 22086 -18452 22106 -18388
rect 15807 -18468 22106 -18452
rect 15807 -18532 22022 -18468
rect 22086 -18532 22106 -18468
rect 15807 -18548 22106 -18532
rect 15807 -18612 22022 -18548
rect 22086 -18612 22106 -18548
rect 15807 -18628 22106 -18612
rect 15807 -18692 22022 -18628
rect 22086 -18692 22106 -18628
rect 15807 -18708 22106 -18692
rect 15807 -18772 22022 -18708
rect 22086 -18772 22106 -18708
rect 15807 -18788 22106 -18772
rect 15807 -18852 22022 -18788
rect 22086 -18852 22106 -18788
rect 15807 -18868 22106 -18852
rect 15807 -18932 22022 -18868
rect 22086 -18932 22106 -18868
rect 15807 -18948 22106 -18932
rect 15807 -19012 22022 -18948
rect 22086 -19012 22106 -18948
rect 15807 -19028 22106 -19012
rect 15807 -19092 22022 -19028
rect 22086 -19092 22106 -19028
rect 15807 -19108 22106 -19092
rect 15807 -19172 22022 -19108
rect 22086 -19172 22106 -19108
rect 15807 -19188 22106 -19172
rect 15807 -19252 22022 -19188
rect 22086 -19252 22106 -19188
rect 15807 -19268 22106 -19252
rect 15807 -19332 22022 -19268
rect 22086 -19332 22106 -19268
rect 15807 -19348 22106 -19332
rect 15807 -19412 22022 -19348
rect 22086 -19412 22106 -19348
rect 15807 -19428 22106 -19412
rect 15807 -19492 22022 -19428
rect 22086 -19492 22106 -19428
rect 15807 -19508 22106 -19492
rect 15807 -19572 22022 -19508
rect 22086 -19572 22106 -19508
rect 15807 -19588 22106 -19572
rect 15807 -19652 22022 -19588
rect 22086 -19652 22106 -19588
rect 15807 -19668 22106 -19652
rect 15807 -19732 22022 -19668
rect 22086 -19732 22106 -19668
rect 15807 -19748 22106 -19732
rect 15807 -19812 22022 -19748
rect 22086 -19812 22106 -19748
rect 15807 -19828 22106 -19812
rect 15807 -19892 22022 -19828
rect 22086 -19892 22106 -19828
rect 15807 -19908 22106 -19892
rect 15807 -19972 22022 -19908
rect 22086 -19972 22106 -19908
rect 15807 -19988 22106 -19972
rect 15807 -20052 22022 -19988
rect 22086 -20052 22106 -19988
rect 15807 -20068 22106 -20052
rect 15807 -20132 22022 -20068
rect 22086 -20132 22106 -20068
rect 15807 -20148 22106 -20132
rect 15807 -20212 22022 -20148
rect 22086 -20212 22106 -20148
rect 15807 -20228 22106 -20212
rect 15807 -20292 22022 -20228
rect 22086 -20292 22106 -20228
rect 15807 -20308 22106 -20292
rect 15807 -20372 22022 -20308
rect 22086 -20372 22106 -20308
rect 15807 -20388 22106 -20372
rect 15807 -20452 22022 -20388
rect 22086 -20452 22106 -20388
rect 15807 -20468 22106 -20452
rect 15807 -20532 22022 -20468
rect 22086 -20532 22106 -20468
rect 15807 -20548 22106 -20532
rect 15807 -20612 22022 -20548
rect 22086 -20612 22106 -20548
rect 15807 -20628 22106 -20612
rect 15807 -20692 22022 -20628
rect 22086 -20692 22106 -20628
rect 15807 -20708 22106 -20692
rect 15807 -20772 22022 -20708
rect 22086 -20772 22106 -20708
rect 15807 -20788 22106 -20772
rect 15807 -20852 22022 -20788
rect 22086 -20852 22106 -20788
rect 15807 -20868 22106 -20852
rect 15807 -20932 22022 -20868
rect 22086 -20932 22106 -20868
rect 15807 -20948 22106 -20932
rect 15807 -21012 22022 -20948
rect 22086 -21012 22106 -20948
rect 15807 -21028 22106 -21012
rect 15807 -21092 22022 -21028
rect 22086 -21092 22106 -21028
rect 15807 -21108 22106 -21092
rect 15807 -21172 22022 -21108
rect 22086 -21172 22106 -21108
rect 15807 -21188 22106 -21172
rect 15807 -21252 22022 -21188
rect 22086 -21252 22106 -21188
rect 15807 -21268 22106 -21252
rect 15807 -21332 22022 -21268
rect 22086 -21332 22106 -21268
rect 15807 -21348 22106 -21332
rect 15807 -21412 22022 -21348
rect 22086 -21412 22106 -21348
rect 15807 -21428 22106 -21412
rect 15807 -21492 22022 -21428
rect 22086 -21492 22106 -21428
rect 15807 -21508 22106 -21492
rect 15807 -21572 22022 -21508
rect 22086 -21572 22106 -21508
rect 15807 -21588 22106 -21572
rect 15807 -21652 22022 -21588
rect 22086 -21652 22106 -21588
rect 15807 -21668 22106 -21652
rect 15807 -21732 22022 -21668
rect 22086 -21732 22106 -21668
rect 15807 -21748 22106 -21732
rect 15807 -21812 22022 -21748
rect 22086 -21812 22106 -21748
rect 15807 -21828 22106 -21812
rect 15807 -21892 22022 -21828
rect 22086 -21892 22106 -21828
rect 15807 -21908 22106 -21892
rect 15807 -21972 22022 -21908
rect 22086 -21972 22106 -21908
rect 15807 -22000 22106 -21972
rect 22126 -15828 28425 -15800
rect 22126 -15892 28341 -15828
rect 28405 -15892 28425 -15828
rect 22126 -15908 28425 -15892
rect 22126 -15972 28341 -15908
rect 28405 -15972 28425 -15908
rect 22126 -15988 28425 -15972
rect 22126 -16052 28341 -15988
rect 28405 -16052 28425 -15988
rect 22126 -16068 28425 -16052
rect 22126 -16132 28341 -16068
rect 28405 -16132 28425 -16068
rect 22126 -16148 28425 -16132
rect 22126 -16212 28341 -16148
rect 28405 -16212 28425 -16148
rect 22126 -16228 28425 -16212
rect 22126 -16292 28341 -16228
rect 28405 -16292 28425 -16228
rect 22126 -16308 28425 -16292
rect 22126 -16372 28341 -16308
rect 28405 -16372 28425 -16308
rect 22126 -16388 28425 -16372
rect 22126 -16452 28341 -16388
rect 28405 -16452 28425 -16388
rect 22126 -16468 28425 -16452
rect 22126 -16532 28341 -16468
rect 28405 -16532 28425 -16468
rect 22126 -16548 28425 -16532
rect 22126 -16612 28341 -16548
rect 28405 -16612 28425 -16548
rect 22126 -16628 28425 -16612
rect 22126 -16692 28341 -16628
rect 28405 -16692 28425 -16628
rect 22126 -16708 28425 -16692
rect 22126 -16772 28341 -16708
rect 28405 -16772 28425 -16708
rect 22126 -16788 28425 -16772
rect 22126 -16852 28341 -16788
rect 28405 -16852 28425 -16788
rect 22126 -16868 28425 -16852
rect 22126 -16932 28341 -16868
rect 28405 -16932 28425 -16868
rect 22126 -16948 28425 -16932
rect 22126 -17012 28341 -16948
rect 28405 -17012 28425 -16948
rect 22126 -17028 28425 -17012
rect 22126 -17092 28341 -17028
rect 28405 -17092 28425 -17028
rect 22126 -17108 28425 -17092
rect 22126 -17172 28341 -17108
rect 28405 -17172 28425 -17108
rect 22126 -17188 28425 -17172
rect 22126 -17252 28341 -17188
rect 28405 -17252 28425 -17188
rect 22126 -17268 28425 -17252
rect 22126 -17332 28341 -17268
rect 28405 -17332 28425 -17268
rect 22126 -17348 28425 -17332
rect 22126 -17412 28341 -17348
rect 28405 -17412 28425 -17348
rect 22126 -17428 28425 -17412
rect 22126 -17492 28341 -17428
rect 28405 -17492 28425 -17428
rect 22126 -17508 28425 -17492
rect 22126 -17572 28341 -17508
rect 28405 -17572 28425 -17508
rect 22126 -17588 28425 -17572
rect 22126 -17652 28341 -17588
rect 28405 -17652 28425 -17588
rect 22126 -17668 28425 -17652
rect 22126 -17732 28341 -17668
rect 28405 -17732 28425 -17668
rect 22126 -17748 28425 -17732
rect 22126 -17812 28341 -17748
rect 28405 -17812 28425 -17748
rect 22126 -17828 28425 -17812
rect 22126 -17892 28341 -17828
rect 28405 -17892 28425 -17828
rect 22126 -17908 28425 -17892
rect 22126 -17972 28341 -17908
rect 28405 -17972 28425 -17908
rect 22126 -17988 28425 -17972
rect 22126 -18052 28341 -17988
rect 28405 -18052 28425 -17988
rect 22126 -18068 28425 -18052
rect 22126 -18132 28341 -18068
rect 28405 -18132 28425 -18068
rect 22126 -18148 28425 -18132
rect 22126 -18212 28341 -18148
rect 28405 -18212 28425 -18148
rect 22126 -18228 28425 -18212
rect 22126 -18292 28341 -18228
rect 28405 -18292 28425 -18228
rect 22126 -18308 28425 -18292
rect 22126 -18372 28341 -18308
rect 28405 -18372 28425 -18308
rect 22126 -18388 28425 -18372
rect 22126 -18452 28341 -18388
rect 28405 -18452 28425 -18388
rect 22126 -18468 28425 -18452
rect 22126 -18532 28341 -18468
rect 28405 -18532 28425 -18468
rect 22126 -18548 28425 -18532
rect 22126 -18612 28341 -18548
rect 28405 -18612 28425 -18548
rect 22126 -18628 28425 -18612
rect 22126 -18692 28341 -18628
rect 28405 -18692 28425 -18628
rect 22126 -18708 28425 -18692
rect 22126 -18772 28341 -18708
rect 28405 -18772 28425 -18708
rect 22126 -18788 28425 -18772
rect 22126 -18852 28341 -18788
rect 28405 -18852 28425 -18788
rect 22126 -18868 28425 -18852
rect 22126 -18932 28341 -18868
rect 28405 -18932 28425 -18868
rect 22126 -18948 28425 -18932
rect 22126 -19012 28341 -18948
rect 28405 -19012 28425 -18948
rect 22126 -19028 28425 -19012
rect 22126 -19092 28341 -19028
rect 28405 -19092 28425 -19028
rect 22126 -19108 28425 -19092
rect 22126 -19172 28341 -19108
rect 28405 -19172 28425 -19108
rect 22126 -19188 28425 -19172
rect 22126 -19252 28341 -19188
rect 28405 -19252 28425 -19188
rect 22126 -19268 28425 -19252
rect 22126 -19332 28341 -19268
rect 28405 -19332 28425 -19268
rect 22126 -19348 28425 -19332
rect 22126 -19412 28341 -19348
rect 28405 -19412 28425 -19348
rect 22126 -19428 28425 -19412
rect 22126 -19492 28341 -19428
rect 28405 -19492 28425 -19428
rect 22126 -19508 28425 -19492
rect 22126 -19572 28341 -19508
rect 28405 -19572 28425 -19508
rect 22126 -19588 28425 -19572
rect 22126 -19652 28341 -19588
rect 28405 -19652 28425 -19588
rect 22126 -19668 28425 -19652
rect 22126 -19732 28341 -19668
rect 28405 -19732 28425 -19668
rect 22126 -19748 28425 -19732
rect 22126 -19812 28341 -19748
rect 28405 -19812 28425 -19748
rect 22126 -19828 28425 -19812
rect 22126 -19892 28341 -19828
rect 28405 -19892 28425 -19828
rect 22126 -19908 28425 -19892
rect 22126 -19972 28341 -19908
rect 28405 -19972 28425 -19908
rect 22126 -19988 28425 -19972
rect 22126 -20052 28341 -19988
rect 28405 -20052 28425 -19988
rect 22126 -20068 28425 -20052
rect 22126 -20132 28341 -20068
rect 28405 -20132 28425 -20068
rect 22126 -20148 28425 -20132
rect 22126 -20212 28341 -20148
rect 28405 -20212 28425 -20148
rect 22126 -20228 28425 -20212
rect 22126 -20292 28341 -20228
rect 28405 -20292 28425 -20228
rect 22126 -20308 28425 -20292
rect 22126 -20372 28341 -20308
rect 28405 -20372 28425 -20308
rect 22126 -20388 28425 -20372
rect 22126 -20452 28341 -20388
rect 28405 -20452 28425 -20388
rect 22126 -20468 28425 -20452
rect 22126 -20532 28341 -20468
rect 28405 -20532 28425 -20468
rect 22126 -20548 28425 -20532
rect 22126 -20612 28341 -20548
rect 28405 -20612 28425 -20548
rect 22126 -20628 28425 -20612
rect 22126 -20692 28341 -20628
rect 28405 -20692 28425 -20628
rect 22126 -20708 28425 -20692
rect 22126 -20772 28341 -20708
rect 28405 -20772 28425 -20708
rect 22126 -20788 28425 -20772
rect 22126 -20852 28341 -20788
rect 28405 -20852 28425 -20788
rect 22126 -20868 28425 -20852
rect 22126 -20932 28341 -20868
rect 28405 -20932 28425 -20868
rect 22126 -20948 28425 -20932
rect 22126 -21012 28341 -20948
rect 28405 -21012 28425 -20948
rect 22126 -21028 28425 -21012
rect 22126 -21092 28341 -21028
rect 28405 -21092 28425 -21028
rect 22126 -21108 28425 -21092
rect 22126 -21172 28341 -21108
rect 28405 -21172 28425 -21108
rect 22126 -21188 28425 -21172
rect 22126 -21252 28341 -21188
rect 28405 -21252 28425 -21188
rect 22126 -21268 28425 -21252
rect 22126 -21332 28341 -21268
rect 28405 -21332 28425 -21268
rect 22126 -21348 28425 -21332
rect 22126 -21412 28341 -21348
rect 28405 -21412 28425 -21348
rect 22126 -21428 28425 -21412
rect 22126 -21492 28341 -21428
rect 28405 -21492 28425 -21428
rect 22126 -21508 28425 -21492
rect 22126 -21572 28341 -21508
rect 28405 -21572 28425 -21508
rect 22126 -21588 28425 -21572
rect 22126 -21652 28341 -21588
rect 28405 -21652 28425 -21588
rect 22126 -21668 28425 -21652
rect 22126 -21732 28341 -21668
rect 28405 -21732 28425 -21668
rect 22126 -21748 28425 -21732
rect 22126 -21812 28341 -21748
rect 28405 -21812 28425 -21748
rect 22126 -21828 28425 -21812
rect 22126 -21892 28341 -21828
rect 28405 -21892 28425 -21828
rect 22126 -21908 28425 -21892
rect 22126 -21972 28341 -21908
rect 28405 -21972 28425 -21908
rect 22126 -22000 28425 -21972
rect 28445 -15828 34744 -15800
rect 28445 -15892 34660 -15828
rect 34724 -15892 34744 -15828
rect 28445 -15908 34744 -15892
rect 28445 -15972 34660 -15908
rect 34724 -15972 34744 -15908
rect 28445 -15988 34744 -15972
rect 28445 -16052 34660 -15988
rect 34724 -16052 34744 -15988
rect 28445 -16068 34744 -16052
rect 28445 -16132 34660 -16068
rect 34724 -16132 34744 -16068
rect 28445 -16148 34744 -16132
rect 28445 -16212 34660 -16148
rect 34724 -16212 34744 -16148
rect 28445 -16228 34744 -16212
rect 28445 -16292 34660 -16228
rect 34724 -16292 34744 -16228
rect 28445 -16308 34744 -16292
rect 28445 -16372 34660 -16308
rect 34724 -16372 34744 -16308
rect 28445 -16388 34744 -16372
rect 28445 -16452 34660 -16388
rect 34724 -16452 34744 -16388
rect 28445 -16468 34744 -16452
rect 28445 -16532 34660 -16468
rect 34724 -16532 34744 -16468
rect 28445 -16548 34744 -16532
rect 28445 -16612 34660 -16548
rect 34724 -16612 34744 -16548
rect 28445 -16628 34744 -16612
rect 28445 -16692 34660 -16628
rect 34724 -16692 34744 -16628
rect 28445 -16708 34744 -16692
rect 28445 -16772 34660 -16708
rect 34724 -16772 34744 -16708
rect 28445 -16788 34744 -16772
rect 28445 -16852 34660 -16788
rect 34724 -16852 34744 -16788
rect 28445 -16868 34744 -16852
rect 28445 -16932 34660 -16868
rect 34724 -16932 34744 -16868
rect 28445 -16948 34744 -16932
rect 28445 -17012 34660 -16948
rect 34724 -17012 34744 -16948
rect 28445 -17028 34744 -17012
rect 28445 -17092 34660 -17028
rect 34724 -17092 34744 -17028
rect 28445 -17108 34744 -17092
rect 28445 -17172 34660 -17108
rect 34724 -17172 34744 -17108
rect 28445 -17188 34744 -17172
rect 28445 -17252 34660 -17188
rect 34724 -17252 34744 -17188
rect 28445 -17268 34744 -17252
rect 28445 -17332 34660 -17268
rect 34724 -17332 34744 -17268
rect 28445 -17348 34744 -17332
rect 28445 -17412 34660 -17348
rect 34724 -17412 34744 -17348
rect 28445 -17428 34744 -17412
rect 28445 -17492 34660 -17428
rect 34724 -17492 34744 -17428
rect 28445 -17508 34744 -17492
rect 28445 -17572 34660 -17508
rect 34724 -17572 34744 -17508
rect 28445 -17588 34744 -17572
rect 28445 -17652 34660 -17588
rect 34724 -17652 34744 -17588
rect 28445 -17668 34744 -17652
rect 28445 -17732 34660 -17668
rect 34724 -17732 34744 -17668
rect 28445 -17748 34744 -17732
rect 28445 -17812 34660 -17748
rect 34724 -17812 34744 -17748
rect 28445 -17828 34744 -17812
rect 28445 -17892 34660 -17828
rect 34724 -17892 34744 -17828
rect 28445 -17908 34744 -17892
rect 28445 -17972 34660 -17908
rect 34724 -17972 34744 -17908
rect 28445 -17988 34744 -17972
rect 28445 -18052 34660 -17988
rect 34724 -18052 34744 -17988
rect 28445 -18068 34744 -18052
rect 28445 -18132 34660 -18068
rect 34724 -18132 34744 -18068
rect 28445 -18148 34744 -18132
rect 28445 -18212 34660 -18148
rect 34724 -18212 34744 -18148
rect 28445 -18228 34744 -18212
rect 28445 -18292 34660 -18228
rect 34724 -18292 34744 -18228
rect 28445 -18308 34744 -18292
rect 28445 -18372 34660 -18308
rect 34724 -18372 34744 -18308
rect 28445 -18388 34744 -18372
rect 28445 -18452 34660 -18388
rect 34724 -18452 34744 -18388
rect 28445 -18468 34744 -18452
rect 28445 -18532 34660 -18468
rect 34724 -18532 34744 -18468
rect 28445 -18548 34744 -18532
rect 28445 -18612 34660 -18548
rect 34724 -18612 34744 -18548
rect 28445 -18628 34744 -18612
rect 28445 -18692 34660 -18628
rect 34724 -18692 34744 -18628
rect 28445 -18708 34744 -18692
rect 28445 -18772 34660 -18708
rect 34724 -18772 34744 -18708
rect 28445 -18788 34744 -18772
rect 28445 -18852 34660 -18788
rect 34724 -18852 34744 -18788
rect 28445 -18868 34744 -18852
rect 28445 -18932 34660 -18868
rect 34724 -18932 34744 -18868
rect 28445 -18948 34744 -18932
rect 28445 -19012 34660 -18948
rect 34724 -19012 34744 -18948
rect 28445 -19028 34744 -19012
rect 28445 -19092 34660 -19028
rect 34724 -19092 34744 -19028
rect 28445 -19108 34744 -19092
rect 28445 -19172 34660 -19108
rect 34724 -19172 34744 -19108
rect 28445 -19188 34744 -19172
rect 28445 -19252 34660 -19188
rect 34724 -19252 34744 -19188
rect 28445 -19268 34744 -19252
rect 28445 -19332 34660 -19268
rect 34724 -19332 34744 -19268
rect 28445 -19348 34744 -19332
rect 28445 -19412 34660 -19348
rect 34724 -19412 34744 -19348
rect 28445 -19428 34744 -19412
rect 28445 -19492 34660 -19428
rect 34724 -19492 34744 -19428
rect 28445 -19508 34744 -19492
rect 28445 -19572 34660 -19508
rect 34724 -19572 34744 -19508
rect 28445 -19588 34744 -19572
rect 28445 -19652 34660 -19588
rect 34724 -19652 34744 -19588
rect 28445 -19668 34744 -19652
rect 28445 -19732 34660 -19668
rect 34724 -19732 34744 -19668
rect 28445 -19748 34744 -19732
rect 28445 -19812 34660 -19748
rect 34724 -19812 34744 -19748
rect 28445 -19828 34744 -19812
rect 28445 -19892 34660 -19828
rect 34724 -19892 34744 -19828
rect 28445 -19908 34744 -19892
rect 28445 -19972 34660 -19908
rect 34724 -19972 34744 -19908
rect 28445 -19988 34744 -19972
rect 28445 -20052 34660 -19988
rect 34724 -20052 34744 -19988
rect 28445 -20068 34744 -20052
rect 28445 -20132 34660 -20068
rect 34724 -20132 34744 -20068
rect 28445 -20148 34744 -20132
rect 28445 -20212 34660 -20148
rect 34724 -20212 34744 -20148
rect 28445 -20228 34744 -20212
rect 28445 -20292 34660 -20228
rect 34724 -20292 34744 -20228
rect 28445 -20308 34744 -20292
rect 28445 -20372 34660 -20308
rect 34724 -20372 34744 -20308
rect 28445 -20388 34744 -20372
rect 28445 -20452 34660 -20388
rect 34724 -20452 34744 -20388
rect 28445 -20468 34744 -20452
rect 28445 -20532 34660 -20468
rect 34724 -20532 34744 -20468
rect 28445 -20548 34744 -20532
rect 28445 -20612 34660 -20548
rect 34724 -20612 34744 -20548
rect 28445 -20628 34744 -20612
rect 28445 -20692 34660 -20628
rect 34724 -20692 34744 -20628
rect 28445 -20708 34744 -20692
rect 28445 -20772 34660 -20708
rect 34724 -20772 34744 -20708
rect 28445 -20788 34744 -20772
rect 28445 -20852 34660 -20788
rect 34724 -20852 34744 -20788
rect 28445 -20868 34744 -20852
rect 28445 -20932 34660 -20868
rect 34724 -20932 34744 -20868
rect 28445 -20948 34744 -20932
rect 28445 -21012 34660 -20948
rect 34724 -21012 34744 -20948
rect 28445 -21028 34744 -21012
rect 28445 -21092 34660 -21028
rect 34724 -21092 34744 -21028
rect 28445 -21108 34744 -21092
rect 28445 -21172 34660 -21108
rect 34724 -21172 34744 -21108
rect 28445 -21188 34744 -21172
rect 28445 -21252 34660 -21188
rect 34724 -21252 34744 -21188
rect 28445 -21268 34744 -21252
rect 28445 -21332 34660 -21268
rect 34724 -21332 34744 -21268
rect 28445 -21348 34744 -21332
rect 28445 -21412 34660 -21348
rect 34724 -21412 34744 -21348
rect 28445 -21428 34744 -21412
rect 28445 -21492 34660 -21428
rect 34724 -21492 34744 -21428
rect 28445 -21508 34744 -21492
rect 28445 -21572 34660 -21508
rect 34724 -21572 34744 -21508
rect 28445 -21588 34744 -21572
rect 28445 -21652 34660 -21588
rect 34724 -21652 34744 -21588
rect 28445 -21668 34744 -21652
rect 28445 -21732 34660 -21668
rect 34724 -21732 34744 -21668
rect 28445 -21748 34744 -21732
rect 28445 -21812 34660 -21748
rect 34724 -21812 34744 -21748
rect 28445 -21828 34744 -21812
rect 28445 -21892 34660 -21828
rect 34724 -21892 34744 -21828
rect 28445 -21908 34744 -21892
rect 28445 -21972 34660 -21908
rect 34724 -21972 34744 -21908
rect 28445 -22000 34744 -21972
rect 34764 -15828 41063 -15800
rect 34764 -15892 40979 -15828
rect 41043 -15892 41063 -15828
rect 34764 -15908 41063 -15892
rect 34764 -15972 40979 -15908
rect 41043 -15972 41063 -15908
rect 34764 -15988 41063 -15972
rect 34764 -16052 40979 -15988
rect 41043 -16052 41063 -15988
rect 34764 -16068 41063 -16052
rect 34764 -16132 40979 -16068
rect 41043 -16132 41063 -16068
rect 34764 -16148 41063 -16132
rect 34764 -16212 40979 -16148
rect 41043 -16212 41063 -16148
rect 34764 -16228 41063 -16212
rect 34764 -16292 40979 -16228
rect 41043 -16292 41063 -16228
rect 34764 -16308 41063 -16292
rect 34764 -16372 40979 -16308
rect 41043 -16372 41063 -16308
rect 34764 -16388 41063 -16372
rect 34764 -16452 40979 -16388
rect 41043 -16452 41063 -16388
rect 34764 -16468 41063 -16452
rect 34764 -16532 40979 -16468
rect 41043 -16532 41063 -16468
rect 34764 -16548 41063 -16532
rect 34764 -16612 40979 -16548
rect 41043 -16612 41063 -16548
rect 34764 -16628 41063 -16612
rect 34764 -16692 40979 -16628
rect 41043 -16692 41063 -16628
rect 34764 -16708 41063 -16692
rect 34764 -16772 40979 -16708
rect 41043 -16772 41063 -16708
rect 34764 -16788 41063 -16772
rect 34764 -16852 40979 -16788
rect 41043 -16852 41063 -16788
rect 34764 -16868 41063 -16852
rect 34764 -16932 40979 -16868
rect 41043 -16932 41063 -16868
rect 34764 -16948 41063 -16932
rect 34764 -17012 40979 -16948
rect 41043 -17012 41063 -16948
rect 34764 -17028 41063 -17012
rect 34764 -17092 40979 -17028
rect 41043 -17092 41063 -17028
rect 34764 -17108 41063 -17092
rect 34764 -17172 40979 -17108
rect 41043 -17172 41063 -17108
rect 34764 -17188 41063 -17172
rect 34764 -17252 40979 -17188
rect 41043 -17252 41063 -17188
rect 34764 -17268 41063 -17252
rect 34764 -17332 40979 -17268
rect 41043 -17332 41063 -17268
rect 34764 -17348 41063 -17332
rect 34764 -17412 40979 -17348
rect 41043 -17412 41063 -17348
rect 34764 -17428 41063 -17412
rect 34764 -17492 40979 -17428
rect 41043 -17492 41063 -17428
rect 34764 -17508 41063 -17492
rect 34764 -17572 40979 -17508
rect 41043 -17572 41063 -17508
rect 34764 -17588 41063 -17572
rect 34764 -17652 40979 -17588
rect 41043 -17652 41063 -17588
rect 34764 -17668 41063 -17652
rect 34764 -17732 40979 -17668
rect 41043 -17732 41063 -17668
rect 34764 -17748 41063 -17732
rect 34764 -17812 40979 -17748
rect 41043 -17812 41063 -17748
rect 34764 -17828 41063 -17812
rect 34764 -17892 40979 -17828
rect 41043 -17892 41063 -17828
rect 34764 -17908 41063 -17892
rect 34764 -17972 40979 -17908
rect 41043 -17972 41063 -17908
rect 34764 -17988 41063 -17972
rect 34764 -18052 40979 -17988
rect 41043 -18052 41063 -17988
rect 34764 -18068 41063 -18052
rect 34764 -18132 40979 -18068
rect 41043 -18132 41063 -18068
rect 34764 -18148 41063 -18132
rect 34764 -18212 40979 -18148
rect 41043 -18212 41063 -18148
rect 34764 -18228 41063 -18212
rect 34764 -18292 40979 -18228
rect 41043 -18292 41063 -18228
rect 34764 -18308 41063 -18292
rect 34764 -18372 40979 -18308
rect 41043 -18372 41063 -18308
rect 34764 -18388 41063 -18372
rect 34764 -18452 40979 -18388
rect 41043 -18452 41063 -18388
rect 34764 -18468 41063 -18452
rect 34764 -18532 40979 -18468
rect 41043 -18532 41063 -18468
rect 34764 -18548 41063 -18532
rect 34764 -18612 40979 -18548
rect 41043 -18612 41063 -18548
rect 34764 -18628 41063 -18612
rect 34764 -18692 40979 -18628
rect 41043 -18692 41063 -18628
rect 34764 -18708 41063 -18692
rect 34764 -18772 40979 -18708
rect 41043 -18772 41063 -18708
rect 34764 -18788 41063 -18772
rect 34764 -18852 40979 -18788
rect 41043 -18852 41063 -18788
rect 34764 -18868 41063 -18852
rect 34764 -18932 40979 -18868
rect 41043 -18932 41063 -18868
rect 34764 -18948 41063 -18932
rect 34764 -19012 40979 -18948
rect 41043 -19012 41063 -18948
rect 34764 -19028 41063 -19012
rect 34764 -19092 40979 -19028
rect 41043 -19092 41063 -19028
rect 34764 -19108 41063 -19092
rect 34764 -19172 40979 -19108
rect 41043 -19172 41063 -19108
rect 34764 -19188 41063 -19172
rect 34764 -19252 40979 -19188
rect 41043 -19252 41063 -19188
rect 34764 -19268 41063 -19252
rect 34764 -19332 40979 -19268
rect 41043 -19332 41063 -19268
rect 34764 -19348 41063 -19332
rect 34764 -19412 40979 -19348
rect 41043 -19412 41063 -19348
rect 34764 -19428 41063 -19412
rect 34764 -19492 40979 -19428
rect 41043 -19492 41063 -19428
rect 34764 -19508 41063 -19492
rect 34764 -19572 40979 -19508
rect 41043 -19572 41063 -19508
rect 34764 -19588 41063 -19572
rect 34764 -19652 40979 -19588
rect 41043 -19652 41063 -19588
rect 34764 -19668 41063 -19652
rect 34764 -19732 40979 -19668
rect 41043 -19732 41063 -19668
rect 34764 -19748 41063 -19732
rect 34764 -19812 40979 -19748
rect 41043 -19812 41063 -19748
rect 34764 -19828 41063 -19812
rect 34764 -19892 40979 -19828
rect 41043 -19892 41063 -19828
rect 34764 -19908 41063 -19892
rect 34764 -19972 40979 -19908
rect 41043 -19972 41063 -19908
rect 34764 -19988 41063 -19972
rect 34764 -20052 40979 -19988
rect 41043 -20052 41063 -19988
rect 34764 -20068 41063 -20052
rect 34764 -20132 40979 -20068
rect 41043 -20132 41063 -20068
rect 34764 -20148 41063 -20132
rect 34764 -20212 40979 -20148
rect 41043 -20212 41063 -20148
rect 34764 -20228 41063 -20212
rect 34764 -20292 40979 -20228
rect 41043 -20292 41063 -20228
rect 34764 -20308 41063 -20292
rect 34764 -20372 40979 -20308
rect 41043 -20372 41063 -20308
rect 34764 -20388 41063 -20372
rect 34764 -20452 40979 -20388
rect 41043 -20452 41063 -20388
rect 34764 -20468 41063 -20452
rect 34764 -20532 40979 -20468
rect 41043 -20532 41063 -20468
rect 34764 -20548 41063 -20532
rect 34764 -20612 40979 -20548
rect 41043 -20612 41063 -20548
rect 34764 -20628 41063 -20612
rect 34764 -20692 40979 -20628
rect 41043 -20692 41063 -20628
rect 34764 -20708 41063 -20692
rect 34764 -20772 40979 -20708
rect 41043 -20772 41063 -20708
rect 34764 -20788 41063 -20772
rect 34764 -20852 40979 -20788
rect 41043 -20852 41063 -20788
rect 34764 -20868 41063 -20852
rect 34764 -20932 40979 -20868
rect 41043 -20932 41063 -20868
rect 34764 -20948 41063 -20932
rect 34764 -21012 40979 -20948
rect 41043 -21012 41063 -20948
rect 34764 -21028 41063 -21012
rect 34764 -21092 40979 -21028
rect 41043 -21092 41063 -21028
rect 34764 -21108 41063 -21092
rect 34764 -21172 40979 -21108
rect 41043 -21172 41063 -21108
rect 34764 -21188 41063 -21172
rect 34764 -21252 40979 -21188
rect 41043 -21252 41063 -21188
rect 34764 -21268 41063 -21252
rect 34764 -21332 40979 -21268
rect 41043 -21332 41063 -21268
rect 34764 -21348 41063 -21332
rect 34764 -21412 40979 -21348
rect 41043 -21412 41063 -21348
rect 34764 -21428 41063 -21412
rect 34764 -21492 40979 -21428
rect 41043 -21492 41063 -21428
rect 34764 -21508 41063 -21492
rect 34764 -21572 40979 -21508
rect 41043 -21572 41063 -21508
rect 34764 -21588 41063 -21572
rect 34764 -21652 40979 -21588
rect 41043 -21652 41063 -21588
rect 34764 -21668 41063 -21652
rect 34764 -21732 40979 -21668
rect 41043 -21732 41063 -21668
rect 34764 -21748 41063 -21732
rect 34764 -21812 40979 -21748
rect 41043 -21812 41063 -21748
rect 34764 -21828 41063 -21812
rect 34764 -21892 40979 -21828
rect 41043 -21892 41063 -21828
rect 34764 -21908 41063 -21892
rect 34764 -21972 40979 -21908
rect 41043 -21972 41063 -21908
rect 34764 -22000 41063 -21972
rect 41083 -15828 47382 -15800
rect 41083 -15892 47298 -15828
rect 47362 -15892 47382 -15828
rect 41083 -15908 47382 -15892
rect 41083 -15972 47298 -15908
rect 47362 -15972 47382 -15908
rect 41083 -15988 47382 -15972
rect 41083 -16052 47298 -15988
rect 47362 -16052 47382 -15988
rect 41083 -16068 47382 -16052
rect 41083 -16132 47298 -16068
rect 47362 -16132 47382 -16068
rect 41083 -16148 47382 -16132
rect 41083 -16212 47298 -16148
rect 47362 -16212 47382 -16148
rect 41083 -16228 47382 -16212
rect 41083 -16292 47298 -16228
rect 47362 -16292 47382 -16228
rect 41083 -16308 47382 -16292
rect 41083 -16372 47298 -16308
rect 47362 -16372 47382 -16308
rect 41083 -16388 47382 -16372
rect 41083 -16452 47298 -16388
rect 47362 -16452 47382 -16388
rect 41083 -16468 47382 -16452
rect 41083 -16532 47298 -16468
rect 47362 -16532 47382 -16468
rect 41083 -16548 47382 -16532
rect 41083 -16612 47298 -16548
rect 47362 -16612 47382 -16548
rect 41083 -16628 47382 -16612
rect 41083 -16692 47298 -16628
rect 47362 -16692 47382 -16628
rect 41083 -16708 47382 -16692
rect 41083 -16772 47298 -16708
rect 47362 -16772 47382 -16708
rect 41083 -16788 47382 -16772
rect 41083 -16852 47298 -16788
rect 47362 -16852 47382 -16788
rect 41083 -16868 47382 -16852
rect 41083 -16932 47298 -16868
rect 47362 -16932 47382 -16868
rect 41083 -16948 47382 -16932
rect 41083 -17012 47298 -16948
rect 47362 -17012 47382 -16948
rect 41083 -17028 47382 -17012
rect 41083 -17092 47298 -17028
rect 47362 -17092 47382 -17028
rect 41083 -17108 47382 -17092
rect 41083 -17172 47298 -17108
rect 47362 -17172 47382 -17108
rect 41083 -17188 47382 -17172
rect 41083 -17252 47298 -17188
rect 47362 -17252 47382 -17188
rect 41083 -17268 47382 -17252
rect 41083 -17332 47298 -17268
rect 47362 -17332 47382 -17268
rect 41083 -17348 47382 -17332
rect 41083 -17412 47298 -17348
rect 47362 -17412 47382 -17348
rect 41083 -17428 47382 -17412
rect 41083 -17492 47298 -17428
rect 47362 -17492 47382 -17428
rect 41083 -17508 47382 -17492
rect 41083 -17572 47298 -17508
rect 47362 -17572 47382 -17508
rect 41083 -17588 47382 -17572
rect 41083 -17652 47298 -17588
rect 47362 -17652 47382 -17588
rect 41083 -17668 47382 -17652
rect 41083 -17732 47298 -17668
rect 47362 -17732 47382 -17668
rect 41083 -17748 47382 -17732
rect 41083 -17812 47298 -17748
rect 47362 -17812 47382 -17748
rect 41083 -17828 47382 -17812
rect 41083 -17892 47298 -17828
rect 47362 -17892 47382 -17828
rect 41083 -17908 47382 -17892
rect 41083 -17972 47298 -17908
rect 47362 -17972 47382 -17908
rect 41083 -17988 47382 -17972
rect 41083 -18052 47298 -17988
rect 47362 -18052 47382 -17988
rect 41083 -18068 47382 -18052
rect 41083 -18132 47298 -18068
rect 47362 -18132 47382 -18068
rect 41083 -18148 47382 -18132
rect 41083 -18212 47298 -18148
rect 47362 -18212 47382 -18148
rect 41083 -18228 47382 -18212
rect 41083 -18292 47298 -18228
rect 47362 -18292 47382 -18228
rect 41083 -18308 47382 -18292
rect 41083 -18372 47298 -18308
rect 47362 -18372 47382 -18308
rect 41083 -18388 47382 -18372
rect 41083 -18452 47298 -18388
rect 47362 -18452 47382 -18388
rect 41083 -18468 47382 -18452
rect 41083 -18532 47298 -18468
rect 47362 -18532 47382 -18468
rect 41083 -18548 47382 -18532
rect 41083 -18612 47298 -18548
rect 47362 -18612 47382 -18548
rect 41083 -18628 47382 -18612
rect 41083 -18692 47298 -18628
rect 47362 -18692 47382 -18628
rect 41083 -18708 47382 -18692
rect 41083 -18772 47298 -18708
rect 47362 -18772 47382 -18708
rect 41083 -18788 47382 -18772
rect 41083 -18852 47298 -18788
rect 47362 -18852 47382 -18788
rect 41083 -18868 47382 -18852
rect 41083 -18932 47298 -18868
rect 47362 -18932 47382 -18868
rect 41083 -18948 47382 -18932
rect 41083 -19012 47298 -18948
rect 47362 -19012 47382 -18948
rect 41083 -19028 47382 -19012
rect 41083 -19092 47298 -19028
rect 47362 -19092 47382 -19028
rect 41083 -19108 47382 -19092
rect 41083 -19172 47298 -19108
rect 47362 -19172 47382 -19108
rect 41083 -19188 47382 -19172
rect 41083 -19252 47298 -19188
rect 47362 -19252 47382 -19188
rect 41083 -19268 47382 -19252
rect 41083 -19332 47298 -19268
rect 47362 -19332 47382 -19268
rect 41083 -19348 47382 -19332
rect 41083 -19412 47298 -19348
rect 47362 -19412 47382 -19348
rect 41083 -19428 47382 -19412
rect 41083 -19492 47298 -19428
rect 47362 -19492 47382 -19428
rect 41083 -19508 47382 -19492
rect 41083 -19572 47298 -19508
rect 47362 -19572 47382 -19508
rect 41083 -19588 47382 -19572
rect 41083 -19652 47298 -19588
rect 47362 -19652 47382 -19588
rect 41083 -19668 47382 -19652
rect 41083 -19732 47298 -19668
rect 47362 -19732 47382 -19668
rect 41083 -19748 47382 -19732
rect 41083 -19812 47298 -19748
rect 47362 -19812 47382 -19748
rect 41083 -19828 47382 -19812
rect 41083 -19892 47298 -19828
rect 47362 -19892 47382 -19828
rect 41083 -19908 47382 -19892
rect 41083 -19972 47298 -19908
rect 47362 -19972 47382 -19908
rect 41083 -19988 47382 -19972
rect 41083 -20052 47298 -19988
rect 47362 -20052 47382 -19988
rect 41083 -20068 47382 -20052
rect 41083 -20132 47298 -20068
rect 47362 -20132 47382 -20068
rect 41083 -20148 47382 -20132
rect 41083 -20212 47298 -20148
rect 47362 -20212 47382 -20148
rect 41083 -20228 47382 -20212
rect 41083 -20292 47298 -20228
rect 47362 -20292 47382 -20228
rect 41083 -20308 47382 -20292
rect 41083 -20372 47298 -20308
rect 47362 -20372 47382 -20308
rect 41083 -20388 47382 -20372
rect 41083 -20452 47298 -20388
rect 47362 -20452 47382 -20388
rect 41083 -20468 47382 -20452
rect 41083 -20532 47298 -20468
rect 47362 -20532 47382 -20468
rect 41083 -20548 47382 -20532
rect 41083 -20612 47298 -20548
rect 47362 -20612 47382 -20548
rect 41083 -20628 47382 -20612
rect 41083 -20692 47298 -20628
rect 47362 -20692 47382 -20628
rect 41083 -20708 47382 -20692
rect 41083 -20772 47298 -20708
rect 47362 -20772 47382 -20708
rect 41083 -20788 47382 -20772
rect 41083 -20852 47298 -20788
rect 47362 -20852 47382 -20788
rect 41083 -20868 47382 -20852
rect 41083 -20932 47298 -20868
rect 47362 -20932 47382 -20868
rect 41083 -20948 47382 -20932
rect 41083 -21012 47298 -20948
rect 47362 -21012 47382 -20948
rect 41083 -21028 47382 -21012
rect 41083 -21092 47298 -21028
rect 47362 -21092 47382 -21028
rect 41083 -21108 47382 -21092
rect 41083 -21172 47298 -21108
rect 47362 -21172 47382 -21108
rect 41083 -21188 47382 -21172
rect 41083 -21252 47298 -21188
rect 47362 -21252 47382 -21188
rect 41083 -21268 47382 -21252
rect 41083 -21332 47298 -21268
rect 47362 -21332 47382 -21268
rect 41083 -21348 47382 -21332
rect 41083 -21412 47298 -21348
rect 47362 -21412 47382 -21348
rect 41083 -21428 47382 -21412
rect 41083 -21492 47298 -21428
rect 47362 -21492 47382 -21428
rect 41083 -21508 47382 -21492
rect 41083 -21572 47298 -21508
rect 47362 -21572 47382 -21508
rect 41083 -21588 47382 -21572
rect 41083 -21652 47298 -21588
rect 47362 -21652 47382 -21588
rect 41083 -21668 47382 -21652
rect 41083 -21732 47298 -21668
rect 47362 -21732 47382 -21668
rect 41083 -21748 47382 -21732
rect 41083 -21812 47298 -21748
rect 47362 -21812 47382 -21748
rect 41083 -21828 47382 -21812
rect 41083 -21892 47298 -21828
rect 47362 -21892 47382 -21828
rect 41083 -21908 47382 -21892
rect 41083 -21972 47298 -21908
rect 47362 -21972 47382 -21908
rect 41083 -22000 47382 -21972
rect -47383 -22128 -41084 -22100
rect -47383 -22192 -41168 -22128
rect -41104 -22192 -41084 -22128
rect -47383 -22208 -41084 -22192
rect -47383 -22272 -41168 -22208
rect -41104 -22272 -41084 -22208
rect -47383 -22288 -41084 -22272
rect -47383 -22352 -41168 -22288
rect -41104 -22352 -41084 -22288
rect -47383 -22368 -41084 -22352
rect -47383 -22432 -41168 -22368
rect -41104 -22432 -41084 -22368
rect -47383 -22448 -41084 -22432
rect -47383 -22512 -41168 -22448
rect -41104 -22512 -41084 -22448
rect -47383 -22528 -41084 -22512
rect -47383 -22592 -41168 -22528
rect -41104 -22592 -41084 -22528
rect -47383 -22608 -41084 -22592
rect -47383 -22672 -41168 -22608
rect -41104 -22672 -41084 -22608
rect -47383 -22688 -41084 -22672
rect -47383 -22752 -41168 -22688
rect -41104 -22752 -41084 -22688
rect -47383 -22768 -41084 -22752
rect -47383 -22832 -41168 -22768
rect -41104 -22832 -41084 -22768
rect -47383 -22848 -41084 -22832
rect -47383 -22912 -41168 -22848
rect -41104 -22912 -41084 -22848
rect -47383 -22928 -41084 -22912
rect -47383 -22992 -41168 -22928
rect -41104 -22992 -41084 -22928
rect -47383 -23008 -41084 -22992
rect -47383 -23072 -41168 -23008
rect -41104 -23072 -41084 -23008
rect -47383 -23088 -41084 -23072
rect -47383 -23152 -41168 -23088
rect -41104 -23152 -41084 -23088
rect -47383 -23168 -41084 -23152
rect -47383 -23232 -41168 -23168
rect -41104 -23232 -41084 -23168
rect -47383 -23248 -41084 -23232
rect -47383 -23312 -41168 -23248
rect -41104 -23312 -41084 -23248
rect -47383 -23328 -41084 -23312
rect -47383 -23392 -41168 -23328
rect -41104 -23392 -41084 -23328
rect -47383 -23408 -41084 -23392
rect -47383 -23472 -41168 -23408
rect -41104 -23472 -41084 -23408
rect -47383 -23488 -41084 -23472
rect -47383 -23552 -41168 -23488
rect -41104 -23552 -41084 -23488
rect -47383 -23568 -41084 -23552
rect -47383 -23632 -41168 -23568
rect -41104 -23632 -41084 -23568
rect -47383 -23648 -41084 -23632
rect -47383 -23712 -41168 -23648
rect -41104 -23712 -41084 -23648
rect -47383 -23728 -41084 -23712
rect -47383 -23792 -41168 -23728
rect -41104 -23792 -41084 -23728
rect -47383 -23808 -41084 -23792
rect -47383 -23872 -41168 -23808
rect -41104 -23872 -41084 -23808
rect -47383 -23888 -41084 -23872
rect -47383 -23952 -41168 -23888
rect -41104 -23952 -41084 -23888
rect -47383 -23968 -41084 -23952
rect -47383 -24032 -41168 -23968
rect -41104 -24032 -41084 -23968
rect -47383 -24048 -41084 -24032
rect -47383 -24112 -41168 -24048
rect -41104 -24112 -41084 -24048
rect -47383 -24128 -41084 -24112
rect -47383 -24192 -41168 -24128
rect -41104 -24192 -41084 -24128
rect -47383 -24208 -41084 -24192
rect -47383 -24272 -41168 -24208
rect -41104 -24272 -41084 -24208
rect -47383 -24288 -41084 -24272
rect -47383 -24352 -41168 -24288
rect -41104 -24352 -41084 -24288
rect -47383 -24368 -41084 -24352
rect -47383 -24432 -41168 -24368
rect -41104 -24432 -41084 -24368
rect -47383 -24448 -41084 -24432
rect -47383 -24512 -41168 -24448
rect -41104 -24512 -41084 -24448
rect -47383 -24528 -41084 -24512
rect -47383 -24592 -41168 -24528
rect -41104 -24592 -41084 -24528
rect -47383 -24608 -41084 -24592
rect -47383 -24672 -41168 -24608
rect -41104 -24672 -41084 -24608
rect -47383 -24688 -41084 -24672
rect -47383 -24752 -41168 -24688
rect -41104 -24752 -41084 -24688
rect -47383 -24768 -41084 -24752
rect -47383 -24832 -41168 -24768
rect -41104 -24832 -41084 -24768
rect -47383 -24848 -41084 -24832
rect -47383 -24912 -41168 -24848
rect -41104 -24912 -41084 -24848
rect -47383 -24928 -41084 -24912
rect -47383 -24992 -41168 -24928
rect -41104 -24992 -41084 -24928
rect -47383 -25008 -41084 -24992
rect -47383 -25072 -41168 -25008
rect -41104 -25072 -41084 -25008
rect -47383 -25088 -41084 -25072
rect -47383 -25152 -41168 -25088
rect -41104 -25152 -41084 -25088
rect -47383 -25168 -41084 -25152
rect -47383 -25232 -41168 -25168
rect -41104 -25232 -41084 -25168
rect -47383 -25248 -41084 -25232
rect -47383 -25312 -41168 -25248
rect -41104 -25312 -41084 -25248
rect -47383 -25328 -41084 -25312
rect -47383 -25392 -41168 -25328
rect -41104 -25392 -41084 -25328
rect -47383 -25408 -41084 -25392
rect -47383 -25472 -41168 -25408
rect -41104 -25472 -41084 -25408
rect -47383 -25488 -41084 -25472
rect -47383 -25552 -41168 -25488
rect -41104 -25552 -41084 -25488
rect -47383 -25568 -41084 -25552
rect -47383 -25632 -41168 -25568
rect -41104 -25632 -41084 -25568
rect -47383 -25648 -41084 -25632
rect -47383 -25712 -41168 -25648
rect -41104 -25712 -41084 -25648
rect -47383 -25728 -41084 -25712
rect -47383 -25792 -41168 -25728
rect -41104 -25792 -41084 -25728
rect -47383 -25808 -41084 -25792
rect -47383 -25872 -41168 -25808
rect -41104 -25872 -41084 -25808
rect -47383 -25888 -41084 -25872
rect -47383 -25952 -41168 -25888
rect -41104 -25952 -41084 -25888
rect -47383 -25968 -41084 -25952
rect -47383 -26032 -41168 -25968
rect -41104 -26032 -41084 -25968
rect -47383 -26048 -41084 -26032
rect -47383 -26112 -41168 -26048
rect -41104 -26112 -41084 -26048
rect -47383 -26128 -41084 -26112
rect -47383 -26192 -41168 -26128
rect -41104 -26192 -41084 -26128
rect -47383 -26208 -41084 -26192
rect -47383 -26272 -41168 -26208
rect -41104 -26272 -41084 -26208
rect -47383 -26288 -41084 -26272
rect -47383 -26352 -41168 -26288
rect -41104 -26352 -41084 -26288
rect -47383 -26368 -41084 -26352
rect -47383 -26432 -41168 -26368
rect -41104 -26432 -41084 -26368
rect -47383 -26448 -41084 -26432
rect -47383 -26512 -41168 -26448
rect -41104 -26512 -41084 -26448
rect -47383 -26528 -41084 -26512
rect -47383 -26592 -41168 -26528
rect -41104 -26592 -41084 -26528
rect -47383 -26608 -41084 -26592
rect -47383 -26672 -41168 -26608
rect -41104 -26672 -41084 -26608
rect -47383 -26688 -41084 -26672
rect -47383 -26752 -41168 -26688
rect -41104 -26752 -41084 -26688
rect -47383 -26768 -41084 -26752
rect -47383 -26832 -41168 -26768
rect -41104 -26832 -41084 -26768
rect -47383 -26848 -41084 -26832
rect -47383 -26912 -41168 -26848
rect -41104 -26912 -41084 -26848
rect -47383 -26928 -41084 -26912
rect -47383 -26992 -41168 -26928
rect -41104 -26992 -41084 -26928
rect -47383 -27008 -41084 -26992
rect -47383 -27072 -41168 -27008
rect -41104 -27072 -41084 -27008
rect -47383 -27088 -41084 -27072
rect -47383 -27152 -41168 -27088
rect -41104 -27152 -41084 -27088
rect -47383 -27168 -41084 -27152
rect -47383 -27232 -41168 -27168
rect -41104 -27232 -41084 -27168
rect -47383 -27248 -41084 -27232
rect -47383 -27312 -41168 -27248
rect -41104 -27312 -41084 -27248
rect -47383 -27328 -41084 -27312
rect -47383 -27392 -41168 -27328
rect -41104 -27392 -41084 -27328
rect -47383 -27408 -41084 -27392
rect -47383 -27472 -41168 -27408
rect -41104 -27472 -41084 -27408
rect -47383 -27488 -41084 -27472
rect -47383 -27552 -41168 -27488
rect -41104 -27552 -41084 -27488
rect -47383 -27568 -41084 -27552
rect -47383 -27632 -41168 -27568
rect -41104 -27632 -41084 -27568
rect -47383 -27648 -41084 -27632
rect -47383 -27712 -41168 -27648
rect -41104 -27712 -41084 -27648
rect -47383 -27728 -41084 -27712
rect -47383 -27792 -41168 -27728
rect -41104 -27792 -41084 -27728
rect -47383 -27808 -41084 -27792
rect -47383 -27872 -41168 -27808
rect -41104 -27872 -41084 -27808
rect -47383 -27888 -41084 -27872
rect -47383 -27952 -41168 -27888
rect -41104 -27952 -41084 -27888
rect -47383 -27968 -41084 -27952
rect -47383 -28032 -41168 -27968
rect -41104 -28032 -41084 -27968
rect -47383 -28048 -41084 -28032
rect -47383 -28112 -41168 -28048
rect -41104 -28112 -41084 -28048
rect -47383 -28128 -41084 -28112
rect -47383 -28192 -41168 -28128
rect -41104 -28192 -41084 -28128
rect -47383 -28208 -41084 -28192
rect -47383 -28272 -41168 -28208
rect -41104 -28272 -41084 -28208
rect -47383 -28300 -41084 -28272
rect -41064 -22128 -34765 -22100
rect -41064 -22192 -34849 -22128
rect -34785 -22192 -34765 -22128
rect -41064 -22208 -34765 -22192
rect -41064 -22272 -34849 -22208
rect -34785 -22272 -34765 -22208
rect -41064 -22288 -34765 -22272
rect -41064 -22352 -34849 -22288
rect -34785 -22352 -34765 -22288
rect -41064 -22368 -34765 -22352
rect -41064 -22432 -34849 -22368
rect -34785 -22432 -34765 -22368
rect -41064 -22448 -34765 -22432
rect -41064 -22512 -34849 -22448
rect -34785 -22512 -34765 -22448
rect -41064 -22528 -34765 -22512
rect -41064 -22592 -34849 -22528
rect -34785 -22592 -34765 -22528
rect -41064 -22608 -34765 -22592
rect -41064 -22672 -34849 -22608
rect -34785 -22672 -34765 -22608
rect -41064 -22688 -34765 -22672
rect -41064 -22752 -34849 -22688
rect -34785 -22752 -34765 -22688
rect -41064 -22768 -34765 -22752
rect -41064 -22832 -34849 -22768
rect -34785 -22832 -34765 -22768
rect -41064 -22848 -34765 -22832
rect -41064 -22912 -34849 -22848
rect -34785 -22912 -34765 -22848
rect -41064 -22928 -34765 -22912
rect -41064 -22992 -34849 -22928
rect -34785 -22992 -34765 -22928
rect -41064 -23008 -34765 -22992
rect -41064 -23072 -34849 -23008
rect -34785 -23072 -34765 -23008
rect -41064 -23088 -34765 -23072
rect -41064 -23152 -34849 -23088
rect -34785 -23152 -34765 -23088
rect -41064 -23168 -34765 -23152
rect -41064 -23232 -34849 -23168
rect -34785 -23232 -34765 -23168
rect -41064 -23248 -34765 -23232
rect -41064 -23312 -34849 -23248
rect -34785 -23312 -34765 -23248
rect -41064 -23328 -34765 -23312
rect -41064 -23392 -34849 -23328
rect -34785 -23392 -34765 -23328
rect -41064 -23408 -34765 -23392
rect -41064 -23472 -34849 -23408
rect -34785 -23472 -34765 -23408
rect -41064 -23488 -34765 -23472
rect -41064 -23552 -34849 -23488
rect -34785 -23552 -34765 -23488
rect -41064 -23568 -34765 -23552
rect -41064 -23632 -34849 -23568
rect -34785 -23632 -34765 -23568
rect -41064 -23648 -34765 -23632
rect -41064 -23712 -34849 -23648
rect -34785 -23712 -34765 -23648
rect -41064 -23728 -34765 -23712
rect -41064 -23792 -34849 -23728
rect -34785 -23792 -34765 -23728
rect -41064 -23808 -34765 -23792
rect -41064 -23872 -34849 -23808
rect -34785 -23872 -34765 -23808
rect -41064 -23888 -34765 -23872
rect -41064 -23952 -34849 -23888
rect -34785 -23952 -34765 -23888
rect -41064 -23968 -34765 -23952
rect -41064 -24032 -34849 -23968
rect -34785 -24032 -34765 -23968
rect -41064 -24048 -34765 -24032
rect -41064 -24112 -34849 -24048
rect -34785 -24112 -34765 -24048
rect -41064 -24128 -34765 -24112
rect -41064 -24192 -34849 -24128
rect -34785 -24192 -34765 -24128
rect -41064 -24208 -34765 -24192
rect -41064 -24272 -34849 -24208
rect -34785 -24272 -34765 -24208
rect -41064 -24288 -34765 -24272
rect -41064 -24352 -34849 -24288
rect -34785 -24352 -34765 -24288
rect -41064 -24368 -34765 -24352
rect -41064 -24432 -34849 -24368
rect -34785 -24432 -34765 -24368
rect -41064 -24448 -34765 -24432
rect -41064 -24512 -34849 -24448
rect -34785 -24512 -34765 -24448
rect -41064 -24528 -34765 -24512
rect -41064 -24592 -34849 -24528
rect -34785 -24592 -34765 -24528
rect -41064 -24608 -34765 -24592
rect -41064 -24672 -34849 -24608
rect -34785 -24672 -34765 -24608
rect -41064 -24688 -34765 -24672
rect -41064 -24752 -34849 -24688
rect -34785 -24752 -34765 -24688
rect -41064 -24768 -34765 -24752
rect -41064 -24832 -34849 -24768
rect -34785 -24832 -34765 -24768
rect -41064 -24848 -34765 -24832
rect -41064 -24912 -34849 -24848
rect -34785 -24912 -34765 -24848
rect -41064 -24928 -34765 -24912
rect -41064 -24992 -34849 -24928
rect -34785 -24992 -34765 -24928
rect -41064 -25008 -34765 -24992
rect -41064 -25072 -34849 -25008
rect -34785 -25072 -34765 -25008
rect -41064 -25088 -34765 -25072
rect -41064 -25152 -34849 -25088
rect -34785 -25152 -34765 -25088
rect -41064 -25168 -34765 -25152
rect -41064 -25232 -34849 -25168
rect -34785 -25232 -34765 -25168
rect -41064 -25248 -34765 -25232
rect -41064 -25312 -34849 -25248
rect -34785 -25312 -34765 -25248
rect -41064 -25328 -34765 -25312
rect -41064 -25392 -34849 -25328
rect -34785 -25392 -34765 -25328
rect -41064 -25408 -34765 -25392
rect -41064 -25472 -34849 -25408
rect -34785 -25472 -34765 -25408
rect -41064 -25488 -34765 -25472
rect -41064 -25552 -34849 -25488
rect -34785 -25552 -34765 -25488
rect -41064 -25568 -34765 -25552
rect -41064 -25632 -34849 -25568
rect -34785 -25632 -34765 -25568
rect -41064 -25648 -34765 -25632
rect -41064 -25712 -34849 -25648
rect -34785 -25712 -34765 -25648
rect -41064 -25728 -34765 -25712
rect -41064 -25792 -34849 -25728
rect -34785 -25792 -34765 -25728
rect -41064 -25808 -34765 -25792
rect -41064 -25872 -34849 -25808
rect -34785 -25872 -34765 -25808
rect -41064 -25888 -34765 -25872
rect -41064 -25952 -34849 -25888
rect -34785 -25952 -34765 -25888
rect -41064 -25968 -34765 -25952
rect -41064 -26032 -34849 -25968
rect -34785 -26032 -34765 -25968
rect -41064 -26048 -34765 -26032
rect -41064 -26112 -34849 -26048
rect -34785 -26112 -34765 -26048
rect -41064 -26128 -34765 -26112
rect -41064 -26192 -34849 -26128
rect -34785 -26192 -34765 -26128
rect -41064 -26208 -34765 -26192
rect -41064 -26272 -34849 -26208
rect -34785 -26272 -34765 -26208
rect -41064 -26288 -34765 -26272
rect -41064 -26352 -34849 -26288
rect -34785 -26352 -34765 -26288
rect -41064 -26368 -34765 -26352
rect -41064 -26432 -34849 -26368
rect -34785 -26432 -34765 -26368
rect -41064 -26448 -34765 -26432
rect -41064 -26512 -34849 -26448
rect -34785 -26512 -34765 -26448
rect -41064 -26528 -34765 -26512
rect -41064 -26592 -34849 -26528
rect -34785 -26592 -34765 -26528
rect -41064 -26608 -34765 -26592
rect -41064 -26672 -34849 -26608
rect -34785 -26672 -34765 -26608
rect -41064 -26688 -34765 -26672
rect -41064 -26752 -34849 -26688
rect -34785 -26752 -34765 -26688
rect -41064 -26768 -34765 -26752
rect -41064 -26832 -34849 -26768
rect -34785 -26832 -34765 -26768
rect -41064 -26848 -34765 -26832
rect -41064 -26912 -34849 -26848
rect -34785 -26912 -34765 -26848
rect -41064 -26928 -34765 -26912
rect -41064 -26992 -34849 -26928
rect -34785 -26992 -34765 -26928
rect -41064 -27008 -34765 -26992
rect -41064 -27072 -34849 -27008
rect -34785 -27072 -34765 -27008
rect -41064 -27088 -34765 -27072
rect -41064 -27152 -34849 -27088
rect -34785 -27152 -34765 -27088
rect -41064 -27168 -34765 -27152
rect -41064 -27232 -34849 -27168
rect -34785 -27232 -34765 -27168
rect -41064 -27248 -34765 -27232
rect -41064 -27312 -34849 -27248
rect -34785 -27312 -34765 -27248
rect -41064 -27328 -34765 -27312
rect -41064 -27392 -34849 -27328
rect -34785 -27392 -34765 -27328
rect -41064 -27408 -34765 -27392
rect -41064 -27472 -34849 -27408
rect -34785 -27472 -34765 -27408
rect -41064 -27488 -34765 -27472
rect -41064 -27552 -34849 -27488
rect -34785 -27552 -34765 -27488
rect -41064 -27568 -34765 -27552
rect -41064 -27632 -34849 -27568
rect -34785 -27632 -34765 -27568
rect -41064 -27648 -34765 -27632
rect -41064 -27712 -34849 -27648
rect -34785 -27712 -34765 -27648
rect -41064 -27728 -34765 -27712
rect -41064 -27792 -34849 -27728
rect -34785 -27792 -34765 -27728
rect -41064 -27808 -34765 -27792
rect -41064 -27872 -34849 -27808
rect -34785 -27872 -34765 -27808
rect -41064 -27888 -34765 -27872
rect -41064 -27952 -34849 -27888
rect -34785 -27952 -34765 -27888
rect -41064 -27968 -34765 -27952
rect -41064 -28032 -34849 -27968
rect -34785 -28032 -34765 -27968
rect -41064 -28048 -34765 -28032
rect -41064 -28112 -34849 -28048
rect -34785 -28112 -34765 -28048
rect -41064 -28128 -34765 -28112
rect -41064 -28192 -34849 -28128
rect -34785 -28192 -34765 -28128
rect -41064 -28208 -34765 -28192
rect -41064 -28272 -34849 -28208
rect -34785 -28272 -34765 -28208
rect -41064 -28300 -34765 -28272
rect -34745 -22128 -28446 -22100
rect -34745 -22192 -28530 -22128
rect -28466 -22192 -28446 -22128
rect -34745 -22208 -28446 -22192
rect -34745 -22272 -28530 -22208
rect -28466 -22272 -28446 -22208
rect -34745 -22288 -28446 -22272
rect -34745 -22352 -28530 -22288
rect -28466 -22352 -28446 -22288
rect -34745 -22368 -28446 -22352
rect -34745 -22432 -28530 -22368
rect -28466 -22432 -28446 -22368
rect -34745 -22448 -28446 -22432
rect -34745 -22512 -28530 -22448
rect -28466 -22512 -28446 -22448
rect -34745 -22528 -28446 -22512
rect -34745 -22592 -28530 -22528
rect -28466 -22592 -28446 -22528
rect -34745 -22608 -28446 -22592
rect -34745 -22672 -28530 -22608
rect -28466 -22672 -28446 -22608
rect -34745 -22688 -28446 -22672
rect -34745 -22752 -28530 -22688
rect -28466 -22752 -28446 -22688
rect -34745 -22768 -28446 -22752
rect -34745 -22832 -28530 -22768
rect -28466 -22832 -28446 -22768
rect -34745 -22848 -28446 -22832
rect -34745 -22912 -28530 -22848
rect -28466 -22912 -28446 -22848
rect -34745 -22928 -28446 -22912
rect -34745 -22992 -28530 -22928
rect -28466 -22992 -28446 -22928
rect -34745 -23008 -28446 -22992
rect -34745 -23072 -28530 -23008
rect -28466 -23072 -28446 -23008
rect -34745 -23088 -28446 -23072
rect -34745 -23152 -28530 -23088
rect -28466 -23152 -28446 -23088
rect -34745 -23168 -28446 -23152
rect -34745 -23232 -28530 -23168
rect -28466 -23232 -28446 -23168
rect -34745 -23248 -28446 -23232
rect -34745 -23312 -28530 -23248
rect -28466 -23312 -28446 -23248
rect -34745 -23328 -28446 -23312
rect -34745 -23392 -28530 -23328
rect -28466 -23392 -28446 -23328
rect -34745 -23408 -28446 -23392
rect -34745 -23472 -28530 -23408
rect -28466 -23472 -28446 -23408
rect -34745 -23488 -28446 -23472
rect -34745 -23552 -28530 -23488
rect -28466 -23552 -28446 -23488
rect -34745 -23568 -28446 -23552
rect -34745 -23632 -28530 -23568
rect -28466 -23632 -28446 -23568
rect -34745 -23648 -28446 -23632
rect -34745 -23712 -28530 -23648
rect -28466 -23712 -28446 -23648
rect -34745 -23728 -28446 -23712
rect -34745 -23792 -28530 -23728
rect -28466 -23792 -28446 -23728
rect -34745 -23808 -28446 -23792
rect -34745 -23872 -28530 -23808
rect -28466 -23872 -28446 -23808
rect -34745 -23888 -28446 -23872
rect -34745 -23952 -28530 -23888
rect -28466 -23952 -28446 -23888
rect -34745 -23968 -28446 -23952
rect -34745 -24032 -28530 -23968
rect -28466 -24032 -28446 -23968
rect -34745 -24048 -28446 -24032
rect -34745 -24112 -28530 -24048
rect -28466 -24112 -28446 -24048
rect -34745 -24128 -28446 -24112
rect -34745 -24192 -28530 -24128
rect -28466 -24192 -28446 -24128
rect -34745 -24208 -28446 -24192
rect -34745 -24272 -28530 -24208
rect -28466 -24272 -28446 -24208
rect -34745 -24288 -28446 -24272
rect -34745 -24352 -28530 -24288
rect -28466 -24352 -28446 -24288
rect -34745 -24368 -28446 -24352
rect -34745 -24432 -28530 -24368
rect -28466 -24432 -28446 -24368
rect -34745 -24448 -28446 -24432
rect -34745 -24512 -28530 -24448
rect -28466 -24512 -28446 -24448
rect -34745 -24528 -28446 -24512
rect -34745 -24592 -28530 -24528
rect -28466 -24592 -28446 -24528
rect -34745 -24608 -28446 -24592
rect -34745 -24672 -28530 -24608
rect -28466 -24672 -28446 -24608
rect -34745 -24688 -28446 -24672
rect -34745 -24752 -28530 -24688
rect -28466 -24752 -28446 -24688
rect -34745 -24768 -28446 -24752
rect -34745 -24832 -28530 -24768
rect -28466 -24832 -28446 -24768
rect -34745 -24848 -28446 -24832
rect -34745 -24912 -28530 -24848
rect -28466 -24912 -28446 -24848
rect -34745 -24928 -28446 -24912
rect -34745 -24992 -28530 -24928
rect -28466 -24992 -28446 -24928
rect -34745 -25008 -28446 -24992
rect -34745 -25072 -28530 -25008
rect -28466 -25072 -28446 -25008
rect -34745 -25088 -28446 -25072
rect -34745 -25152 -28530 -25088
rect -28466 -25152 -28446 -25088
rect -34745 -25168 -28446 -25152
rect -34745 -25232 -28530 -25168
rect -28466 -25232 -28446 -25168
rect -34745 -25248 -28446 -25232
rect -34745 -25312 -28530 -25248
rect -28466 -25312 -28446 -25248
rect -34745 -25328 -28446 -25312
rect -34745 -25392 -28530 -25328
rect -28466 -25392 -28446 -25328
rect -34745 -25408 -28446 -25392
rect -34745 -25472 -28530 -25408
rect -28466 -25472 -28446 -25408
rect -34745 -25488 -28446 -25472
rect -34745 -25552 -28530 -25488
rect -28466 -25552 -28446 -25488
rect -34745 -25568 -28446 -25552
rect -34745 -25632 -28530 -25568
rect -28466 -25632 -28446 -25568
rect -34745 -25648 -28446 -25632
rect -34745 -25712 -28530 -25648
rect -28466 -25712 -28446 -25648
rect -34745 -25728 -28446 -25712
rect -34745 -25792 -28530 -25728
rect -28466 -25792 -28446 -25728
rect -34745 -25808 -28446 -25792
rect -34745 -25872 -28530 -25808
rect -28466 -25872 -28446 -25808
rect -34745 -25888 -28446 -25872
rect -34745 -25952 -28530 -25888
rect -28466 -25952 -28446 -25888
rect -34745 -25968 -28446 -25952
rect -34745 -26032 -28530 -25968
rect -28466 -26032 -28446 -25968
rect -34745 -26048 -28446 -26032
rect -34745 -26112 -28530 -26048
rect -28466 -26112 -28446 -26048
rect -34745 -26128 -28446 -26112
rect -34745 -26192 -28530 -26128
rect -28466 -26192 -28446 -26128
rect -34745 -26208 -28446 -26192
rect -34745 -26272 -28530 -26208
rect -28466 -26272 -28446 -26208
rect -34745 -26288 -28446 -26272
rect -34745 -26352 -28530 -26288
rect -28466 -26352 -28446 -26288
rect -34745 -26368 -28446 -26352
rect -34745 -26432 -28530 -26368
rect -28466 -26432 -28446 -26368
rect -34745 -26448 -28446 -26432
rect -34745 -26512 -28530 -26448
rect -28466 -26512 -28446 -26448
rect -34745 -26528 -28446 -26512
rect -34745 -26592 -28530 -26528
rect -28466 -26592 -28446 -26528
rect -34745 -26608 -28446 -26592
rect -34745 -26672 -28530 -26608
rect -28466 -26672 -28446 -26608
rect -34745 -26688 -28446 -26672
rect -34745 -26752 -28530 -26688
rect -28466 -26752 -28446 -26688
rect -34745 -26768 -28446 -26752
rect -34745 -26832 -28530 -26768
rect -28466 -26832 -28446 -26768
rect -34745 -26848 -28446 -26832
rect -34745 -26912 -28530 -26848
rect -28466 -26912 -28446 -26848
rect -34745 -26928 -28446 -26912
rect -34745 -26992 -28530 -26928
rect -28466 -26992 -28446 -26928
rect -34745 -27008 -28446 -26992
rect -34745 -27072 -28530 -27008
rect -28466 -27072 -28446 -27008
rect -34745 -27088 -28446 -27072
rect -34745 -27152 -28530 -27088
rect -28466 -27152 -28446 -27088
rect -34745 -27168 -28446 -27152
rect -34745 -27232 -28530 -27168
rect -28466 -27232 -28446 -27168
rect -34745 -27248 -28446 -27232
rect -34745 -27312 -28530 -27248
rect -28466 -27312 -28446 -27248
rect -34745 -27328 -28446 -27312
rect -34745 -27392 -28530 -27328
rect -28466 -27392 -28446 -27328
rect -34745 -27408 -28446 -27392
rect -34745 -27472 -28530 -27408
rect -28466 -27472 -28446 -27408
rect -34745 -27488 -28446 -27472
rect -34745 -27552 -28530 -27488
rect -28466 -27552 -28446 -27488
rect -34745 -27568 -28446 -27552
rect -34745 -27632 -28530 -27568
rect -28466 -27632 -28446 -27568
rect -34745 -27648 -28446 -27632
rect -34745 -27712 -28530 -27648
rect -28466 -27712 -28446 -27648
rect -34745 -27728 -28446 -27712
rect -34745 -27792 -28530 -27728
rect -28466 -27792 -28446 -27728
rect -34745 -27808 -28446 -27792
rect -34745 -27872 -28530 -27808
rect -28466 -27872 -28446 -27808
rect -34745 -27888 -28446 -27872
rect -34745 -27952 -28530 -27888
rect -28466 -27952 -28446 -27888
rect -34745 -27968 -28446 -27952
rect -34745 -28032 -28530 -27968
rect -28466 -28032 -28446 -27968
rect -34745 -28048 -28446 -28032
rect -34745 -28112 -28530 -28048
rect -28466 -28112 -28446 -28048
rect -34745 -28128 -28446 -28112
rect -34745 -28192 -28530 -28128
rect -28466 -28192 -28446 -28128
rect -34745 -28208 -28446 -28192
rect -34745 -28272 -28530 -28208
rect -28466 -28272 -28446 -28208
rect -34745 -28300 -28446 -28272
rect -28426 -22128 -22127 -22100
rect -28426 -22192 -22211 -22128
rect -22147 -22192 -22127 -22128
rect -28426 -22208 -22127 -22192
rect -28426 -22272 -22211 -22208
rect -22147 -22272 -22127 -22208
rect -28426 -22288 -22127 -22272
rect -28426 -22352 -22211 -22288
rect -22147 -22352 -22127 -22288
rect -28426 -22368 -22127 -22352
rect -28426 -22432 -22211 -22368
rect -22147 -22432 -22127 -22368
rect -28426 -22448 -22127 -22432
rect -28426 -22512 -22211 -22448
rect -22147 -22512 -22127 -22448
rect -28426 -22528 -22127 -22512
rect -28426 -22592 -22211 -22528
rect -22147 -22592 -22127 -22528
rect -28426 -22608 -22127 -22592
rect -28426 -22672 -22211 -22608
rect -22147 -22672 -22127 -22608
rect -28426 -22688 -22127 -22672
rect -28426 -22752 -22211 -22688
rect -22147 -22752 -22127 -22688
rect -28426 -22768 -22127 -22752
rect -28426 -22832 -22211 -22768
rect -22147 -22832 -22127 -22768
rect -28426 -22848 -22127 -22832
rect -28426 -22912 -22211 -22848
rect -22147 -22912 -22127 -22848
rect -28426 -22928 -22127 -22912
rect -28426 -22992 -22211 -22928
rect -22147 -22992 -22127 -22928
rect -28426 -23008 -22127 -22992
rect -28426 -23072 -22211 -23008
rect -22147 -23072 -22127 -23008
rect -28426 -23088 -22127 -23072
rect -28426 -23152 -22211 -23088
rect -22147 -23152 -22127 -23088
rect -28426 -23168 -22127 -23152
rect -28426 -23232 -22211 -23168
rect -22147 -23232 -22127 -23168
rect -28426 -23248 -22127 -23232
rect -28426 -23312 -22211 -23248
rect -22147 -23312 -22127 -23248
rect -28426 -23328 -22127 -23312
rect -28426 -23392 -22211 -23328
rect -22147 -23392 -22127 -23328
rect -28426 -23408 -22127 -23392
rect -28426 -23472 -22211 -23408
rect -22147 -23472 -22127 -23408
rect -28426 -23488 -22127 -23472
rect -28426 -23552 -22211 -23488
rect -22147 -23552 -22127 -23488
rect -28426 -23568 -22127 -23552
rect -28426 -23632 -22211 -23568
rect -22147 -23632 -22127 -23568
rect -28426 -23648 -22127 -23632
rect -28426 -23712 -22211 -23648
rect -22147 -23712 -22127 -23648
rect -28426 -23728 -22127 -23712
rect -28426 -23792 -22211 -23728
rect -22147 -23792 -22127 -23728
rect -28426 -23808 -22127 -23792
rect -28426 -23872 -22211 -23808
rect -22147 -23872 -22127 -23808
rect -28426 -23888 -22127 -23872
rect -28426 -23952 -22211 -23888
rect -22147 -23952 -22127 -23888
rect -28426 -23968 -22127 -23952
rect -28426 -24032 -22211 -23968
rect -22147 -24032 -22127 -23968
rect -28426 -24048 -22127 -24032
rect -28426 -24112 -22211 -24048
rect -22147 -24112 -22127 -24048
rect -28426 -24128 -22127 -24112
rect -28426 -24192 -22211 -24128
rect -22147 -24192 -22127 -24128
rect -28426 -24208 -22127 -24192
rect -28426 -24272 -22211 -24208
rect -22147 -24272 -22127 -24208
rect -28426 -24288 -22127 -24272
rect -28426 -24352 -22211 -24288
rect -22147 -24352 -22127 -24288
rect -28426 -24368 -22127 -24352
rect -28426 -24432 -22211 -24368
rect -22147 -24432 -22127 -24368
rect -28426 -24448 -22127 -24432
rect -28426 -24512 -22211 -24448
rect -22147 -24512 -22127 -24448
rect -28426 -24528 -22127 -24512
rect -28426 -24592 -22211 -24528
rect -22147 -24592 -22127 -24528
rect -28426 -24608 -22127 -24592
rect -28426 -24672 -22211 -24608
rect -22147 -24672 -22127 -24608
rect -28426 -24688 -22127 -24672
rect -28426 -24752 -22211 -24688
rect -22147 -24752 -22127 -24688
rect -28426 -24768 -22127 -24752
rect -28426 -24832 -22211 -24768
rect -22147 -24832 -22127 -24768
rect -28426 -24848 -22127 -24832
rect -28426 -24912 -22211 -24848
rect -22147 -24912 -22127 -24848
rect -28426 -24928 -22127 -24912
rect -28426 -24992 -22211 -24928
rect -22147 -24992 -22127 -24928
rect -28426 -25008 -22127 -24992
rect -28426 -25072 -22211 -25008
rect -22147 -25072 -22127 -25008
rect -28426 -25088 -22127 -25072
rect -28426 -25152 -22211 -25088
rect -22147 -25152 -22127 -25088
rect -28426 -25168 -22127 -25152
rect -28426 -25232 -22211 -25168
rect -22147 -25232 -22127 -25168
rect -28426 -25248 -22127 -25232
rect -28426 -25312 -22211 -25248
rect -22147 -25312 -22127 -25248
rect -28426 -25328 -22127 -25312
rect -28426 -25392 -22211 -25328
rect -22147 -25392 -22127 -25328
rect -28426 -25408 -22127 -25392
rect -28426 -25472 -22211 -25408
rect -22147 -25472 -22127 -25408
rect -28426 -25488 -22127 -25472
rect -28426 -25552 -22211 -25488
rect -22147 -25552 -22127 -25488
rect -28426 -25568 -22127 -25552
rect -28426 -25632 -22211 -25568
rect -22147 -25632 -22127 -25568
rect -28426 -25648 -22127 -25632
rect -28426 -25712 -22211 -25648
rect -22147 -25712 -22127 -25648
rect -28426 -25728 -22127 -25712
rect -28426 -25792 -22211 -25728
rect -22147 -25792 -22127 -25728
rect -28426 -25808 -22127 -25792
rect -28426 -25872 -22211 -25808
rect -22147 -25872 -22127 -25808
rect -28426 -25888 -22127 -25872
rect -28426 -25952 -22211 -25888
rect -22147 -25952 -22127 -25888
rect -28426 -25968 -22127 -25952
rect -28426 -26032 -22211 -25968
rect -22147 -26032 -22127 -25968
rect -28426 -26048 -22127 -26032
rect -28426 -26112 -22211 -26048
rect -22147 -26112 -22127 -26048
rect -28426 -26128 -22127 -26112
rect -28426 -26192 -22211 -26128
rect -22147 -26192 -22127 -26128
rect -28426 -26208 -22127 -26192
rect -28426 -26272 -22211 -26208
rect -22147 -26272 -22127 -26208
rect -28426 -26288 -22127 -26272
rect -28426 -26352 -22211 -26288
rect -22147 -26352 -22127 -26288
rect -28426 -26368 -22127 -26352
rect -28426 -26432 -22211 -26368
rect -22147 -26432 -22127 -26368
rect -28426 -26448 -22127 -26432
rect -28426 -26512 -22211 -26448
rect -22147 -26512 -22127 -26448
rect -28426 -26528 -22127 -26512
rect -28426 -26592 -22211 -26528
rect -22147 -26592 -22127 -26528
rect -28426 -26608 -22127 -26592
rect -28426 -26672 -22211 -26608
rect -22147 -26672 -22127 -26608
rect -28426 -26688 -22127 -26672
rect -28426 -26752 -22211 -26688
rect -22147 -26752 -22127 -26688
rect -28426 -26768 -22127 -26752
rect -28426 -26832 -22211 -26768
rect -22147 -26832 -22127 -26768
rect -28426 -26848 -22127 -26832
rect -28426 -26912 -22211 -26848
rect -22147 -26912 -22127 -26848
rect -28426 -26928 -22127 -26912
rect -28426 -26992 -22211 -26928
rect -22147 -26992 -22127 -26928
rect -28426 -27008 -22127 -26992
rect -28426 -27072 -22211 -27008
rect -22147 -27072 -22127 -27008
rect -28426 -27088 -22127 -27072
rect -28426 -27152 -22211 -27088
rect -22147 -27152 -22127 -27088
rect -28426 -27168 -22127 -27152
rect -28426 -27232 -22211 -27168
rect -22147 -27232 -22127 -27168
rect -28426 -27248 -22127 -27232
rect -28426 -27312 -22211 -27248
rect -22147 -27312 -22127 -27248
rect -28426 -27328 -22127 -27312
rect -28426 -27392 -22211 -27328
rect -22147 -27392 -22127 -27328
rect -28426 -27408 -22127 -27392
rect -28426 -27472 -22211 -27408
rect -22147 -27472 -22127 -27408
rect -28426 -27488 -22127 -27472
rect -28426 -27552 -22211 -27488
rect -22147 -27552 -22127 -27488
rect -28426 -27568 -22127 -27552
rect -28426 -27632 -22211 -27568
rect -22147 -27632 -22127 -27568
rect -28426 -27648 -22127 -27632
rect -28426 -27712 -22211 -27648
rect -22147 -27712 -22127 -27648
rect -28426 -27728 -22127 -27712
rect -28426 -27792 -22211 -27728
rect -22147 -27792 -22127 -27728
rect -28426 -27808 -22127 -27792
rect -28426 -27872 -22211 -27808
rect -22147 -27872 -22127 -27808
rect -28426 -27888 -22127 -27872
rect -28426 -27952 -22211 -27888
rect -22147 -27952 -22127 -27888
rect -28426 -27968 -22127 -27952
rect -28426 -28032 -22211 -27968
rect -22147 -28032 -22127 -27968
rect -28426 -28048 -22127 -28032
rect -28426 -28112 -22211 -28048
rect -22147 -28112 -22127 -28048
rect -28426 -28128 -22127 -28112
rect -28426 -28192 -22211 -28128
rect -22147 -28192 -22127 -28128
rect -28426 -28208 -22127 -28192
rect -28426 -28272 -22211 -28208
rect -22147 -28272 -22127 -28208
rect -28426 -28300 -22127 -28272
rect -22107 -22128 -15808 -22100
rect -22107 -22192 -15892 -22128
rect -15828 -22192 -15808 -22128
rect -22107 -22208 -15808 -22192
rect -22107 -22272 -15892 -22208
rect -15828 -22272 -15808 -22208
rect -22107 -22288 -15808 -22272
rect -22107 -22352 -15892 -22288
rect -15828 -22352 -15808 -22288
rect -22107 -22368 -15808 -22352
rect -22107 -22432 -15892 -22368
rect -15828 -22432 -15808 -22368
rect -22107 -22448 -15808 -22432
rect -22107 -22512 -15892 -22448
rect -15828 -22512 -15808 -22448
rect -22107 -22528 -15808 -22512
rect -22107 -22592 -15892 -22528
rect -15828 -22592 -15808 -22528
rect -22107 -22608 -15808 -22592
rect -22107 -22672 -15892 -22608
rect -15828 -22672 -15808 -22608
rect -22107 -22688 -15808 -22672
rect -22107 -22752 -15892 -22688
rect -15828 -22752 -15808 -22688
rect -22107 -22768 -15808 -22752
rect -22107 -22832 -15892 -22768
rect -15828 -22832 -15808 -22768
rect -22107 -22848 -15808 -22832
rect -22107 -22912 -15892 -22848
rect -15828 -22912 -15808 -22848
rect -22107 -22928 -15808 -22912
rect -22107 -22992 -15892 -22928
rect -15828 -22992 -15808 -22928
rect -22107 -23008 -15808 -22992
rect -22107 -23072 -15892 -23008
rect -15828 -23072 -15808 -23008
rect -22107 -23088 -15808 -23072
rect -22107 -23152 -15892 -23088
rect -15828 -23152 -15808 -23088
rect -22107 -23168 -15808 -23152
rect -22107 -23232 -15892 -23168
rect -15828 -23232 -15808 -23168
rect -22107 -23248 -15808 -23232
rect -22107 -23312 -15892 -23248
rect -15828 -23312 -15808 -23248
rect -22107 -23328 -15808 -23312
rect -22107 -23392 -15892 -23328
rect -15828 -23392 -15808 -23328
rect -22107 -23408 -15808 -23392
rect -22107 -23472 -15892 -23408
rect -15828 -23472 -15808 -23408
rect -22107 -23488 -15808 -23472
rect -22107 -23552 -15892 -23488
rect -15828 -23552 -15808 -23488
rect -22107 -23568 -15808 -23552
rect -22107 -23632 -15892 -23568
rect -15828 -23632 -15808 -23568
rect -22107 -23648 -15808 -23632
rect -22107 -23712 -15892 -23648
rect -15828 -23712 -15808 -23648
rect -22107 -23728 -15808 -23712
rect -22107 -23792 -15892 -23728
rect -15828 -23792 -15808 -23728
rect -22107 -23808 -15808 -23792
rect -22107 -23872 -15892 -23808
rect -15828 -23872 -15808 -23808
rect -22107 -23888 -15808 -23872
rect -22107 -23952 -15892 -23888
rect -15828 -23952 -15808 -23888
rect -22107 -23968 -15808 -23952
rect -22107 -24032 -15892 -23968
rect -15828 -24032 -15808 -23968
rect -22107 -24048 -15808 -24032
rect -22107 -24112 -15892 -24048
rect -15828 -24112 -15808 -24048
rect -22107 -24128 -15808 -24112
rect -22107 -24192 -15892 -24128
rect -15828 -24192 -15808 -24128
rect -22107 -24208 -15808 -24192
rect -22107 -24272 -15892 -24208
rect -15828 -24272 -15808 -24208
rect -22107 -24288 -15808 -24272
rect -22107 -24352 -15892 -24288
rect -15828 -24352 -15808 -24288
rect -22107 -24368 -15808 -24352
rect -22107 -24432 -15892 -24368
rect -15828 -24432 -15808 -24368
rect -22107 -24448 -15808 -24432
rect -22107 -24512 -15892 -24448
rect -15828 -24512 -15808 -24448
rect -22107 -24528 -15808 -24512
rect -22107 -24592 -15892 -24528
rect -15828 -24592 -15808 -24528
rect -22107 -24608 -15808 -24592
rect -22107 -24672 -15892 -24608
rect -15828 -24672 -15808 -24608
rect -22107 -24688 -15808 -24672
rect -22107 -24752 -15892 -24688
rect -15828 -24752 -15808 -24688
rect -22107 -24768 -15808 -24752
rect -22107 -24832 -15892 -24768
rect -15828 -24832 -15808 -24768
rect -22107 -24848 -15808 -24832
rect -22107 -24912 -15892 -24848
rect -15828 -24912 -15808 -24848
rect -22107 -24928 -15808 -24912
rect -22107 -24992 -15892 -24928
rect -15828 -24992 -15808 -24928
rect -22107 -25008 -15808 -24992
rect -22107 -25072 -15892 -25008
rect -15828 -25072 -15808 -25008
rect -22107 -25088 -15808 -25072
rect -22107 -25152 -15892 -25088
rect -15828 -25152 -15808 -25088
rect -22107 -25168 -15808 -25152
rect -22107 -25232 -15892 -25168
rect -15828 -25232 -15808 -25168
rect -22107 -25248 -15808 -25232
rect -22107 -25312 -15892 -25248
rect -15828 -25312 -15808 -25248
rect -22107 -25328 -15808 -25312
rect -22107 -25392 -15892 -25328
rect -15828 -25392 -15808 -25328
rect -22107 -25408 -15808 -25392
rect -22107 -25472 -15892 -25408
rect -15828 -25472 -15808 -25408
rect -22107 -25488 -15808 -25472
rect -22107 -25552 -15892 -25488
rect -15828 -25552 -15808 -25488
rect -22107 -25568 -15808 -25552
rect -22107 -25632 -15892 -25568
rect -15828 -25632 -15808 -25568
rect -22107 -25648 -15808 -25632
rect -22107 -25712 -15892 -25648
rect -15828 -25712 -15808 -25648
rect -22107 -25728 -15808 -25712
rect -22107 -25792 -15892 -25728
rect -15828 -25792 -15808 -25728
rect -22107 -25808 -15808 -25792
rect -22107 -25872 -15892 -25808
rect -15828 -25872 -15808 -25808
rect -22107 -25888 -15808 -25872
rect -22107 -25952 -15892 -25888
rect -15828 -25952 -15808 -25888
rect -22107 -25968 -15808 -25952
rect -22107 -26032 -15892 -25968
rect -15828 -26032 -15808 -25968
rect -22107 -26048 -15808 -26032
rect -22107 -26112 -15892 -26048
rect -15828 -26112 -15808 -26048
rect -22107 -26128 -15808 -26112
rect -22107 -26192 -15892 -26128
rect -15828 -26192 -15808 -26128
rect -22107 -26208 -15808 -26192
rect -22107 -26272 -15892 -26208
rect -15828 -26272 -15808 -26208
rect -22107 -26288 -15808 -26272
rect -22107 -26352 -15892 -26288
rect -15828 -26352 -15808 -26288
rect -22107 -26368 -15808 -26352
rect -22107 -26432 -15892 -26368
rect -15828 -26432 -15808 -26368
rect -22107 -26448 -15808 -26432
rect -22107 -26512 -15892 -26448
rect -15828 -26512 -15808 -26448
rect -22107 -26528 -15808 -26512
rect -22107 -26592 -15892 -26528
rect -15828 -26592 -15808 -26528
rect -22107 -26608 -15808 -26592
rect -22107 -26672 -15892 -26608
rect -15828 -26672 -15808 -26608
rect -22107 -26688 -15808 -26672
rect -22107 -26752 -15892 -26688
rect -15828 -26752 -15808 -26688
rect -22107 -26768 -15808 -26752
rect -22107 -26832 -15892 -26768
rect -15828 -26832 -15808 -26768
rect -22107 -26848 -15808 -26832
rect -22107 -26912 -15892 -26848
rect -15828 -26912 -15808 -26848
rect -22107 -26928 -15808 -26912
rect -22107 -26992 -15892 -26928
rect -15828 -26992 -15808 -26928
rect -22107 -27008 -15808 -26992
rect -22107 -27072 -15892 -27008
rect -15828 -27072 -15808 -27008
rect -22107 -27088 -15808 -27072
rect -22107 -27152 -15892 -27088
rect -15828 -27152 -15808 -27088
rect -22107 -27168 -15808 -27152
rect -22107 -27232 -15892 -27168
rect -15828 -27232 -15808 -27168
rect -22107 -27248 -15808 -27232
rect -22107 -27312 -15892 -27248
rect -15828 -27312 -15808 -27248
rect -22107 -27328 -15808 -27312
rect -22107 -27392 -15892 -27328
rect -15828 -27392 -15808 -27328
rect -22107 -27408 -15808 -27392
rect -22107 -27472 -15892 -27408
rect -15828 -27472 -15808 -27408
rect -22107 -27488 -15808 -27472
rect -22107 -27552 -15892 -27488
rect -15828 -27552 -15808 -27488
rect -22107 -27568 -15808 -27552
rect -22107 -27632 -15892 -27568
rect -15828 -27632 -15808 -27568
rect -22107 -27648 -15808 -27632
rect -22107 -27712 -15892 -27648
rect -15828 -27712 -15808 -27648
rect -22107 -27728 -15808 -27712
rect -22107 -27792 -15892 -27728
rect -15828 -27792 -15808 -27728
rect -22107 -27808 -15808 -27792
rect -22107 -27872 -15892 -27808
rect -15828 -27872 -15808 -27808
rect -22107 -27888 -15808 -27872
rect -22107 -27952 -15892 -27888
rect -15828 -27952 -15808 -27888
rect -22107 -27968 -15808 -27952
rect -22107 -28032 -15892 -27968
rect -15828 -28032 -15808 -27968
rect -22107 -28048 -15808 -28032
rect -22107 -28112 -15892 -28048
rect -15828 -28112 -15808 -28048
rect -22107 -28128 -15808 -28112
rect -22107 -28192 -15892 -28128
rect -15828 -28192 -15808 -28128
rect -22107 -28208 -15808 -28192
rect -22107 -28272 -15892 -28208
rect -15828 -28272 -15808 -28208
rect -22107 -28300 -15808 -28272
rect -15788 -22128 -9489 -22100
rect -15788 -22192 -9573 -22128
rect -9509 -22192 -9489 -22128
rect -15788 -22208 -9489 -22192
rect -15788 -22272 -9573 -22208
rect -9509 -22272 -9489 -22208
rect -15788 -22288 -9489 -22272
rect -15788 -22352 -9573 -22288
rect -9509 -22352 -9489 -22288
rect -15788 -22368 -9489 -22352
rect -15788 -22432 -9573 -22368
rect -9509 -22432 -9489 -22368
rect -15788 -22448 -9489 -22432
rect -15788 -22512 -9573 -22448
rect -9509 -22512 -9489 -22448
rect -15788 -22528 -9489 -22512
rect -15788 -22592 -9573 -22528
rect -9509 -22592 -9489 -22528
rect -15788 -22608 -9489 -22592
rect -15788 -22672 -9573 -22608
rect -9509 -22672 -9489 -22608
rect -15788 -22688 -9489 -22672
rect -15788 -22752 -9573 -22688
rect -9509 -22752 -9489 -22688
rect -15788 -22768 -9489 -22752
rect -15788 -22832 -9573 -22768
rect -9509 -22832 -9489 -22768
rect -15788 -22848 -9489 -22832
rect -15788 -22912 -9573 -22848
rect -9509 -22912 -9489 -22848
rect -15788 -22928 -9489 -22912
rect -15788 -22992 -9573 -22928
rect -9509 -22992 -9489 -22928
rect -15788 -23008 -9489 -22992
rect -15788 -23072 -9573 -23008
rect -9509 -23072 -9489 -23008
rect -15788 -23088 -9489 -23072
rect -15788 -23152 -9573 -23088
rect -9509 -23152 -9489 -23088
rect -15788 -23168 -9489 -23152
rect -15788 -23232 -9573 -23168
rect -9509 -23232 -9489 -23168
rect -15788 -23248 -9489 -23232
rect -15788 -23312 -9573 -23248
rect -9509 -23312 -9489 -23248
rect -15788 -23328 -9489 -23312
rect -15788 -23392 -9573 -23328
rect -9509 -23392 -9489 -23328
rect -15788 -23408 -9489 -23392
rect -15788 -23472 -9573 -23408
rect -9509 -23472 -9489 -23408
rect -15788 -23488 -9489 -23472
rect -15788 -23552 -9573 -23488
rect -9509 -23552 -9489 -23488
rect -15788 -23568 -9489 -23552
rect -15788 -23632 -9573 -23568
rect -9509 -23632 -9489 -23568
rect -15788 -23648 -9489 -23632
rect -15788 -23712 -9573 -23648
rect -9509 -23712 -9489 -23648
rect -15788 -23728 -9489 -23712
rect -15788 -23792 -9573 -23728
rect -9509 -23792 -9489 -23728
rect -15788 -23808 -9489 -23792
rect -15788 -23872 -9573 -23808
rect -9509 -23872 -9489 -23808
rect -15788 -23888 -9489 -23872
rect -15788 -23952 -9573 -23888
rect -9509 -23952 -9489 -23888
rect -15788 -23968 -9489 -23952
rect -15788 -24032 -9573 -23968
rect -9509 -24032 -9489 -23968
rect -15788 -24048 -9489 -24032
rect -15788 -24112 -9573 -24048
rect -9509 -24112 -9489 -24048
rect -15788 -24128 -9489 -24112
rect -15788 -24192 -9573 -24128
rect -9509 -24192 -9489 -24128
rect -15788 -24208 -9489 -24192
rect -15788 -24272 -9573 -24208
rect -9509 -24272 -9489 -24208
rect -15788 -24288 -9489 -24272
rect -15788 -24352 -9573 -24288
rect -9509 -24352 -9489 -24288
rect -15788 -24368 -9489 -24352
rect -15788 -24432 -9573 -24368
rect -9509 -24432 -9489 -24368
rect -15788 -24448 -9489 -24432
rect -15788 -24512 -9573 -24448
rect -9509 -24512 -9489 -24448
rect -15788 -24528 -9489 -24512
rect -15788 -24592 -9573 -24528
rect -9509 -24592 -9489 -24528
rect -15788 -24608 -9489 -24592
rect -15788 -24672 -9573 -24608
rect -9509 -24672 -9489 -24608
rect -15788 -24688 -9489 -24672
rect -15788 -24752 -9573 -24688
rect -9509 -24752 -9489 -24688
rect -15788 -24768 -9489 -24752
rect -15788 -24832 -9573 -24768
rect -9509 -24832 -9489 -24768
rect -15788 -24848 -9489 -24832
rect -15788 -24912 -9573 -24848
rect -9509 -24912 -9489 -24848
rect -15788 -24928 -9489 -24912
rect -15788 -24992 -9573 -24928
rect -9509 -24992 -9489 -24928
rect -15788 -25008 -9489 -24992
rect -15788 -25072 -9573 -25008
rect -9509 -25072 -9489 -25008
rect -15788 -25088 -9489 -25072
rect -15788 -25152 -9573 -25088
rect -9509 -25152 -9489 -25088
rect -15788 -25168 -9489 -25152
rect -15788 -25232 -9573 -25168
rect -9509 -25232 -9489 -25168
rect -15788 -25248 -9489 -25232
rect -15788 -25312 -9573 -25248
rect -9509 -25312 -9489 -25248
rect -15788 -25328 -9489 -25312
rect -15788 -25392 -9573 -25328
rect -9509 -25392 -9489 -25328
rect -15788 -25408 -9489 -25392
rect -15788 -25472 -9573 -25408
rect -9509 -25472 -9489 -25408
rect -15788 -25488 -9489 -25472
rect -15788 -25552 -9573 -25488
rect -9509 -25552 -9489 -25488
rect -15788 -25568 -9489 -25552
rect -15788 -25632 -9573 -25568
rect -9509 -25632 -9489 -25568
rect -15788 -25648 -9489 -25632
rect -15788 -25712 -9573 -25648
rect -9509 -25712 -9489 -25648
rect -15788 -25728 -9489 -25712
rect -15788 -25792 -9573 -25728
rect -9509 -25792 -9489 -25728
rect -15788 -25808 -9489 -25792
rect -15788 -25872 -9573 -25808
rect -9509 -25872 -9489 -25808
rect -15788 -25888 -9489 -25872
rect -15788 -25952 -9573 -25888
rect -9509 -25952 -9489 -25888
rect -15788 -25968 -9489 -25952
rect -15788 -26032 -9573 -25968
rect -9509 -26032 -9489 -25968
rect -15788 -26048 -9489 -26032
rect -15788 -26112 -9573 -26048
rect -9509 -26112 -9489 -26048
rect -15788 -26128 -9489 -26112
rect -15788 -26192 -9573 -26128
rect -9509 -26192 -9489 -26128
rect -15788 -26208 -9489 -26192
rect -15788 -26272 -9573 -26208
rect -9509 -26272 -9489 -26208
rect -15788 -26288 -9489 -26272
rect -15788 -26352 -9573 -26288
rect -9509 -26352 -9489 -26288
rect -15788 -26368 -9489 -26352
rect -15788 -26432 -9573 -26368
rect -9509 -26432 -9489 -26368
rect -15788 -26448 -9489 -26432
rect -15788 -26512 -9573 -26448
rect -9509 -26512 -9489 -26448
rect -15788 -26528 -9489 -26512
rect -15788 -26592 -9573 -26528
rect -9509 -26592 -9489 -26528
rect -15788 -26608 -9489 -26592
rect -15788 -26672 -9573 -26608
rect -9509 -26672 -9489 -26608
rect -15788 -26688 -9489 -26672
rect -15788 -26752 -9573 -26688
rect -9509 -26752 -9489 -26688
rect -15788 -26768 -9489 -26752
rect -15788 -26832 -9573 -26768
rect -9509 -26832 -9489 -26768
rect -15788 -26848 -9489 -26832
rect -15788 -26912 -9573 -26848
rect -9509 -26912 -9489 -26848
rect -15788 -26928 -9489 -26912
rect -15788 -26992 -9573 -26928
rect -9509 -26992 -9489 -26928
rect -15788 -27008 -9489 -26992
rect -15788 -27072 -9573 -27008
rect -9509 -27072 -9489 -27008
rect -15788 -27088 -9489 -27072
rect -15788 -27152 -9573 -27088
rect -9509 -27152 -9489 -27088
rect -15788 -27168 -9489 -27152
rect -15788 -27232 -9573 -27168
rect -9509 -27232 -9489 -27168
rect -15788 -27248 -9489 -27232
rect -15788 -27312 -9573 -27248
rect -9509 -27312 -9489 -27248
rect -15788 -27328 -9489 -27312
rect -15788 -27392 -9573 -27328
rect -9509 -27392 -9489 -27328
rect -15788 -27408 -9489 -27392
rect -15788 -27472 -9573 -27408
rect -9509 -27472 -9489 -27408
rect -15788 -27488 -9489 -27472
rect -15788 -27552 -9573 -27488
rect -9509 -27552 -9489 -27488
rect -15788 -27568 -9489 -27552
rect -15788 -27632 -9573 -27568
rect -9509 -27632 -9489 -27568
rect -15788 -27648 -9489 -27632
rect -15788 -27712 -9573 -27648
rect -9509 -27712 -9489 -27648
rect -15788 -27728 -9489 -27712
rect -15788 -27792 -9573 -27728
rect -9509 -27792 -9489 -27728
rect -15788 -27808 -9489 -27792
rect -15788 -27872 -9573 -27808
rect -9509 -27872 -9489 -27808
rect -15788 -27888 -9489 -27872
rect -15788 -27952 -9573 -27888
rect -9509 -27952 -9489 -27888
rect -15788 -27968 -9489 -27952
rect -15788 -28032 -9573 -27968
rect -9509 -28032 -9489 -27968
rect -15788 -28048 -9489 -28032
rect -15788 -28112 -9573 -28048
rect -9509 -28112 -9489 -28048
rect -15788 -28128 -9489 -28112
rect -15788 -28192 -9573 -28128
rect -9509 -28192 -9489 -28128
rect -15788 -28208 -9489 -28192
rect -15788 -28272 -9573 -28208
rect -9509 -28272 -9489 -28208
rect -15788 -28300 -9489 -28272
rect -9469 -22128 -3170 -22100
rect -9469 -22192 -3254 -22128
rect -3190 -22192 -3170 -22128
rect -9469 -22208 -3170 -22192
rect -9469 -22272 -3254 -22208
rect -3190 -22272 -3170 -22208
rect -9469 -22288 -3170 -22272
rect -9469 -22352 -3254 -22288
rect -3190 -22352 -3170 -22288
rect -9469 -22368 -3170 -22352
rect -9469 -22432 -3254 -22368
rect -3190 -22432 -3170 -22368
rect -9469 -22448 -3170 -22432
rect -9469 -22512 -3254 -22448
rect -3190 -22512 -3170 -22448
rect -9469 -22528 -3170 -22512
rect -9469 -22592 -3254 -22528
rect -3190 -22592 -3170 -22528
rect -9469 -22608 -3170 -22592
rect -9469 -22672 -3254 -22608
rect -3190 -22672 -3170 -22608
rect -9469 -22688 -3170 -22672
rect -9469 -22752 -3254 -22688
rect -3190 -22752 -3170 -22688
rect -9469 -22768 -3170 -22752
rect -9469 -22832 -3254 -22768
rect -3190 -22832 -3170 -22768
rect -9469 -22848 -3170 -22832
rect -9469 -22912 -3254 -22848
rect -3190 -22912 -3170 -22848
rect -9469 -22928 -3170 -22912
rect -9469 -22992 -3254 -22928
rect -3190 -22992 -3170 -22928
rect -9469 -23008 -3170 -22992
rect -9469 -23072 -3254 -23008
rect -3190 -23072 -3170 -23008
rect -9469 -23088 -3170 -23072
rect -9469 -23152 -3254 -23088
rect -3190 -23152 -3170 -23088
rect -9469 -23168 -3170 -23152
rect -9469 -23232 -3254 -23168
rect -3190 -23232 -3170 -23168
rect -9469 -23248 -3170 -23232
rect -9469 -23312 -3254 -23248
rect -3190 -23312 -3170 -23248
rect -9469 -23328 -3170 -23312
rect -9469 -23392 -3254 -23328
rect -3190 -23392 -3170 -23328
rect -9469 -23408 -3170 -23392
rect -9469 -23472 -3254 -23408
rect -3190 -23472 -3170 -23408
rect -9469 -23488 -3170 -23472
rect -9469 -23552 -3254 -23488
rect -3190 -23552 -3170 -23488
rect -9469 -23568 -3170 -23552
rect -9469 -23632 -3254 -23568
rect -3190 -23632 -3170 -23568
rect -9469 -23648 -3170 -23632
rect -9469 -23712 -3254 -23648
rect -3190 -23712 -3170 -23648
rect -9469 -23728 -3170 -23712
rect -9469 -23792 -3254 -23728
rect -3190 -23792 -3170 -23728
rect -9469 -23808 -3170 -23792
rect -9469 -23872 -3254 -23808
rect -3190 -23872 -3170 -23808
rect -9469 -23888 -3170 -23872
rect -9469 -23952 -3254 -23888
rect -3190 -23952 -3170 -23888
rect -9469 -23968 -3170 -23952
rect -9469 -24032 -3254 -23968
rect -3190 -24032 -3170 -23968
rect -9469 -24048 -3170 -24032
rect -9469 -24112 -3254 -24048
rect -3190 -24112 -3170 -24048
rect -9469 -24128 -3170 -24112
rect -9469 -24192 -3254 -24128
rect -3190 -24192 -3170 -24128
rect -9469 -24208 -3170 -24192
rect -9469 -24272 -3254 -24208
rect -3190 -24272 -3170 -24208
rect -9469 -24288 -3170 -24272
rect -9469 -24352 -3254 -24288
rect -3190 -24352 -3170 -24288
rect -9469 -24368 -3170 -24352
rect -9469 -24432 -3254 -24368
rect -3190 -24432 -3170 -24368
rect -9469 -24448 -3170 -24432
rect -9469 -24512 -3254 -24448
rect -3190 -24512 -3170 -24448
rect -9469 -24528 -3170 -24512
rect -9469 -24592 -3254 -24528
rect -3190 -24592 -3170 -24528
rect -9469 -24608 -3170 -24592
rect -9469 -24672 -3254 -24608
rect -3190 -24672 -3170 -24608
rect -9469 -24688 -3170 -24672
rect -9469 -24752 -3254 -24688
rect -3190 -24752 -3170 -24688
rect -9469 -24768 -3170 -24752
rect -9469 -24832 -3254 -24768
rect -3190 -24832 -3170 -24768
rect -9469 -24848 -3170 -24832
rect -9469 -24912 -3254 -24848
rect -3190 -24912 -3170 -24848
rect -9469 -24928 -3170 -24912
rect -9469 -24992 -3254 -24928
rect -3190 -24992 -3170 -24928
rect -9469 -25008 -3170 -24992
rect -9469 -25072 -3254 -25008
rect -3190 -25072 -3170 -25008
rect -9469 -25088 -3170 -25072
rect -9469 -25152 -3254 -25088
rect -3190 -25152 -3170 -25088
rect -9469 -25168 -3170 -25152
rect -9469 -25232 -3254 -25168
rect -3190 -25232 -3170 -25168
rect -9469 -25248 -3170 -25232
rect -9469 -25312 -3254 -25248
rect -3190 -25312 -3170 -25248
rect -9469 -25328 -3170 -25312
rect -9469 -25392 -3254 -25328
rect -3190 -25392 -3170 -25328
rect -9469 -25408 -3170 -25392
rect -9469 -25472 -3254 -25408
rect -3190 -25472 -3170 -25408
rect -9469 -25488 -3170 -25472
rect -9469 -25552 -3254 -25488
rect -3190 -25552 -3170 -25488
rect -9469 -25568 -3170 -25552
rect -9469 -25632 -3254 -25568
rect -3190 -25632 -3170 -25568
rect -9469 -25648 -3170 -25632
rect -9469 -25712 -3254 -25648
rect -3190 -25712 -3170 -25648
rect -9469 -25728 -3170 -25712
rect -9469 -25792 -3254 -25728
rect -3190 -25792 -3170 -25728
rect -9469 -25808 -3170 -25792
rect -9469 -25872 -3254 -25808
rect -3190 -25872 -3170 -25808
rect -9469 -25888 -3170 -25872
rect -9469 -25952 -3254 -25888
rect -3190 -25952 -3170 -25888
rect -9469 -25968 -3170 -25952
rect -9469 -26032 -3254 -25968
rect -3190 -26032 -3170 -25968
rect -9469 -26048 -3170 -26032
rect -9469 -26112 -3254 -26048
rect -3190 -26112 -3170 -26048
rect -9469 -26128 -3170 -26112
rect -9469 -26192 -3254 -26128
rect -3190 -26192 -3170 -26128
rect -9469 -26208 -3170 -26192
rect -9469 -26272 -3254 -26208
rect -3190 -26272 -3170 -26208
rect -9469 -26288 -3170 -26272
rect -9469 -26352 -3254 -26288
rect -3190 -26352 -3170 -26288
rect -9469 -26368 -3170 -26352
rect -9469 -26432 -3254 -26368
rect -3190 -26432 -3170 -26368
rect -9469 -26448 -3170 -26432
rect -9469 -26512 -3254 -26448
rect -3190 -26512 -3170 -26448
rect -9469 -26528 -3170 -26512
rect -9469 -26592 -3254 -26528
rect -3190 -26592 -3170 -26528
rect -9469 -26608 -3170 -26592
rect -9469 -26672 -3254 -26608
rect -3190 -26672 -3170 -26608
rect -9469 -26688 -3170 -26672
rect -9469 -26752 -3254 -26688
rect -3190 -26752 -3170 -26688
rect -9469 -26768 -3170 -26752
rect -9469 -26832 -3254 -26768
rect -3190 -26832 -3170 -26768
rect -9469 -26848 -3170 -26832
rect -9469 -26912 -3254 -26848
rect -3190 -26912 -3170 -26848
rect -9469 -26928 -3170 -26912
rect -9469 -26992 -3254 -26928
rect -3190 -26992 -3170 -26928
rect -9469 -27008 -3170 -26992
rect -9469 -27072 -3254 -27008
rect -3190 -27072 -3170 -27008
rect -9469 -27088 -3170 -27072
rect -9469 -27152 -3254 -27088
rect -3190 -27152 -3170 -27088
rect -9469 -27168 -3170 -27152
rect -9469 -27232 -3254 -27168
rect -3190 -27232 -3170 -27168
rect -9469 -27248 -3170 -27232
rect -9469 -27312 -3254 -27248
rect -3190 -27312 -3170 -27248
rect -9469 -27328 -3170 -27312
rect -9469 -27392 -3254 -27328
rect -3190 -27392 -3170 -27328
rect -9469 -27408 -3170 -27392
rect -9469 -27472 -3254 -27408
rect -3190 -27472 -3170 -27408
rect -9469 -27488 -3170 -27472
rect -9469 -27552 -3254 -27488
rect -3190 -27552 -3170 -27488
rect -9469 -27568 -3170 -27552
rect -9469 -27632 -3254 -27568
rect -3190 -27632 -3170 -27568
rect -9469 -27648 -3170 -27632
rect -9469 -27712 -3254 -27648
rect -3190 -27712 -3170 -27648
rect -9469 -27728 -3170 -27712
rect -9469 -27792 -3254 -27728
rect -3190 -27792 -3170 -27728
rect -9469 -27808 -3170 -27792
rect -9469 -27872 -3254 -27808
rect -3190 -27872 -3170 -27808
rect -9469 -27888 -3170 -27872
rect -9469 -27952 -3254 -27888
rect -3190 -27952 -3170 -27888
rect -9469 -27968 -3170 -27952
rect -9469 -28032 -3254 -27968
rect -3190 -28032 -3170 -27968
rect -9469 -28048 -3170 -28032
rect -9469 -28112 -3254 -28048
rect -3190 -28112 -3170 -28048
rect -9469 -28128 -3170 -28112
rect -9469 -28192 -3254 -28128
rect -3190 -28192 -3170 -28128
rect -9469 -28208 -3170 -28192
rect -9469 -28272 -3254 -28208
rect -3190 -28272 -3170 -28208
rect -9469 -28300 -3170 -28272
rect -3150 -22128 3149 -22100
rect -3150 -22192 3065 -22128
rect 3129 -22192 3149 -22128
rect -3150 -22208 3149 -22192
rect -3150 -22272 3065 -22208
rect 3129 -22272 3149 -22208
rect -3150 -22288 3149 -22272
rect -3150 -22352 3065 -22288
rect 3129 -22352 3149 -22288
rect -3150 -22368 3149 -22352
rect -3150 -22432 3065 -22368
rect 3129 -22432 3149 -22368
rect -3150 -22448 3149 -22432
rect -3150 -22512 3065 -22448
rect 3129 -22512 3149 -22448
rect -3150 -22528 3149 -22512
rect -3150 -22592 3065 -22528
rect 3129 -22592 3149 -22528
rect -3150 -22608 3149 -22592
rect -3150 -22672 3065 -22608
rect 3129 -22672 3149 -22608
rect -3150 -22688 3149 -22672
rect -3150 -22752 3065 -22688
rect 3129 -22752 3149 -22688
rect -3150 -22768 3149 -22752
rect -3150 -22832 3065 -22768
rect 3129 -22832 3149 -22768
rect -3150 -22848 3149 -22832
rect -3150 -22912 3065 -22848
rect 3129 -22912 3149 -22848
rect -3150 -22928 3149 -22912
rect -3150 -22992 3065 -22928
rect 3129 -22992 3149 -22928
rect -3150 -23008 3149 -22992
rect -3150 -23072 3065 -23008
rect 3129 -23072 3149 -23008
rect -3150 -23088 3149 -23072
rect -3150 -23152 3065 -23088
rect 3129 -23152 3149 -23088
rect -3150 -23168 3149 -23152
rect -3150 -23232 3065 -23168
rect 3129 -23232 3149 -23168
rect -3150 -23248 3149 -23232
rect -3150 -23312 3065 -23248
rect 3129 -23312 3149 -23248
rect -3150 -23328 3149 -23312
rect -3150 -23392 3065 -23328
rect 3129 -23392 3149 -23328
rect -3150 -23408 3149 -23392
rect -3150 -23472 3065 -23408
rect 3129 -23472 3149 -23408
rect -3150 -23488 3149 -23472
rect -3150 -23552 3065 -23488
rect 3129 -23552 3149 -23488
rect -3150 -23568 3149 -23552
rect -3150 -23632 3065 -23568
rect 3129 -23632 3149 -23568
rect -3150 -23648 3149 -23632
rect -3150 -23712 3065 -23648
rect 3129 -23712 3149 -23648
rect -3150 -23728 3149 -23712
rect -3150 -23792 3065 -23728
rect 3129 -23792 3149 -23728
rect -3150 -23808 3149 -23792
rect -3150 -23872 3065 -23808
rect 3129 -23872 3149 -23808
rect -3150 -23888 3149 -23872
rect -3150 -23952 3065 -23888
rect 3129 -23952 3149 -23888
rect -3150 -23968 3149 -23952
rect -3150 -24032 3065 -23968
rect 3129 -24032 3149 -23968
rect -3150 -24048 3149 -24032
rect -3150 -24112 3065 -24048
rect 3129 -24112 3149 -24048
rect -3150 -24128 3149 -24112
rect -3150 -24192 3065 -24128
rect 3129 -24192 3149 -24128
rect -3150 -24208 3149 -24192
rect -3150 -24272 3065 -24208
rect 3129 -24272 3149 -24208
rect -3150 -24288 3149 -24272
rect -3150 -24352 3065 -24288
rect 3129 -24352 3149 -24288
rect -3150 -24368 3149 -24352
rect -3150 -24432 3065 -24368
rect 3129 -24432 3149 -24368
rect -3150 -24448 3149 -24432
rect -3150 -24512 3065 -24448
rect 3129 -24512 3149 -24448
rect -3150 -24528 3149 -24512
rect -3150 -24592 3065 -24528
rect 3129 -24592 3149 -24528
rect -3150 -24608 3149 -24592
rect -3150 -24672 3065 -24608
rect 3129 -24672 3149 -24608
rect -3150 -24688 3149 -24672
rect -3150 -24752 3065 -24688
rect 3129 -24752 3149 -24688
rect -3150 -24768 3149 -24752
rect -3150 -24832 3065 -24768
rect 3129 -24832 3149 -24768
rect -3150 -24848 3149 -24832
rect -3150 -24912 3065 -24848
rect 3129 -24912 3149 -24848
rect -3150 -24928 3149 -24912
rect -3150 -24992 3065 -24928
rect 3129 -24992 3149 -24928
rect -3150 -25008 3149 -24992
rect -3150 -25072 3065 -25008
rect 3129 -25072 3149 -25008
rect -3150 -25088 3149 -25072
rect -3150 -25152 3065 -25088
rect 3129 -25152 3149 -25088
rect -3150 -25168 3149 -25152
rect -3150 -25232 3065 -25168
rect 3129 -25232 3149 -25168
rect -3150 -25248 3149 -25232
rect -3150 -25312 3065 -25248
rect 3129 -25312 3149 -25248
rect -3150 -25328 3149 -25312
rect -3150 -25392 3065 -25328
rect 3129 -25392 3149 -25328
rect -3150 -25408 3149 -25392
rect -3150 -25472 3065 -25408
rect 3129 -25472 3149 -25408
rect -3150 -25488 3149 -25472
rect -3150 -25552 3065 -25488
rect 3129 -25552 3149 -25488
rect -3150 -25568 3149 -25552
rect -3150 -25632 3065 -25568
rect 3129 -25632 3149 -25568
rect -3150 -25648 3149 -25632
rect -3150 -25712 3065 -25648
rect 3129 -25712 3149 -25648
rect -3150 -25728 3149 -25712
rect -3150 -25792 3065 -25728
rect 3129 -25792 3149 -25728
rect -3150 -25808 3149 -25792
rect -3150 -25872 3065 -25808
rect 3129 -25872 3149 -25808
rect -3150 -25888 3149 -25872
rect -3150 -25952 3065 -25888
rect 3129 -25952 3149 -25888
rect -3150 -25968 3149 -25952
rect -3150 -26032 3065 -25968
rect 3129 -26032 3149 -25968
rect -3150 -26048 3149 -26032
rect -3150 -26112 3065 -26048
rect 3129 -26112 3149 -26048
rect -3150 -26128 3149 -26112
rect -3150 -26192 3065 -26128
rect 3129 -26192 3149 -26128
rect -3150 -26208 3149 -26192
rect -3150 -26272 3065 -26208
rect 3129 -26272 3149 -26208
rect -3150 -26288 3149 -26272
rect -3150 -26352 3065 -26288
rect 3129 -26352 3149 -26288
rect -3150 -26368 3149 -26352
rect -3150 -26432 3065 -26368
rect 3129 -26432 3149 -26368
rect -3150 -26448 3149 -26432
rect -3150 -26512 3065 -26448
rect 3129 -26512 3149 -26448
rect -3150 -26528 3149 -26512
rect -3150 -26592 3065 -26528
rect 3129 -26592 3149 -26528
rect -3150 -26608 3149 -26592
rect -3150 -26672 3065 -26608
rect 3129 -26672 3149 -26608
rect -3150 -26688 3149 -26672
rect -3150 -26752 3065 -26688
rect 3129 -26752 3149 -26688
rect -3150 -26768 3149 -26752
rect -3150 -26832 3065 -26768
rect 3129 -26832 3149 -26768
rect -3150 -26848 3149 -26832
rect -3150 -26912 3065 -26848
rect 3129 -26912 3149 -26848
rect -3150 -26928 3149 -26912
rect -3150 -26992 3065 -26928
rect 3129 -26992 3149 -26928
rect -3150 -27008 3149 -26992
rect -3150 -27072 3065 -27008
rect 3129 -27072 3149 -27008
rect -3150 -27088 3149 -27072
rect -3150 -27152 3065 -27088
rect 3129 -27152 3149 -27088
rect -3150 -27168 3149 -27152
rect -3150 -27232 3065 -27168
rect 3129 -27232 3149 -27168
rect -3150 -27248 3149 -27232
rect -3150 -27312 3065 -27248
rect 3129 -27312 3149 -27248
rect -3150 -27328 3149 -27312
rect -3150 -27392 3065 -27328
rect 3129 -27392 3149 -27328
rect -3150 -27408 3149 -27392
rect -3150 -27472 3065 -27408
rect 3129 -27472 3149 -27408
rect -3150 -27488 3149 -27472
rect -3150 -27552 3065 -27488
rect 3129 -27552 3149 -27488
rect -3150 -27568 3149 -27552
rect -3150 -27632 3065 -27568
rect 3129 -27632 3149 -27568
rect -3150 -27648 3149 -27632
rect -3150 -27712 3065 -27648
rect 3129 -27712 3149 -27648
rect -3150 -27728 3149 -27712
rect -3150 -27792 3065 -27728
rect 3129 -27792 3149 -27728
rect -3150 -27808 3149 -27792
rect -3150 -27872 3065 -27808
rect 3129 -27872 3149 -27808
rect -3150 -27888 3149 -27872
rect -3150 -27952 3065 -27888
rect 3129 -27952 3149 -27888
rect -3150 -27968 3149 -27952
rect -3150 -28032 3065 -27968
rect 3129 -28032 3149 -27968
rect -3150 -28048 3149 -28032
rect -3150 -28112 3065 -28048
rect 3129 -28112 3149 -28048
rect -3150 -28128 3149 -28112
rect -3150 -28192 3065 -28128
rect 3129 -28192 3149 -28128
rect -3150 -28208 3149 -28192
rect -3150 -28272 3065 -28208
rect 3129 -28272 3149 -28208
rect -3150 -28300 3149 -28272
rect 3169 -22128 9468 -22100
rect 3169 -22192 9384 -22128
rect 9448 -22192 9468 -22128
rect 3169 -22208 9468 -22192
rect 3169 -22272 9384 -22208
rect 9448 -22272 9468 -22208
rect 3169 -22288 9468 -22272
rect 3169 -22352 9384 -22288
rect 9448 -22352 9468 -22288
rect 3169 -22368 9468 -22352
rect 3169 -22432 9384 -22368
rect 9448 -22432 9468 -22368
rect 3169 -22448 9468 -22432
rect 3169 -22512 9384 -22448
rect 9448 -22512 9468 -22448
rect 3169 -22528 9468 -22512
rect 3169 -22592 9384 -22528
rect 9448 -22592 9468 -22528
rect 3169 -22608 9468 -22592
rect 3169 -22672 9384 -22608
rect 9448 -22672 9468 -22608
rect 3169 -22688 9468 -22672
rect 3169 -22752 9384 -22688
rect 9448 -22752 9468 -22688
rect 3169 -22768 9468 -22752
rect 3169 -22832 9384 -22768
rect 9448 -22832 9468 -22768
rect 3169 -22848 9468 -22832
rect 3169 -22912 9384 -22848
rect 9448 -22912 9468 -22848
rect 3169 -22928 9468 -22912
rect 3169 -22992 9384 -22928
rect 9448 -22992 9468 -22928
rect 3169 -23008 9468 -22992
rect 3169 -23072 9384 -23008
rect 9448 -23072 9468 -23008
rect 3169 -23088 9468 -23072
rect 3169 -23152 9384 -23088
rect 9448 -23152 9468 -23088
rect 3169 -23168 9468 -23152
rect 3169 -23232 9384 -23168
rect 9448 -23232 9468 -23168
rect 3169 -23248 9468 -23232
rect 3169 -23312 9384 -23248
rect 9448 -23312 9468 -23248
rect 3169 -23328 9468 -23312
rect 3169 -23392 9384 -23328
rect 9448 -23392 9468 -23328
rect 3169 -23408 9468 -23392
rect 3169 -23472 9384 -23408
rect 9448 -23472 9468 -23408
rect 3169 -23488 9468 -23472
rect 3169 -23552 9384 -23488
rect 9448 -23552 9468 -23488
rect 3169 -23568 9468 -23552
rect 3169 -23632 9384 -23568
rect 9448 -23632 9468 -23568
rect 3169 -23648 9468 -23632
rect 3169 -23712 9384 -23648
rect 9448 -23712 9468 -23648
rect 3169 -23728 9468 -23712
rect 3169 -23792 9384 -23728
rect 9448 -23792 9468 -23728
rect 3169 -23808 9468 -23792
rect 3169 -23872 9384 -23808
rect 9448 -23872 9468 -23808
rect 3169 -23888 9468 -23872
rect 3169 -23952 9384 -23888
rect 9448 -23952 9468 -23888
rect 3169 -23968 9468 -23952
rect 3169 -24032 9384 -23968
rect 9448 -24032 9468 -23968
rect 3169 -24048 9468 -24032
rect 3169 -24112 9384 -24048
rect 9448 -24112 9468 -24048
rect 3169 -24128 9468 -24112
rect 3169 -24192 9384 -24128
rect 9448 -24192 9468 -24128
rect 3169 -24208 9468 -24192
rect 3169 -24272 9384 -24208
rect 9448 -24272 9468 -24208
rect 3169 -24288 9468 -24272
rect 3169 -24352 9384 -24288
rect 9448 -24352 9468 -24288
rect 3169 -24368 9468 -24352
rect 3169 -24432 9384 -24368
rect 9448 -24432 9468 -24368
rect 3169 -24448 9468 -24432
rect 3169 -24512 9384 -24448
rect 9448 -24512 9468 -24448
rect 3169 -24528 9468 -24512
rect 3169 -24592 9384 -24528
rect 9448 -24592 9468 -24528
rect 3169 -24608 9468 -24592
rect 3169 -24672 9384 -24608
rect 9448 -24672 9468 -24608
rect 3169 -24688 9468 -24672
rect 3169 -24752 9384 -24688
rect 9448 -24752 9468 -24688
rect 3169 -24768 9468 -24752
rect 3169 -24832 9384 -24768
rect 9448 -24832 9468 -24768
rect 3169 -24848 9468 -24832
rect 3169 -24912 9384 -24848
rect 9448 -24912 9468 -24848
rect 3169 -24928 9468 -24912
rect 3169 -24992 9384 -24928
rect 9448 -24992 9468 -24928
rect 3169 -25008 9468 -24992
rect 3169 -25072 9384 -25008
rect 9448 -25072 9468 -25008
rect 3169 -25088 9468 -25072
rect 3169 -25152 9384 -25088
rect 9448 -25152 9468 -25088
rect 3169 -25168 9468 -25152
rect 3169 -25232 9384 -25168
rect 9448 -25232 9468 -25168
rect 3169 -25248 9468 -25232
rect 3169 -25312 9384 -25248
rect 9448 -25312 9468 -25248
rect 3169 -25328 9468 -25312
rect 3169 -25392 9384 -25328
rect 9448 -25392 9468 -25328
rect 3169 -25408 9468 -25392
rect 3169 -25472 9384 -25408
rect 9448 -25472 9468 -25408
rect 3169 -25488 9468 -25472
rect 3169 -25552 9384 -25488
rect 9448 -25552 9468 -25488
rect 3169 -25568 9468 -25552
rect 3169 -25632 9384 -25568
rect 9448 -25632 9468 -25568
rect 3169 -25648 9468 -25632
rect 3169 -25712 9384 -25648
rect 9448 -25712 9468 -25648
rect 3169 -25728 9468 -25712
rect 3169 -25792 9384 -25728
rect 9448 -25792 9468 -25728
rect 3169 -25808 9468 -25792
rect 3169 -25872 9384 -25808
rect 9448 -25872 9468 -25808
rect 3169 -25888 9468 -25872
rect 3169 -25952 9384 -25888
rect 9448 -25952 9468 -25888
rect 3169 -25968 9468 -25952
rect 3169 -26032 9384 -25968
rect 9448 -26032 9468 -25968
rect 3169 -26048 9468 -26032
rect 3169 -26112 9384 -26048
rect 9448 -26112 9468 -26048
rect 3169 -26128 9468 -26112
rect 3169 -26192 9384 -26128
rect 9448 -26192 9468 -26128
rect 3169 -26208 9468 -26192
rect 3169 -26272 9384 -26208
rect 9448 -26272 9468 -26208
rect 3169 -26288 9468 -26272
rect 3169 -26352 9384 -26288
rect 9448 -26352 9468 -26288
rect 3169 -26368 9468 -26352
rect 3169 -26432 9384 -26368
rect 9448 -26432 9468 -26368
rect 3169 -26448 9468 -26432
rect 3169 -26512 9384 -26448
rect 9448 -26512 9468 -26448
rect 3169 -26528 9468 -26512
rect 3169 -26592 9384 -26528
rect 9448 -26592 9468 -26528
rect 3169 -26608 9468 -26592
rect 3169 -26672 9384 -26608
rect 9448 -26672 9468 -26608
rect 3169 -26688 9468 -26672
rect 3169 -26752 9384 -26688
rect 9448 -26752 9468 -26688
rect 3169 -26768 9468 -26752
rect 3169 -26832 9384 -26768
rect 9448 -26832 9468 -26768
rect 3169 -26848 9468 -26832
rect 3169 -26912 9384 -26848
rect 9448 -26912 9468 -26848
rect 3169 -26928 9468 -26912
rect 3169 -26992 9384 -26928
rect 9448 -26992 9468 -26928
rect 3169 -27008 9468 -26992
rect 3169 -27072 9384 -27008
rect 9448 -27072 9468 -27008
rect 3169 -27088 9468 -27072
rect 3169 -27152 9384 -27088
rect 9448 -27152 9468 -27088
rect 3169 -27168 9468 -27152
rect 3169 -27232 9384 -27168
rect 9448 -27232 9468 -27168
rect 3169 -27248 9468 -27232
rect 3169 -27312 9384 -27248
rect 9448 -27312 9468 -27248
rect 3169 -27328 9468 -27312
rect 3169 -27392 9384 -27328
rect 9448 -27392 9468 -27328
rect 3169 -27408 9468 -27392
rect 3169 -27472 9384 -27408
rect 9448 -27472 9468 -27408
rect 3169 -27488 9468 -27472
rect 3169 -27552 9384 -27488
rect 9448 -27552 9468 -27488
rect 3169 -27568 9468 -27552
rect 3169 -27632 9384 -27568
rect 9448 -27632 9468 -27568
rect 3169 -27648 9468 -27632
rect 3169 -27712 9384 -27648
rect 9448 -27712 9468 -27648
rect 3169 -27728 9468 -27712
rect 3169 -27792 9384 -27728
rect 9448 -27792 9468 -27728
rect 3169 -27808 9468 -27792
rect 3169 -27872 9384 -27808
rect 9448 -27872 9468 -27808
rect 3169 -27888 9468 -27872
rect 3169 -27952 9384 -27888
rect 9448 -27952 9468 -27888
rect 3169 -27968 9468 -27952
rect 3169 -28032 9384 -27968
rect 9448 -28032 9468 -27968
rect 3169 -28048 9468 -28032
rect 3169 -28112 9384 -28048
rect 9448 -28112 9468 -28048
rect 3169 -28128 9468 -28112
rect 3169 -28192 9384 -28128
rect 9448 -28192 9468 -28128
rect 3169 -28208 9468 -28192
rect 3169 -28272 9384 -28208
rect 9448 -28272 9468 -28208
rect 3169 -28300 9468 -28272
rect 9488 -22128 15787 -22100
rect 9488 -22192 15703 -22128
rect 15767 -22192 15787 -22128
rect 9488 -22208 15787 -22192
rect 9488 -22272 15703 -22208
rect 15767 -22272 15787 -22208
rect 9488 -22288 15787 -22272
rect 9488 -22352 15703 -22288
rect 15767 -22352 15787 -22288
rect 9488 -22368 15787 -22352
rect 9488 -22432 15703 -22368
rect 15767 -22432 15787 -22368
rect 9488 -22448 15787 -22432
rect 9488 -22512 15703 -22448
rect 15767 -22512 15787 -22448
rect 9488 -22528 15787 -22512
rect 9488 -22592 15703 -22528
rect 15767 -22592 15787 -22528
rect 9488 -22608 15787 -22592
rect 9488 -22672 15703 -22608
rect 15767 -22672 15787 -22608
rect 9488 -22688 15787 -22672
rect 9488 -22752 15703 -22688
rect 15767 -22752 15787 -22688
rect 9488 -22768 15787 -22752
rect 9488 -22832 15703 -22768
rect 15767 -22832 15787 -22768
rect 9488 -22848 15787 -22832
rect 9488 -22912 15703 -22848
rect 15767 -22912 15787 -22848
rect 9488 -22928 15787 -22912
rect 9488 -22992 15703 -22928
rect 15767 -22992 15787 -22928
rect 9488 -23008 15787 -22992
rect 9488 -23072 15703 -23008
rect 15767 -23072 15787 -23008
rect 9488 -23088 15787 -23072
rect 9488 -23152 15703 -23088
rect 15767 -23152 15787 -23088
rect 9488 -23168 15787 -23152
rect 9488 -23232 15703 -23168
rect 15767 -23232 15787 -23168
rect 9488 -23248 15787 -23232
rect 9488 -23312 15703 -23248
rect 15767 -23312 15787 -23248
rect 9488 -23328 15787 -23312
rect 9488 -23392 15703 -23328
rect 15767 -23392 15787 -23328
rect 9488 -23408 15787 -23392
rect 9488 -23472 15703 -23408
rect 15767 -23472 15787 -23408
rect 9488 -23488 15787 -23472
rect 9488 -23552 15703 -23488
rect 15767 -23552 15787 -23488
rect 9488 -23568 15787 -23552
rect 9488 -23632 15703 -23568
rect 15767 -23632 15787 -23568
rect 9488 -23648 15787 -23632
rect 9488 -23712 15703 -23648
rect 15767 -23712 15787 -23648
rect 9488 -23728 15787 -23712
rect 9488 -23792 15703 -23728
rect 15767 -23792 15787 -23728
rect 9488 -23808 15787 -23792
rect 9488 -23872 15703 -23808
rect 15767 -23872 15787 -23808
rect 9488 -23888 15787 -23872
rect 9488 -23952 15703 -23888
rect 15767 -23952 15787 -23888
rect 9488 -23968 15787 -23952
rect 9488 -24032 15703 -23968
rect 15767 -24032 15787 -23968
rect 9488 -24048 15787 -24032
rect 9488 -24112 15703 -24048
rect 15767 -24112 15787 -24048
rect 9488 -24128 15787 -24112
rect 9488 -24192 15703 -24128
rect 15767 -24192 15787 -24128
rect 9488 -24208 15787 -24192
rect 9488 -24272 15703 -24208
rect 15767 -24272 15787 -24208
rect 9488 -24288 15787 -24272
rect 9488 -24352 15703 -24288
rect 15767 -24352 15787 -24288
rect 9488 -24368 15787 -24352
rect 9488 -24432 15703 -24368
rect 15767 -24432 15787 -24368
rect 9488 -24448 15787 -24432
rect 9488 -24512 15703 -24448
rect 15767 -24512 15787 -24448
rect 9488 -24528 15787 -24512
rect 9488 -24592 15703 -24528
rect 15767 -24592 15787 -24528
rect 9488 -24608 15787 -24592
rect 9488 -24672 15703 -24608
rect 15767 -24672 15787 -24608
rect 9488 -24688 15787 -24672
rect 9488 -24752 15703 -24688
rect 15767 -24752 15787 -24688
rect 9488 -24768 15787 -24752
rect 9488 -24832 15703 -24768
rect 15767 -24832 15787 -24768
rect 9488 -24848 15787 -24832
rect 9488 -24912 15703 -24848
rect 15767 -24912 15787 -24848
rect 9488 -24928 15787 -24912
rect 9488 -24992 15703 -24928
rect 15767 -24992 15787 -24928
rect 9488 -25008 15787 -24992
rect 9488 -25072 15703 -25008
rect 15767 -25072 15787 -25008
rect 9488 -25088 15787 -25072
rect 9488 -25152 15703 -25088
rect 15767 -25152 15787 -25088
rect 9488 -25168 15787 -25152
rect 9488 -25232 15703 -25168
rect 15767 -25232 15787 -25168
rect 9488 -25248 15787 -25232
rect 9488 -25312 15703 -25248
rect 15767 -25312 15787 -25248
rect 9488 -25328 15787 -25312
rect 9488 -25392 15703 -25328
rect 15767 -25392 15787 -25328
rect 9488 -25408 15787 -25392
rect 9488 -25472 15703 -25408
rect 15767 -25472 15787 -25408
rect 9488 -25488 15787 -25472
rect 9488 -25552 15703 -25488
rect 15767 -25552 15787 -25488
rect 9488 -25568 15787 -25552
rect 9488 -25632 15703 -25568
rect 15767 -25632 15787 -25568
rect 9488 -25648 15787 -25632
rect 9488 -25712 15703 -25648
rect 15767 -25712 15787 -25648
rect 9488 -25728 15787 -25712
rect 9488 -25792 15703 -25728
rect 15767 -25792 15787 -25728
rect 9488 -25808 15787 -25792
rect 9488 -25872 15703 -25808
rect 15767 -25872 15787 -25808
rect 9488 -25888 15787 -25872
rect 9488 -25952 15703 -25888
rect 15767 -25952 15787 -25888
rect 9488 -25968 15787 -25952
rect 9488 -26032 15703 -25968
rect 15767 -26032 15787 -25968
rect 9488 -26048 15787 -26032
rect 9488 -26112 15703 -26048
rect 15767 -26112 15787 -26048
rect 9488 -26128 15787 -26112
rect 9488 -26192 15703 -26128
rect 15767 -26192 15787 -26128
rect 9488 -26208 15787 -26192
rect 9488 -26272 15703 -26208
rect 15767 -26272 15787 -26208
rect 9488 -26288 15787 -26272
rect 9488 -26352 15703 -26288
rect 15767 -26352 15787 -26288
rect 9488 -26368 15787 -26352
rect 9488 -26432 15703 -26368
rect 15767 -26432 15787 -26368
rect 9488 -26448 15787 -26432
rect 9488 -26512 15703 -26448
rect 15767 -26512 15787 -26448
rect 9488 -26528 15787 -26512
rect 9488 -26592 15703 -26528
rect 15767 -26592 15787 -26528
rect 9488 -26608 15787 -26592
rect 9488 -26672 15703 -26608
rect 15767 -26672 15787 -26608
rect 9488 -26688 15787 -26672
rect 9488 -26752 15703 -26688
rect 15767 -26752 15787 -26688
rect 9488 -26768 15787 -26752
rect 9488 -26832 15703 -26768
rect 15767 -26832 15787 -26768
rect 9488 -26848 15787 -26832
rect 9488 -26912 15703 -26848
rect 15767 -26912 15787 -26848
rect 9488 -26928 15787 -26912
rect 9488 -26992 15703 -26928
rect 15767 -26992 15787 -26928
rect 9488 -27008 15787 -26992
rect 9488 -27072 15703 -27008
rect 15767 -27072 15787 -27008
rect 9488 -27088 15787 -27072
rect 9488 -27152 15703 -27088
rect 15767 -27152 15787 -27088
rect 9488 -27168 15787 -27152
rect 9488 -27232 15703 -27168
rect 15767 -27232 15787 -27168
rect 9488 -27248 15787 -27232
rect 9488 -27312 15703 -27248
rect 15767 -27312 15787 -27248
rect 9488 -27328 15787 -27312
rect 9488 -27392 15703 -27328
rect 15767 -27392 15787 -27328
rect 9488 -27408 15787 -27392
rect 9488 -27472 15703 -27408
rect 15767 -27472 15787 -27408
rect 9488 -27488 15787 -27472
rect 9488 -27552 15703 -27488
rect 15767 -27552 15787 -27488
rect 9488 -27568 15787 -27552
rect 9488 -27632 15703 -27568
rect 15767 -27632 15787 -27568
rect 9488 -27648 15787 -27632
rect 9488 -27712 15703 -27648
rect 15767 -27712 15787 -27648
rect 9488 -27728 15787 -27712
rect 9488 -27792 15703 -27728
rect 15767 -27792 15787 -27728
rect 9488 -27808 15787 -27792
rect 9488 -27872 15703 -27808
rect 15767 -27872 15787 -27808
rect 9488 -27888 15787 -27872
rect 9488 -27952 15703 -27888
rect 15767 -27952 15787 -27888
rect 9488 -27968 15787 -27952
rect 9488 -28032 15703 -27968
rect 15767 -28032 15787 -27968
rect 9488 -28048 15787 -28032
rect 9488 -28112 15703 -28048
rect 15767 -28112 15787 -28048
rect 9488 -28128 15787 -28112
rect 9488 -28192 15703 -28128
rect 15767 -28192 15787 -28128
rect 9488 -28208 15787 -28192
rect 9488 -28272 15703 -28208
rect 15767 -28272 15787 -28208
rect 9488 -28300 15787 -28272
rect 15807 -22128 22106 -22100
rect 15807 -22192 22022 -22128
rect 22086 -22192 22106 -22128
rect 15807 -22208 22106 -22192
rect 15807 -22272 22022 -22208
rect 22086 -22272 22106 -22208
rect 15807 -22288 22106 -22272
rect 15807 -22352 22022 -22288
rect 22086 -22352 22106 -22288
rect 15807 -22368 22106 -22352
rect 15807 -22432 22022 -22368
rect 22086 -22432 22106 -22368
rect 15807 -22448 22106 -22432
rect 15807 -22512 22022 -22448
rect 22086 -22512 22106 -22448
rect 15807 -22528 22106 -22512
rect 15807 -22592 22022 -22528
rect 22086 -22592 22106 -22528
rect 15807 -22608 22106 -22592
rect 15807 -22672 22022 -22608
rect 22086 -22672 22106 -22608
rect 15807 -22688 22106 -22672
rect 15807 -22752 22022 -22688
rect 22086 -22752 22106 -22688
rect 15807 -22768 22106 -22752
rect 15807 -22832 22022 -22768
rect 22086 -22832 22106 -22768
rect 15807 -22848 22106 -22832
rect 15807 -22912 22022 -22848
rect 22086 -22912 22106 -22848
rect 15807 -22928 22106 -22912
rect 15807 -22992 22022 -22928
rect 22086 -22992 22106 -22928
rect 15807 -23008 22106 -22992
rect 15807 -23072 22022 -23008
rect 22086 -23072 22106 -23008
rect 15807 -23088 22106 -23072
rect 15807 -23152 22022 -23088
rect 22086 -23152 22106 -23088
rect 15807 -23168 22106 -23152
rect 15807 -23232 22022 -23168
rect 22086 -23232 22106 -23168
rect 15807 -23248 22106 -23232
rect 15807 -23312 22022 -23248
rect 22086 -23312 22106 -23248
rect 15807 -23328 22106 -23312
rect 15807 -23392 22022 -23328
rect 22086 -23392 22106 -23328
rect 15807 -23408 22106 -23392
rect 15807 -23472 22022 -23408
rect 22086 -23472 22106 -23408
rect 15807 -23488 22106 -23472
rect 15807 -23552 22022 -23488
rect 22086 -23552 22106 -23488
rect 15807 -23568 22106 -23552
rect 15807 -23632 22022 -23568
rect 22086 -23632 22106 -23568
rect 15807 -23648 22106 -23632
rect 15807 -23712 22022 -23648
rect 22086 -23712 22106 -23648
rect 15807 -23728 22106 -23712
rect 15807 -23792 22022 -23728
rect 22086 -23792 22106 -23728
rect 15807 -23808 22106 -23792
rect 15807 -23872 22022 -23808
rect 22086 -23872 22106 -23808
rect 15807 -23888 22106 -23872
rect 15807 -23952 22022 -23888
rect 22086 -23952 22106 -23888
rect 15807 -23968 22106 -23952
rect 15807 -24032 22022 -23968
rect 22086 -24032 22106 -23968
rect 15807 -24048 22106 -24032
rect 15807 -24112 22022 -24048
rect 22086 -24112 22106 -24048
rect 15807 -24128 22106 -24112
rect 15807 -24192 22022 -24128
rect 22086 -24192 22106 -24128
rect 15807 -24208 22106 -24192
rect 15807 -24272 22022 -24208
rect 22086 -24272 22106 -24208
rect 15807 -24288 22106 -24272
rect 15807 -24352 22022 -24288
rect 22086 -24352 22106 -24288
rect 15807 -24368 22106 -24352
rect 15807 -24432 22022 -24368
rect 22086 -24432 22106 -24368
rect 15807 -24448 22106 -24432
rect 15807 -24512 22022 -24448
rect 22086 -24512 22106 -24448
rect 15807 -24528 22106 -24512
rect 15807 -24592 22022 -24528
rect 22086 -24592 22106 -24528
rect 15807 -24608 22106 -24592
rect 15807 -24672 22022 -24608
rect 22086 -24672 22106 -24608
rect 15807 -24688 22106 -24672
rect 15807 -24752 22022 -24688
rect 22086 -24752 22106 -24688
rect 15807 -24768 22106 -24752
rect 15807 -24832 22022 -24768
rect 22086 -24832 22106 -24768
rect 15807 -24848 22106 -24832
rect 15807 -24912 22022 -24848
rect 22086 -24912 22106 -24848
rect 15807 -24928 22106 -24912
rect 15807 -24992 22022 -24928
rect 22086 -24992 22106 -24928
rect 15807 -25008 22106 -24992
rect 15807 -25072 22022 -25008
rect 22086 -25072 22106 -25008
rect 15807 -25088 22106 -25072
rect 15807 -25152 22022 -25088
rect 22086 -25152 22106 -25088
rect 15807 -25168 22106 -25152
rect 15807 -25232 22022 -25168
rect 22086 -25232 22106 -25168
rect 15807 -25248 22106 -25232
rect 15807 -25312 22022 -25248
rect 22086 -25312 22106 -25248
rect 15807 -25328 22106 -25312
rect 15807 -25392 22022 -25328
rect 22086 -25392 22106 -25328
rect 15807 -25408 22106 -25392
rect 15807 -25472 22022 -25408
rect 22086 -25472 22106 -25408
rect 15807 -25488 22106 -25472
rect 15807 -25552 22022 -25488
rect 22086 -25552 22106 -25488
rect 15807 -25568 22106 -25552
rect 15807 -25632 22022 -25568
rect 22086 -25632 22106 -25568
rect 15807 -25648 22106 -25632
rect 15807 -25712 22022 -25648
rect 22086 -25712 22106 -25648
rect 15807 -25728 22106 -25712
rect 15807 -25792 22022 -25728
rect 22086 -25792 22106 -25728
rect 15807 -25808 22106 -25792
rect 15807 -25872 22022 -25808
rect 22086 -25872 22106 -25808
rect 15807 -25888 22106 -25872
rect 15807 -25952 22022 -25888
rect 22086 -25952 22106 -25888
rect 15807 -25968 22106 -25952
rect 15807 -26032 22022 -25968
rect 22086 -26032 22106 -25968
rect 15807 -26048 22106 -26032
rect 15807 -26112 22022 -26048
rect 22086 -26112 22106 -26048
rect 15807 -26128 22106 -26112
rect 15807 -26192 22022 -26128
rect 22086 -26192 22106 -26128
rect 15807 -26208 22106 -26192
rect 15807 -26272 22022 -26208
rect 22086 -26272 22106 -26208
rect 15807 -26288 22106 -26272
rect 15807 -26352 22022 -26288
rect 22086 -26352 22106 -26288
rect 15807 -26368 22106 -26352
rect 15807 -26432 22022 -26368
rect 22086 -26432 22106 -26368
rect 15807 -26448 22106 -26432
rect 15807 -26512 22022 -26448
rect 22086 -26512 22106 -26448
rect 15807 -26528 22106 -26512
rect 15807 -26592 22022 -26528
rect 22086 -26592 22106 -26528
rect 15807 -26608 22106 -26592
rect 15807 -26672 22022 -26608
rect 22086 -26672 22106 -26608
rect 15807 -26688 22106 -26672
rect 15807 -26752 22022 -26688
rect 22086 -26752 22106 -26688
rect 15807 -26768 22106 -26752
rect 15807 -26832 22022 -26768
rect 22086 -26832 22106 -26768
rect 15807 -26848 22106 -26832
rect 15807 -26912 22022 -26848
rect 22086 -26912 22106 -26848
rect 15807 -26928 22106 -26912
rect 15807 -26992 22022 -26928
rect 22086 -26992 22106 -26928
rect 15807 -27008 22106 -26992
rect 15807 -27072 22022 -27008
rect 22086 -27072 22106 -27008
rect 15807 -27088 22106 -27072
rect 15807 -27152 22022 -27088
rect 22086 -27152 22106 -27088
rect 15807 -27168 22106 -27152
rect 15807 -27232 22022 -27168
rect 22086 -27232 22106 -27168
rect 15807 -27248 22106 -27232
rect 15807 -27312 22022 -27248
rect 22086 -27312 22106 -27248
rect 15807 -27328 22106 -27312
rect 15807 -27392 22022 -27328
rect 22086 -27392 22106 -27328
rect 15807 -27408 22106 -27392
rect 15807 -27472 22022 -27408
rect 22086 -27472 22106 -27408
rect 15807 -27488 22106 -27472
rect 15807 -27552 22022 -27488
rect 22086 -27552 22106 -27488
rect 15807 -27568 22106 -27552
rect 15807 -27632 22022 -27568
rect 22086 -27632 22106 -27568
rect 15807 -27648 22106 -27632
rect 15807 -27712 22022 -27648
rect 22086 -27712 22106 -27648
rect 15807 -27728 22106 -27712
rect 15807 -27792 22022 -27728
rect 22086 -27792 22106 -27728
rect 15807 -27808 22106 -27792
rect 15807 -27872 22022 -27808
rect 22086 -27872 22106 -27808
rect 15807 -27888 22106 -27872
rect 15807 -27952 22022 -27888
rect 22086 -27952 22106 -27888
rect 15807 -27968 22106 -27952
rect 15807 -28032 22022 -27968
rect 22086 -28032 22106 -27968
rect 15807 -28048 22106 -28032
rect 15807 -28112 22022 -28048
rect 22086 -28112 22106 -28048
rect 15807 -28128 22106 -28112
rect 15807 -28192 22022 -28128
rect 22086 -28192 22106 -28128
rect 15807 -28208 22106 -28192
rect 15807 -28272 22022 -28208
rect 22086 -28272 22106 -28208
rect 15807 -28300 22106 -28272
rect 22126 -22128 28425 -22100
rect 22126 -22192 28341 -22128
rect 28405 -22192 28425 -22128
rect 22126 -22208 28425 -22192
rect 22126 -22272 28341 -22208
rect 28405 -22272 28425 -22208
rect 22126 -22288 28425 -22272
rect 22126 -22352 28341 -22288
rect 28405 -22352 28425 -22288
rect 22126 -22368 28425 -22352
rect 22126 -22432 28341 -22368
rect 28405 -22432 28425 -22368
rect 22126 -22448 28425 -22432
rect 22126 -22512 28341 -22448
rect 28405 -22512 28425 -22448
rect 22126 -22528 28425 -22512
rect 22126 -22592 28341 -22528
rect 28405 -22592 28425 -22528
rect 22126 -22608 28425 -22592
rect 22126 -22672 28341 -22608
rect 28405 -22672 28425 -22608
rect 22126 -22688 28425 -22672
rect 22126 -22752 28341 -22688
rect 28405 -22752 28425 -22688
rect 22126 -22768 28425 -22752
rect 22126 -22832 28341 -22768
rect 28405 -22832 28425 -22768
rect 22126 -22848 28425 -22832
rect 22126 -22912 28341 -22848
rect 28405 -22912 28425 -22848
rect 22126 -22928 28425 -22912
rect 22126 -22992 28341 -22928
rect 28405 -22992 28425 -22928
rect 22126 -23008 28425 -22992
rect 22126 -23072 28341 -23008
rect 28405 -23072 28425 -23008
rect 22126 -23088 28425 -23072
rect 22126 -23152 28341 -23088
rect 28405 -23152 28425 -23088
rect 22126 -23168 28425 -23152
rect 22126 -23232 28341 -23168
rect 28405 -23232 28425 -23168
rect 22126 -23248 28425 -23232
rect 22126 -23312 28341 -23248
rect 28405 -23312 28425 -23248
rect 22126 -23328 28425 -23312
rect 22126 -23392 28341 -23328
rect 28405 -23392 28425 -23328
rect 22126 -23408 28425 -23392
rect 22126 -23472 28341 -23408
rect 28405 -23472 28425 -23408
rect 22126 -23488 28425 -23472
rect 22126 -23552 28341 -23488
rect 28405 -23552 28425 -23488
rect 22126 -23568 28425 -23552
rect 22126 -23632 28341 -23568
rect 28405 -23632 28425 -23568
rect 22126 -23648 28425 -23632
rect 22126 -23712 28341 -23648
rect 28405 -23712 28425 -23648
rect 22126 -23728 28425 -23712
rect 22126 -23792 28341 -23728
rect 28405 -23792 28425 -23728
rect 22126 -23808 28425 -23792
rect 22126 -23872 28341 -23808
rect 28405 -23872 28425 -23808
rect 22126 -23888 28425 -23872
rect 22126 -23952 28341 -23888
rect 28405 -23952 28425 -23888
rect 22126 -23968 28425 -23952
rect 22126 -24032 28341 -23968
rect 28405 -24032 28425 -23968
rect 22126 -24048 28425 -24032
rect 22126 -24112 28341 -24048
rect 28405 -24112 28425 -24048
rect 22126 -24128 28425 -24112
rect 22126 -24192 28341 -24128
rect 28405 -24192 28425 -24128
rect 22126 -24208 28425 -24192
rect 22126 -24272 28341 -24208
rect 28405 -24272 28425 -24208
rect 22126 -24288 28425 -24272
rect 22126 -24352 28341 -24288
rect 28405 -24352 28425 -24288
rect 22126 -24368 28425 -24352
rect 22126 -24432 28341 -24368
rect 28405 -24432 28425 -24368
rect 22126 -24448 28425 -24432
rect 22126 -24512 28341 -24448
rect 28405 -24512 28425 -24448
rect 22126 -24528 28425 -24512
rect 22126 -24592 28341 -24528
rect 28405 -24592 28425 -24528
rect 22126 -24608 28425 -24592
rect 22126 -24672 28341 -24608
rect 28405 -24672 28425 -24608
rect 22126 -24688 28425 -24672
rect 22126 -24752 28341 -24688
rect 28405 -24752 28425 -24688
rect 22126 -24768 28425 -24752
rect 22126 -24832 28341 -24768
rect 28405 -24832 28425 -24768
rect 22126 -24848 28425 -24832
rect 22126 -24912 28341 -24848
rect 28405 -24912 28425 -24848
rect 22126 -24928 28425 -24912
rect 22126 -24992 28341 -24928
rect 28405 -24992 28425 -24928
rect 22126 -25008 28425 -24992
rect 22126 -25072 28341 -25008
rect 28405 -25072 28425 -25008
rect 22126 -25088 28425 -25072
rect 22126 -25152 28341 -25088
rect 28405 -25152 28425 -25088
rect 22126 -25168 28425 -25152
rect 22126 -25232 28341 -25168
rect 28405 -25232 28425 -25168
rect 22126 -25248 28425 -25232
rect 22126 -25312 28341 -25248
rect 28405 -25312 28425 -25248
rect 22126 -25328 28425 -25312
rect 22126 -25392 28341 -25328
rect 28405 -25392 28425 -25328
rect 22126 -25408 28425 -25392
rect 22126 -25472 28341 -25408
rect 28405 -25472 28425 -25408
rect 22126 -25488 28425 -25472
rect 22126 -25552 28341 -25488
rect 28405 -25552 28425 -25488
rect 22126 -25568 28425 -25552
rect 22126 -25632 28341 -25568
rect 28405 -25632 28425 -25568
rect 22126 -25648 28425 -25632
rect 22126 -25712 28341 -25648
rect 28405 -25712 28425 -25648
rect 22126 -25728 28425 -25712
rect 22126 -25792 28341 -25728
rect 28405 -25792 28425 -25728
rect 22126 -25808 28425 -25792
rect 22126 -25872 28341 -25808
rect 28405 -25872 28425 -25808
rect 22126 -25888 28425 -25872
rect 22126 -25952 28341 -25888
rect 28405 -25952 28425 -25888
rect 22126 -25968 28425 -25952
rect 22126 -26032 28341 -25968
rect 28405 -26032 28425 -25968
rect 22126 -26048 28425 -26032
rect 22126 -26112 28341 -26048
rect 28405 -26112 28425 -26048
rect 22126 -26128 28425 -26112
rect 22126 -26192 28341 -26128
rect 28405 -26192 28425 -26128
rect 22126 -26208 28425 -26192
rect 22126 -26272 28341 -26208
rect 28405 -26272 28425 -26208
rect 22126 -26288 28425 -26272
rect 22126 -26352 28341 -26288
rect 28405 -26352 28425 -26288
rect 22126 -26368 28425 -26352
rect 22126 -26432 28341 -26368
rect 28405 -26432 28425 -26368
rect 22126 -26448 28425 -26432
rect 22126 -26512 28341 -26448
rect 28405 -26512 28425 -26448
rect 22126 -26528 28425 -26512
rect 22126 -26592 28341 -26528
rect 28405 -26592 28425 -26528
rect 22126 -26608 28425 -26592
rect 22126 -26672 28341 -26608
rect 28405 -26672 28425 -26608
rect 22126 -26688 28425 -26672
rect 22126 -26752 28341 -26688
rect 28405 -26752 28425 -26688
rect 22126 -26768 28425 -26752
rect 22126 -26832 28341 -26768
rect 28405 -26832 28425 -26768
rect 22126 -26848 28425 -26832
rect 22126 -26912 28341 -26848
rect 28405 -26912 28425 -26848
rect 22126 -26928 28425 -26912
rect 22126 -26992 28341 -26928
rect 28405 -26992 28425 -26928
rect 22126 -27008 28425 -26992
rect 22126 -27072 28341 -27008
rect 28405 -27072 28425 -27008
rect 22126 -27088 28425 -27072
rect 22126 -27152 28341 -27088
rect 28405 -27152 28425 -27088
rect 22126 -27168 28425 -27152
rect 22126 -27232 28341 -27168
rect 28405 -27232 28425 -27168
rect 22126 -27248 28425 -27232
rect 22126 -27312 28341 -27248
rect 28405 -27312 28425 -27248
rect 22126 -27328 28425 -27312
rect 22126 -27392 28341 -27328
rect 28405 -27392 28425 -27328
rect 22126 -27408 28425 -27392
rect 22126 -27472 28341 -27408
rect 28405 -27472 28425 -27408
rect 22126 -27488 28425 -27472
rect 22126 -27552 28341 -27488
rect 28405 -27552 28425 -27488
rect 22126 -27568 28425 -27552
rect 22126 -27632 28341 -27568
rect 28405 -27632 28425 -27568
rect 22126 -27648 28425 -27632
rect 22126 -27712 28341 -27648
rect 28405 -27712 28425 -27648
rect 22126 -27728 28425 -27712
rect 22126 -27792 28341 -27728
rect 28405 -27792 28425 -27728
rect 22126 -27808 28425 -27792
rect 22126 -27872 28341 -27808
rect 28405 -27872 28425 -27808
rect 22126 -27888 28425 -27872
rect 22126 -27952 28341 -27888
rect 28405 -27952 28425 -27888
rect 22126 -27968 28425 -27952
rect 22126 -28032 28341 -27968
rect 28405 -28032 28425 -27968
rect 22126 -28048 28425 -28032
rect 22126 -28112 28341 -28048
rect 28405 -28112 28425 -28048
rect 22126 -28128 28425 -28112
rect 22126 -28192 28341 -28128
rect 28405 -28192 28425 -28128
rect 22126 -28208 28425 -28192
rect 22126 -28272 28341 -28208
rect 28405 -28272 28425 -28208
rect 22126 -28300 28425 -28272
rect 28445 -22128 34744 -22100
rect 28445 -22192 34660 -22128
rect 34724 -22192 34744 -22128
rect 28445 -22208 34744 -22192
rect 28445 -22272 34660 -22208
rect 34724 -22272 34744 -22208
rect 28445 -22288 34744 -22272
rect 28445 -22352 34660 -22288
rect 34724 -22352 34744 -22288
rect 28445 -22368 34744 -22352
rect 28445 -22432 34660 -22368
rect 34724 -22432 34744 -22368
rect 28445 -22448 34744 -22432
rect 28445 -22512 34660 -22448
rect 34724 -22512 34744 -22448
rect 28445 -22528 34744 -22512
rect 28445 -22592 34660 -22528
rect 34724 -22592 34744 -22528
rect 28445 -22608 34744 -22592
rect 28445 -22672 34660 -22608
rect 34724 -22672 34744 -22608
rect 28445 -22688 34744 -22672
rect 28445 -22752 34660 -22688
rect 34724 -22752 34744 -22688
rect 28445 -22768 34744 -22752
rect 28445 -22832 34660 -22768
rect 34724 -22832 34744 -22768
rect 28445 -22848 34744 -22832
rect 28445 -22912 34660 -22848
rect 34724 -22912 34744 -22848
rect 28445 -22928 34744 -22912
rect 28445 -22992 34660 -22928
rect 34724 -22992 34744 -22928
rect 28445 -23008 34744 -22992
rect 28445 -23072 34660 -23008
rect 34724 -23072 34744 -23008
rect 28445 -23088 34744 -23072
rect 28445 -23152 34660 -23088
rect 34724 -23152 34744 -23088
rect 28445 -23168 34744 -23152
rect 28445 -23232 34660 -23168
rect 34724 -23232 34744 -23168
rect 28445 -23248 34744 -23232
rect 28445 -23312 34660 -23248
rect 34724 -23312 34744 -23248
rect 28445 -23328 34744 -23312
rect 28445 -23392 34660 -23328
rect 34724 -23392 34744 -23328
rect 28445 -23408 34744 -23392
rect 28445 -23472 34660 -23408
rect 34724 -23472 34744 -23408
rect 28445 -23488 34744 -23472
rect 28445 -23552 34660 -23488
rect 34724 -23552 34744 -23488
rect 28445 -23568 34744 -23552
rect 28445 -23632 34660 -23568
rect 34724 -23632 34744 -23568
rect 28445 -23648 34744 -23632
rect 28445 -23712 34660 -23648
rect 34724 -23712 34744 -23648
rect 28445 -23728 34744 -23712
rect 28445 -23792 34660 -23728
rect 34724 -23792 34744 -23728
rect 28445 -23808 34744 -23792
rect 28445 -23872 34660 -23808
rect 34724 -23872 34744 -23808
rect 28445 -23888 34744 -23872
rect 28445 -23952 34660 -23888
rect 34724 -23952 34744 -23888
rect 28445 -23968 34744 -23952
rect 28445 -24032 34660 -23968
rect 34724 -24032 34744 -23968
rect 28445 -24048 34744 -24032
rect 28445 -24112 34660 -24048
rect 34724 -24112 34744 -24048
rect 28445 -24128 34744 -24112
rect 28445 -24192 34660 -24128
rect 34724 -24192 34744 -24128
rect 28445 -24208 34744 -24192
rect 28445 -24272 34660 -24208
rect 34724 -24272 34744 -24208
rect 28445 -24288 34744 -24272
rect 28445 -24352 34660 -24288
rect 34724 -24352 34744 -24288
rect 28445 -24368 34744 -24352
rect 28445 -24432 34660 -24368
rect 34724 -24432 34744 -24368
rect 28445 -24448 34744 -24432
rect 28445 -24512 34660 -24448
rect 34724 -24512 34744 -24448
rect 28445 -24528 34744 -24512
rect 28445 -24592 34660 -24528
rect 34724 -24592 34744 -24528
rect 28445 -24608 34744 -24592
rect 28445 -24672 34660 -24608
rect 34724 -24672 34744 -24608
rect 28445 -24688 34744 -24672
rect 28445 -24752 34660 -24688
rect 34724 -24752 34744 -24688
rect 28445 -24768 34744 -24752
rect 28445 -24832 34660 -24768
rect 34724 -24832 34744 -24768
rect 28445 -24848 34744 -24832
rect 28445 -24912 34660 -24848
rect 34724 -24912 34744 -24848
rect 28445 -24928 34744 -24912
rect 28445 -24992 34660 -24928
rect 34724 -24992 34744 -24928
rect 28445 -25008 34744 -24992
rect 28445 -25072 34660 -25008
rect 34724 -25072 34744 -25008
rect 28445 -25088 34744 -25072
rect 28445 -25152 34660 -25088
rect 34724 -25152 34744 -25088
rect 28445 -25168 34744 -25152
rect 28445 -25232 34660 -25168
rect 34724 -25232 34744 -25168
rect 28445 -25248 34744 -25232
rect 28445 -25312 34660 -25248
rect 34724 -25312 34744 -25248
rect 28445 -25328 34744 -25312
rect 28445 -25392 34660 -25328
rect 34724 -25392 34744 -25328
rect 28445 -25408 34744 -25392
rect 28445 -25472 34660 -25408
rect 34724 -25472 34744 -25408
rect 28445 -25488 34744 -25472
rect 28445 -25552 34660 -25488
rect 34724 -25552 34744 -25488
rect 28445 -25568 34744 -25552
rect 28445 -25632 34660 -25568
rect 34724 -25632 34744 -25568
rect 28445 -25648 34744 -25632
rect 28445 -25712 34660 -25648
rect 34724 -25712 34744 -25648
rect 28445 -25728 34744 -25712
rect 28445 -25792 34660 -25728
rect 34724 -25792 34744 -25728
rect 28445 -25808 34744 -25792
rect 28445 -25872 34660 -25808
rect 34724 -25872 34744 -25808
rect 28445 -25888 34744 -25872
rect 28445 -25952 34660 -25888
rect 34724 -25952 34744 -25888
rect 28445 -25968 34744 -25952
rect 28445 -26032 34660 -25968
rect 34724 -26032 34744 -25968
rect 28445 -26048 34744 -26032
rect 28445 -26112 34660 -26048
rect 34724 -26112 34744 -26048
rect 28445 -26128 34744 -26112
rect 28445 -26192 34660 -26128
rect 34724 -26192 34744 -26128
rect 28445 -26208 34744 -26192
rect 28445 -26272 34660 -26208
rect 34724 -26272 34744 -26208
rect 28445 -26288 34744 -26272
rect 28445 -26352 34660 -26288
rect 34724 -26352 34744 -26288
rect 28445 -26368 34744 -26352
rect 28445 -26432 34660 -26368
rect 34724 -26432 34744 -26368
rect 28445 -26448 34744 -26432
rect 28445 -26512 34660 -26448
rect 34724 -26512 34744 -26448
rect 28445 -26528 34744 -26512
rect 28445 -26592 34660 -26528
rect 34724 -26592 34744 -26528
rect 28445 -26608 34744 -26592
rect 28445 -26672 34660 -26608
rect 34724 -26672 34744 -26608
rect 28445 -26688 34744 -26672
rect 28445 -26752 34660 -26688
rect 34724 -26752 34744 -26688
rect 28445 -26768 34744 -26752
rect 28445 -26832 34660 -26768
rect 34724 -26832 34744 -26768
rect 28445 -26848 34744 -26832
rect 28445 -26912 34660 -26848
rect 34724 -26912 34744 -26848
rect 28445 -26928 34744 -26912
rect 28445 -26992 34660 -26928
rect 34724 -26992 34744 -26928
rect 28445 -27008 34744 -26992
rect 28445 -27072 34660 -27008
rect 34724 -27072 34744 -27008
rect 28445 -27088 34744 -27072
rect 28445 -27152 34660 -27088
rect 34724 -27152 34744 -27088
rect 28445 -27168 34744 -27152
rect 28445 -27232 34660 -27168
rect 34724 -27232 34744 -27168
rect 28445 -27248 34744 -27232
rect 28445 -27312 34660 -27248
rect 34724 -27312 34744 -27248
rect 28445 -27328 34744 -27312
rect 28445 -27392 34660 -27328
rect 34724 -27392 34744 -27328
rect 28445 -27408 34744 -27392
rect 28445 -27472 34660 -27408
rect 34724 -27472 34744 -27408
rect 28445 -27488 34744 -27472
rect 28445 -27552 34660 -27488
rect 34724 -27552 34744 -27488
rect 28445 -27568 34744 -27552
rect 28445 -27632 34660 -27568
rect 34724 -27632 34744 -27568
rect 28445 -27648 34744 -27632
rect 28445 -27712 34660 -27648
rect 34724 -27712 34744 -27648
rect 28445 -27728 34744 -27712
rect 28445 -27792 34660 -27728
rect 34724 -27792 34744 -27728
rect 28445 -27808 34744 -27792
rect 28445 -27872 34660 -27808
rect 34724 -27872 34744 -27808
rect 28445 -27888 34744 -27872
rect 28445 -27952 34660 -27888
rect 34724 -27952 34744 -27888
rect 28445 -27968 34744 -27952
rect 28445 -28032 34660 -27968
rect 34724 -28032 34744 -27968
rect 28445 -28048 34744 -28032
rect 28445 -28112 34660 -28048
rect 34724 -28112 34744 -28048
rect 28445 -28128 34744 -28112
rect 28445 -28192 34660 -28128
rect 34724 -28192 34744 -28128
rect 28445 -28208 34744 -28192
rect 28445 -28272 34660 -28208
rect 34724 -28272 34744 -28208
rect 28445 -28300 34744 -28272
rect 34764 -22128 41063 -22100
rect 34764 -22192 40979 -22128
rect 41043 -22192 41063 -22128
rect 34764 -22208 41063 -22192
rect 34764 -22272 40979 -22208
rect 41043 -22272 41063 -22208
rect 34764 -22288 41063 -22272
rect 34764 -22352 40979 -22288
rect 41043 -22352 41063 -22288
rect 34764 -22368 41063 -22352
rect 34764 -22432 40979 -22368
rect 41043 -22432 41063 -22368
rect 34764 -22448 41063 -22432
rect 34764 -22512 40979 -22448
rect 41043 -22512 41063 -22448
rect 34764 -22528 41063 -22512
rect 34764 -22592 40979 -22528
rect 41043 -22592 41063 -22528
rect 34764 -22608 41063 -22592
rect 34764 -22672 40979 -22608
rect 41043 -22672 41063 -22608
rect 34764 -22688 41063 -22672
rect 34764 -22752 40979 -22688
rect 41043 -22752 41063 -22688
rect 34764 -22768 41063 -22752
rect 34764 -22832 40979 -22768
rect 41043 -22832 41063 -22768
rect 34764 -22848 41063 -22832
rect 34764 -22912 40979 -22848
rect 41043 -22912 41063 -22848
rect 34764 -22928 41063 -22912
rect 34764 -22992 40979 -22928
rect 41043 -22992 41063 -22928
rect 34764 -23008 41063 -22992
rect 34764 -23072 40979 -23008
rect 41043 -23072 41063 -23008
rect 34764 -23088 41063 -23072
rect 34764 -23152 40979 -23088
rect 41043 -23152 41063 -23088
rect 34764 -23168 41063 -23152
rect 34764 -23232 40979 -23168
rect 41043 -23232 41063 -23168
rect 34764 -23248 41063 -23232
rect 34764 -23312 40979 -23248
rect 41043 -23312 41063 -23248
rect 34764 -23328 41063 -23312
rect 34764 -23392 40979 -23328
rect 41043 -23392 41063 -23328
rect 34764 -23408 41063 -23392
rect 34764 -23472 40979 -23408
rect 41043 -23472 41063 -23408
rect 34764 -23488 41063 -23472
rect 34764 -23552 40979 -23488
rect 41043 -23552 41063 -23488
rect 34764 -23568 41063 -23552
rect 34764 -23632 40979 -23568
rect 41043 -23632 41063 -23568
rect 34764 -23648 41063 -23632
rect 34764 -23712 40979 -23648
rect 41043 -23712 41063 -23648
rect 34764 -23728 41063 -23712
rect 34764 -23792 40979 -23728
rect 41043 -23792 41063 -23728
rect 34764 -23808 41063 -23792
rect 34764 -23872 40979 -23808
rect 41043 -23872 41063 -23808
rect 34764 -23888 41063 -23872
rect 34764 -23952 40979 -23888
rect 41043 -23952 41063 -23888
rect 34764 -23968 41063 -23952
rect 34764 -24032 40979 -23968
rect 41043 -24032 41063 -23968
rect 34764 -24048 41063 -24032
rect 34764 -24112 40979 -24048
rect 41043 -24112 41063 -24048
rect 34764 -24128 41063 -24112
rect 34764 -24192 40979 -24128
rect 41043 -24192 41063 -24128
rect 34764 -24208 41063 -24192
rect 34764 -24272 40979 -24208
rect 41043 -24272 41063 -24208
rect 34764 -24288 41063 -24272
rect 34764 -24352 40979 -24288
rect 41043 -24352 41063 -24288
rect 34764 -24368 41063 -24352
rect 34764 -24432 40979 -24368
rect 41043 -24432 41063 -24368
rect 34764 -24448 41063 -24432
rect 34764 -24512 40979 -24448
rect 41043 -24512 41063 -24448
rect 34764 -24528 41063 -24512
rect 34764 -24592 40979 -24528
rect 41043 -24592 41063 -24528
rect 34764 -24608 41063 -24592
rect 34764 -24672 40979 -24608
rect 41043 -24672 41063 -24608
rect 34764 -24688 41063 -24672
rect 34764 -24752 40979 -24688
rect 41043 -24752 41063 -24688
rect 34764 -24768 41063 -24752
rect 34764 -24832 40979 -24768
rect 41043 -24832 41063 -24768
rect 34764 -24848 41063 -24832
rect 34764 -24912 40979 -24848
rect 41043 -24912 41063 -24848
rect 34764 -24928 41063 -24912
rect 34764 -24992 40979 -24928
rect 41043 -24992 41063 -24928
rect 34764 -25008 41063 -24992
rect 34764 -25072 40979 -25008
rect 41043 -25072 41063 -25008
rect 34764 -25088 41063 -25072
rect 34764 -25152 40979 -25088
rect 41043 -25152 41063 -25088
rect 34764 -25168 41063 -25152
rect 34764 -25232 40979 -25168
rect 41043 -25232 41063 -25168
rect 34764 -25248 41063 -25232
rect 34764 -25312 40979 -25248
rect 41043 -25312 41063 -25248
rect 34764 -25328 41063 -25312
rect 34764 -25392 40979 -25328
rect 41043 -25392 41063 -25328
rect 34764 -25408 41063 -25392
rect 34764 -25472 40979 -25408
rect 41043 -25472 41063 -25408
rect 34764 -25488 41063 -25472
rect 34764 -25552 40979 -25488
rect 41043 -25552 41063 -25488
rect 34764 -25568 41063 -25552
rect 34764 -25632 40979 -25568
rect 41043 -25632 41063 -25568
rect 34764 -25648 41063 -25632
rect 34764 -25712 40979 -25648
rect 41043 -25712 41063 -25648
rect 34764 -25728 41063 -25712
rect 34764 -25792 40979 -25728
rect 41043 -25792 41063 -25728
rect 34764 -25808 41063 -25792
rect 34764 -25872 40979 -25808
rect 41043 -25872 41063 -25808
rect 34764 -25888 41063 -25872
rect 34764 -25952 40979 -25888
rect 41043 -25952 41063 -25888
rect 34764 -25968 41063 -25952
rect 34764 -26032 40979 -25968
rect 41043 -26032 41063 -25968
rect 34764 -26048 41063 -26032
rect 34764 -26112 40979 -26048
rect 41043 -26112 41063 -26048
rect 34764 -26128 41063 -26112
rect 34764 -26192 40979 -26128
rect 41043 -26192 41063 -26128
rect 34764 -26208 41063 -26192
rect 34764 -26272 40979 -26208
rect 41043 -26272 41063 -26208
rect 34764 -26288 41063 -26272
rect 34764 -26352 40979 -26288
rect 41043 -26352 41063 -26288
rect 34764 -26368 41063 -26352
rect 34764 -26432 40979 -26368
rect 41043 -26432 41063 -26368
rect 34764 -26448 41063 -26432
rect 34764 -26512 40979 -26448
rect 41043 -26512 41063 -26448
rect 34764 -26528 41063 -26512
rect 34764 -26592 40979 -26528
rect 41043 -26592 41063 -26528
rect 34764 -26608 41063 -26592
rect 34764 -26672 40979 -26608
rect 41043 -26672 41063 -26608
rect 34764 -26688 41063 -26672
rect 34764 -26752 40979 -26688
rect 41043 -26752 41063 -26688
rect 34764 -26768 41063 -26752
rect 34764 -26832 40979 -26768
rect 41043 -26832 41063 -26768
rect 34764 -26848 41063 -26832
rect 34764 -26912 40979 -26848
rect 41043 -26912 41063 -26848
rect 34764 -26928 41063 -26912
rect 34764 -26992 40979 -26928
rect 41043 -26992 41063 -26928
rect 34764 -27008 41063 -26992
rect 34764 -27072 40979 -27008
rect 41043 -27072 41063 -27008
rect 34764 -27088 41063 -27072
rect 34764 -27152 40979 -27088
rect 41043 -27152 41063 -27088
rect 34764 -27168 41063 -27152
rect 34764 -27232 40979 -27168
rect 41043 -27232 41063 -27168
rect 34764 -27248 41063 -27232
rect 34764 -27312 40979 -27248
rect 41043 -27312 41063 -27248
rect 34764 -27328 41063 -27312
rect 34764 -27392 40979 -27328
rect 41043 -27392 41063 -27328
rect 34764 -27408 41063 -27392
rect 34764 -27472 40979 -27408
rect 41043 -27472 41063 -27408
rect 34764 -27488 41063 -27472
rect 34764 -27552 40979 -27488
rect 41043 -27552 41063 -27488
rect 34764 -27568 41063 -27552
rect 34764 -27632 40979 -27568
rect 41043 -27632 41063 -27568
rect 34764 -27648 41063 -27632
rect 34764 -27712 40979 -27648
rect 41043 -27712 41063 -27648
rect 34764 -27728 41063 -27712
rect 34764 -27792 40979 -27728
rect 41043 -27792 41063 -27728
rect 34764 -27808 41063 -27792
rect 34764 -27872 40979 -27808
rect 41043 -27872 41063 -27808
rect 34764 -27888 41063 -27872
rect 34764 -27952 40979 -27888
rect 41043 -27952 41063 -27888
rect 34764 -27968 41063 -27952
rect 34764 -28032 40979 -27968
rect 41043 -28032 41063 -27968
rect 34764 -28048 41063 -28032
rect 34764 -28112 40979 -28048
rect 41043 -28112 41063 -28048
rect 34764 -28128 41063 -28112
rect 34764 -28192 40979 -28128
rect 41043 -28192 41063 -28128
rect 34764 -28208 41063 -28192
rect 34764 -28272 40979 -28208
rect 41043 -28272 41063 -28208
rect 34764 -28300 41063 -28272
rect 41083 -22128 47382 -22100
rect 41083 -22192 47298 -22128
rect 47362 -22192 47382 -22128
rect 41083 -22208 47382 -22192
rect 41083 -22272 47298 -22208
rect 47362 -22272 47382 -22208
rect 41083 -22288 47382 -22272
rect 41083 -22352 47298 -22288
rect 47362 -22352 47382 -22288
rect 41083 -22368 47382 -22352
rect 41083 -22432 47298 -22368
rect 47362 -22432 47382 -22368
rect 41083 -22448 47382 -22432
rect 41083 -22512 47298 -22448
rect 47362 -22512 47382 -22448
rect 41083 -22528 47382 -22512
rect 41083 -22592 47298 -22528
rect 47362 -22592 47382 -22528
rect 41083 -22608 47382 -22592
rect 41083 -22672 47298 -22608
rect 47362 -22672 47382 -22608
rect 41083 -22688 47382 -22672
rect 41083 -22752 47298 -22688
rect 47362 -22752 47382 -22688
rect 41083 -22768 47382 -22752
rect 41083 -22832 47298 -22768
rect 47362 -22832 47382 -22768
rect 41083 -22848 47382 -22832
rect 41083 -22912 47298 -22848
rect 47362 -22912 47382 -22848
rect 41083 -22928 47382 -22912
rect 41083 -22992 47298 -22928
rect 47362 -22992 47382 -22928
rect 41083 -23008 47382 -22992
rect 41083 -23072 47298 -23008
rect 47362 -23072 47382 -23008
rect 41083 -23088 47382 -23072
rect 41083 -23152 47298 -23088
rect 47362 -23152 47382 -23088
rect 41083 -23168 47382 -23152
rect 41083 -23232 47298 -23168
rect 47362 -23232 47382 -23168
rect 41083 -23248 47382 -23232
rect 41083 -23312 47298 -23248
rect 47362 -23312 47382 -23248
rect 41083 -23328 47382 -23312
rect 41083 -23392 47298 -23328
rect 47362 -23392 47382 -23328
rect 41083 -23408 47382 -23392
rect 41083 -23472 47298 -23408
rect 47362 -23472 47382 -23408
rect 41083 -23488 47382 -23472
rect 41083 -23552 47298 -23488
rect 47362 -23552 47382 -23488
rect 41083 -23568 47382 -23552
rect 41083 -23632 47298 -23568
rect 47362 -23632 47382 -23568
rect 41083 -23648 47382 -23632
rect 41083 -23712 47298 -23648
rect 47362 -23712 47382 -23648
rect 41083 -23728 47382 -23712
rect 41083 -23792 47298 -23728
rect 47362 -23792 47382 -23728
rect 41083 -23808 47382 -23792
rect 41083 -23872 47298 -23808
rect 47362 -23872 47382 -23808
rect 41083 -23888 47382 -23872
rect 41083 -23952 47298 -23888
rect 47362 -23952 47382 -23888
rect 41083 -23968 47382 -23952
rect 41083 -24032 47298 -23968
rect 47362 -24032 47382 -23968
rect 41083 -24048 47382 -24032
rect 41083 -24112 47298 -24048
rect 47362 -24112 47382 -24048
rect 41083 -24128 47382 -24112
rect 41083 -24192 47298 -24128
rect 47362 -24192 47382 -24128
rect 41083 -24208 47382 -24192
rect 41083 -24272 47298 -24208
rect 47362 -24272 47382 -24208
rect 41083 -24288 47382 -24272
rect 41083 -24352 47298 -24288
rect 47362 -24352 47382 -24288
rect 41083 -24368 47382 -24352
rect 41083 -24432 47298 -24368
rect 47362 -24432 47382 -24368
rect 41083 -24448 47382 -24432
rect 41083 -24512 47298 -24448
rect 47362 -24512 47382 -24448
rect 41083 -24528 47382 -24512
rect 41083 -24592 47298 -24528
rect 47362 -24592 47382 -24528
rect 41083 -24608 47382 -24592
rect 41083 -24672 47298 -24608
rect 47362 -24672 47382 -24608
rect 41083 -24688 47382 -24672
rect 41083 -24752 47298 -24688
rect 47362 -24752 47382 -24688
rect 41083 -24768 47382 -24752
rect 41083 -24832 47298 -24768
rect 47362 -24832 47382 -24768
rect 41083 -24848 47382 -24832
rect 41083 -24912 47298 -24848
rect 47362 -24912 47382 -24848
rect 41083 -24928 47382 -24912
rect 41083 -24992 47298 -24928
rect 47362 -24992 47382 -24928
rect 41083 -25008 47382 -24992
rect 41083 -25072 47298 -25008
rect 47362 -25072 47382 -25008
rect 41083 -25088 47382 -25072
rect 41083 -25152 47298 -25088
rect 47362 -25152 47382 -25088
rect 41083 -25168 47382 -25152
rect 41083 -25232 47298 -25168
rect 47362 -25232 47382 -25168
rect 41083 -25248 47382 -25232
rect 41083 -25312 47298 -25248
rect 47362 -25312 47382 -25248
rect 41083 -25328 47382 -25312
rect 41083 -25392 47298 -25328
rect 47362 -25392 47382 -25328
rect 41083 -25408 47382 -25392
rect 41083 -25472 47298 -25408
rect 47362 -25472 47382 -25408
rect 41083 -25488 47382 -25472
rect 41083 -25552 47298 -25488
rect 47362 -25552 47382 -25488
rect 41083 -25568 47382 -25552
rect 41083 -25632 47298 -25568
rect 47362 -25632 47382 -25568
rect 41083 -25648 47382 -25632
rect 41083 -25712 47298 -25648
rect 47362 -25712 47382 -25648
rect 41083 -25728 47382 -25712
rect 41083 -25792 47298 -25728
rect 47362 -25792 47382 -25728
rect 41083 -25808 47382 -25792
rect 41083 -25872 47298 -25808
rect 47362 -25872 47382 -25808
rect 41083 -25888 47382 -25872
rect 41083 -25952 47298 -25888
rect 47362 -25952 47382 -25888
rect 41083 -25968 47382 -25952
rect 41083 -26032 47298 -25968
rect 47362 -26032 47382 -25968
rect 41083 -26048 47382 -26032
rect 41083 -26112 47298 -26048
rect 47362 -26112 47382 -26048
rect 41083 -26128 47382 -26112
rect 41083 -26192 47298 -26128
rect 47362 -26192 47382 -26128
rect 41083 -26208 47382 -26192
rect 41083 -26272 47298 -26208
rect 47362 -26272 47382 -26208
rect 41083 -26288 47382 -26272
rect 41083 -26352 47298 -26288
rect 47362 -26352 47382 -26288
rect 41083 -26368 47382 -26352
rect 41083 -26432 47298 -26368
rect 47362 -26432 47382 -26368
rect 41083 -26448 47382 -26432
rect 41083 -26512 47298 -26448
rect 47362 -26512 47382 -26448
rect 41083 -26528 47382 -26512
rect 41083 -26592 47298 -26528
rect 47362 -26592 47382 -26528
rect 41083 -26608 47382 -26592
rect 41083 -26672 47298 -26608
rect 47362 -26672 47382 -26608
rect 41083 -26688 47382 -26672
rect 41083 -26752 47298 -26688
rect 47362 -26752 47382 -26688
rect 41083 -26768 47382 -26752
rect 41083 -26832 47298 -26768
rect 47362 -26832 47382 -26768
rect 41083 -26848 47382 -26832
rect 41083 -26912 47298 -26848
rect 47362 -26912 47382 -26848
rect 41083 -26928 47382 -26912
rect 41083 -26992 47298 -26928
rect 47362 -26992 47382 -26928
rect 41083 -27008 47382 -26992
rect 41083 -27072 47298 -27008
rect 47362 -27072 47382 -27008
rect 41083 -27088 47382 -27072
rect 41083 -27152 47298 -27088
rect 47362 -27152 47382 -27088
rect 41083 -27168 47382 -27152
rect 41083 -27232 47298 -27168
rect 47362 -27232 47382 -27168
rect 41083 -27248 47382 -27232
rect 41083 -27312 47298 -27248
rect 47362 -27312 47382 -27248
rect 41083 -27328 47382 -27312
rect 41083 -27392 47298 -27328
rect 47362 -27392 47382 -27328
rect 41083 -27408 47382 -27392
rect 41083 -27472 47298 -27408
rect 47362 -27472 47382 -27408
rect 41083 -27488 47382 -27472
rect 41083 -27552 47298 -27488
rect 47362 -27552 47382 -27488
rect 41083 -27568 47382 -27552
rect 41083 -27632 47298 -27568
rect 47362 -27632 47382 -27568
rect 41083 -27648 47382 -27632
rect 41083 -27712 47298 -27648
rect 47362 -27712 47382 -27648
rect 41083 -27728 47382 -27712
rect 41083 -27792 47298 -27728
rect 47362 -27792 47382 -27728
rect 41083 -27808 47382 -27792
rect 41083 -27872 47298 -27808
rect 47362 -27872 47382 -27808
rect 41083 -27888 47382 -27872
rect 41083 -27952 47298 -27888
rect 47362 -27952 47382 -27888
rect 41083 -27968 47382 -27952
rect 41083 -28032 47298 -27968
rect 47362 -28032 47382 -27968
rect 41083 -28048 47382 -28032
rect 41083 -28112 47298 -28048
rect 47362 -28112 47382 -28048
rect 41083 -28128 47382 -28112
rect 41083 -28192 47298 -28128
rect 47362 -28192 47382 -28128
rect 41083 -28208 47382 -28192
rect 41083 -28272 47298 -28208
rect 47362 -28272 47382 -28208
rect 41083 -28300 47382 -28272
rect -47383 -28428 -41084 -28400
rect -47383 -28492 -41168 -28428
rect -41104 -28492 -41084 -28428
rect -47383 -28508 -41084 -28492
rect -47383 -28572 -41168 -28508
rect -41104 -28572 -41084 -28508
rect -47383 -28588 -41084 -28572
rect -47383 -28652 -41168 -28588
rect -41104 -28652 -41084 -28588
rect -47383 -28668 -41084 -28652
rect -47383 -28732 -41168 -28668
rect -41104 -28732 -41084 -28668
rect -47383 -28748 -41084 -28732
rect -47383 -28812 -41168 -28748
rect -41104 -28812 -41084 -28748
rect -47383 -28828 -41084 -28812
rect -47383 -28892 -41168 -28828
rect -41104 -28892 -41084 -28828
rect -47383 -28908 -41084 -28892
rect -47383 -28972 -41168 -28908
rect -41104 -28972 -41084 -28908
rect -47383 -28988 -41084 -28972
rect -47383 -29052 -41168 -28988
rect -41104 -29052 -41084 -28988
rect -47383 -29068 -41084 -29052
rect -47383 -29132 -41168 -29068
rect -41104 -29132 -41084 -29068
rect -47383 -29148 -41084 -29132
rect -47383 -29212 -41168 -29148
rect -41104 -29212 -41084 -29148
rect -47383 -29228 -41084 -29212
rect -47383 -29292 -41168 -29228
rect -41104 -29292 -41084 -29228
rect -47383 -29308 -41084 -29292
rect -47383 -29372 -41168 -29308
rect -41104 -29372 -41084 -29308
rect -47383 -29388 -41084 -29372
rect -47383 -29452 -41168 -29388
rect -41104 -29452 -41084 -29388
rect -47383 -29468 -41084 -29452
rect -47383 -29532 -41168 -29468
rect -41104 -29532 -41084 -29468
rect -47383 -29548 -41084 -29532
rect -47383 -29612 -41168 -29548
rect -41104 -29612 -41084 -29548
rect -47383 -29628 -41084 -29612
rect -47383 -29692 -41168 -29628
rect -41104 -29692 -41084 -29628
rect -47383 -29708 -41084 -29692
rect -47383 -29772 -41168 -29708
rect -41104 -29772 -41084 -29708
rect -47383 -29788 -41084 -29772
rect -47383 -29852 -41168 -29788
rect -41104 -29852 -41084 -29788
rect -47383 -29868 -41084 -29852
rect -47383 -29932 -41168 -29868
rect -41104 -29932 -41084 -29868
rect -47383 -29948 -41084 -29932
rect -47383 -30012 -41168 -29948
rect -41104 -30012 -41084 -29948
rect -47383 -30028 -41084 -30012
rect -47383 -30092 -41168 -30028
rect -41104 -30092 -41084 -30028
rect -47383 -30108 -41084 -30092
rect -47383 -30172 -41168 -30108
rect -41104 -30172 -41084 -30108
rect -47383 -30188 -41084 -30172
rect -47383 -30252 -41168 -30188
rect -41104 -30252 -41084 -30188
rect -47383 -30268 -41084 -30252
rect -47383 -30332 -41168 -30268
rect -41104 -30332 -41084 -30268
rect -47383 -30348 -41084 -30332
rect -47383 -30412 -41168 -30348
rect -41104 -30412 -41084 -30348
rect -47383 -30428 -41084 -30412
rect -47383 -30492 -41168 -30428
rect -41104 -30492 -41084 -30428
rect -47383 -30508 -41084 -30492
rect -47383 -30572 -41168 -30508
rect -41104 -30572 -41084 -30508
rect -47383 -30588 -41084 -30572
rect -47383 -30652 -41168 -30588
rect -41104 -30652 -41084 -30588
rect -47383 -30668 -41084 -30652
rect -47383 -30732 -41168 -30668
rect -41104 -30732 -41084 -30668
rect -47383 -30748 -41084 -30732
rect -47383 -30812 -41168 -30748
rect -41104 -30812 -41084 -30748
rect -47383 -30828 -41084 -30812
rect -47383 -30892 -41168 -30828
rect -41104 -30892 -41084 -30828
rect -47383 -30908 -41084 -30892
rect -47383 -30972 -41168 -30908
rect -41104 -30972 -41084 -30908
rect -47383 -30988 -41084 -30972
rect -47383 -31052 -41168 -30988
rect -41104 -31052 -41084 -30988
rect -47383 -31068 -41084 -31052
rect -47383 -31132 -41168 -31068
rect -41104 -31132 -41084 -31068
rect -47383 -31148 -41084 -31132
rect -47383 -31212 -41168 -31148
rect -41104 -31212 -41084 -31148
rect -47383 -31228 -41084 -31212
rect -47383 -31292 -41168 -31228
rect -41104 -31292 -41084 -31228
rect -47383 -31308 -41084 -31292
rect -47383 -31372 -41168 -31308
rect -41104 -31372 -41084 -31308
rect -47383 -31388 -41084 -31372
rect -47383 -31452 -41168 -31388
rect -41104 -31452 -41084 -31388
rect -47383 -31468 -41084 -31452
rect -47383 -31532 -41168 -31468
rect -41104 -31532 -41084 -31468
rect -47383 -31548 -41084 -31532
rect -47383 -31612 -41168 -31548
rect -41104 -31612 -41084 -31548
rect -47383 -31628 -41084 -31612
rect -47383 -31692 -41168 -31628
rect -41104 -31692 -41084 -31628
rect -47383 -31708 -41084 -31692
rect -47383 -31772 -41168 -31708
rect -41104 -31772 -41084 -31708
rect -47383 -31788 -41084 -31772
rect -47383 -31852 -41168 -31788
rect -41104 -31852 -41084 -31788
rect -47383 -31868 -41084 -31852
rect -47383 -31932 -41168 -31868
rect -41104 -31932 -41084 -31868
rect -47383 -31948 -41084 -31932
rect -47383 -32012 -41168 -31948
rect -41104 -32012 -41084 -31948
rect -47383 -32028 -41084 -32012
rect -47383 -32092 -41168 -32028
rect -41104 -32092 -41084 -32028
rect -47383 -32108 -41084 -32092
rect -47383 -32172 -41168 -32108
rect -41104 -32172 -41084 -32108
rect -47383 -32188 -41084 -32172
rect -47383 -32252 -41168 -32188
rect -41104 -32252 -41084 -32188
rect -47383 -32268 -41084 -32252
rect -47383 -32332 -41168 -32268
rect -41104 -32332 -41084 -32268
rect -47383 -32348 -41084 -32332
rect -47383 -32412 -41168 -32348
rect -41104 -32412 -41084 -32348
rect -47383 -32428 -41084 -32412
rect -47383 -32492 -41168 -32428
rect -41104 -32492 -41084 -32428
rect -47383 -32508 -41084 -32492
rect -47383 -32572 -41168 -32508
rect -41104 -32572 -41084 -32508
rect -47383 -32588 -41084 -32572
rect -47383 -32652 -41168 -32588
rect -41104 -32652 -41084 -32588
rect -47383 -32668 -41084 -32652
rect -47383 -32732 -41168 -32668
rect -41104 -32732 -41084 -32668
rect -47383 -32748 -41084 -32732
rect -47383 -32812 -41168 -32748
rect -41104 -32812 -41084 -32748
rect -47383 -32828 -41084 -32812
rect -47383 -32892 -41168 -32828
rect -41104 -32892 -41084 -32828
rect -47383 -32908 -41084 -32892
rect -47383 -32972 -41168 -32908
rect -41104 -32972 -41084 -32908
rect -47383 -32988 -41084 -32972
rect -47383 -33052 -41168 -32988
rect -41104 -33052 -41084 -32988
rect -47383 -33068 -41084 -33052
rect -47383 -33132 -41168 -33068
rect -41104 -33132 -41084 -33068
rect -47383 -33148 -41084 -33132
rect -47383 -33212 -41168 -33148
rect -41104 -33212 -41084 -33148
rect -47383 -33228 -41084 -33212
rect -47383 -33292 -41168 -33228
rect -41104 -33292 -41084 -33228
rect -47383 -33308 -41084 -33292
rect -47383 -33372 -41168 -33308
rect -41104 -33372 -41084 -33308
rect -47383 -33388 -41084 -33372
rect -47383 -33452 -41168 -33388
rect -41104 -33452 -41084 -33388
rect -47383 -33468 -41084 -33452
rect -47383 -33532 -41168 -33468
rect -41104 -33532 -41084 -33468
rect -47383 -33548 -41084 -33532
rect -47383 -33612 -41168 -33548
rect -41104 -33612 -41084 -33548
rect -47383 -33628 -41084 -33612
rect -47383 -33692 -41168 -33628
rect -41104 -33692 -41084 -33628
rect -47383 -33708 -41084 -33692
rect -47383 -33772 -41168 -33708
rect -41104 -33772 -41084 -33708
rect -47383 -33788 -41084 -33772
rect -47383 -33852 -41168 -33788
rect -41104 -33852 -41084 -33788
rect -47383 -33868 -41084 -33852
rect -47383 -33932 -41168 -33868
rect -41104 -33932 -41084 -33868
rect -47383 -33948 -41084 -33932
rect -47383 -34012 -41168 -33948
rect -41104 -34012 -41084 -33948
rect -47383 -34028 -41084 -34012
rect -47383 -34092 -41168 -34028
rect -41104 -34092 -41084 -34028
rect -47383 -34108 -41084 -34092
rect -47383 -34172 -41168 -34108
rect -41104 -34172 -41084 -34108
rect -47383 -34188 -41084 -34172
rect -47383 -34252 -41168 -34188
rect -41104 -34252 -41084 -34188
rect -47383 -34268 -41084 -34252
rect -47383 -34332 -41168 -34268
rect -41104 -34332 -41084 -34268
rect -47383 -34348 -41084 -34332
rect -47383 -34412 -41168 -34348
rect -41104 -34412 -41084 -34348
rect -47383 -34428 -41084 -34412
rect -47383 -34492 -41168 -34428
rect -41104 -34492 -41084 -34428
rect -47383 -34508 -41084 -34492
rect -47383 -34572 -41168 -34508
rect -41104 -34572 -41084 -34508
rect -47383 -34600 -41084 -34572
rect -41064 -28428 -34765 -28400
rect -41064 -28492 -34849 -28428
rect -34785 -28492 -34765 -28428
rect -41064 -28508 -34765 -28492
rect -41064 -28572 -34849 -28508
rect -34785 -28572 -34765 -28508
rect -41064 -28588 -34765 -28572
rect -41064 -28652 -34849 -28588
rect -34785 -28652 -34765 -28588
rect -41064 -28668 -34765 -28652
rect -41064 -28732 -34849 -28668
rect -34785 -28732 -34765 -28668
rect -41064 -28748 -34765 -28732
rect -41064 -28812 -34849 -28748
rect -34785 -28812 -34765 -28748
rect -41064 -28828 -34765 -28812
rect -41064 -28892 -34849 -28828
rect -34785 -28892 -34765 -28828
rect -41064 -28908 -34765 -28892
rect -41064 -28972 -34849 -28908
rect -34785 -28972 -34765 -28908
rect -41064 -28988 -34765 -28972
rect -41064 -29052 -34849 -28988
rect -34785 -29052 -34765 -28988
rect -41064 -29068 -34765 -29052
rect -41064 -29132 -34849 -29068
rect -34785 -29132 -34765 -29068
rect -41064 -29148 -34765 -29132
rect -41064 -29212 -34849 -29148
rect -34785 -29212 -34765 -29148
rect -41064 -29228 -34765 -29212
rect -41064 -29292 -34849 -29228
rect -34785 -29292 -34765 -29228
rect -41064 -29308 -34765 -29292
rect -41064 -29372 -34849 -29308
rect -34785 -29372 -34765 -29308
rect -41064 -29388 -34765 -29372
rect -41064 -29452 -34849 -29388
rect -34785 -29452 -34765 -29388
rect -41064 -29468 -34765 -29452
rect -41064 -29532 -34849 -29468
rect -34785 -29532 -34765 -29468
rect -41064 -29548 -34765 -29532
rect -41064 -29612 -34849 -29548
rect -34785 -29612 -34765 -29548
rect -41064 -29628 -34765 -29612
rect -41064 -29692 -34849 -29628
rect -34785 -29692 -34765 -29628
rect -41064 -29708 -34765 -29692
rect -41064 -29772 -34849 -29708
rect -34785 -29772 -34765 -29708
rect -41064 -29788 -34765 -29772
rect -41064 -29852 -34849 -29788
rect -34785 -29852 -34765 -29788
rect -41064 -29868 -34765 -29852
rect -41064 -29932 -34849 -29868
rect -34785 -29932 -34765 -29868
rect -41064 -29948 -34765 -29932
rect -41064 -30012 -34849 -29948
rect -34785 -30012 -34765 -29948
rect -41064 -30028 -34765 -30012
rect -41064 -30092 -34849 -30028
rect -34785 -30092 -34765 -30028
rect -41064 -30108 -34765 -30092
rect -41064 -30172 -34849 -30108
rect -34785 -30172 -34765 -30108
rect -41064 -30188 -34765 -30172
rect -41064 -30252 -34849 -30188
rect -34785 -30252 -34765 -30188
rect -41064 -30268 -34765 -30252
rect -41064 -30332 -34849 -30268
rect -34785 -30332 -34765 -30268
rect -41064 -30348 -34765 -30332
rect -41064 -30412 -34849 -30348
rect -34785 -30412 -34765 -30348
rect -41064 -30428 -34765 -30412
rect -41064 -30492 -34849 -30428
rect -34785 -30492 -34765 -30428
rect -41064 -30508 -34765 -30492
rect -41064 -30572 -34849 -30508
rect -34785 -30572 -34765 -30508
rect -41064 -30588 -34765 -30572
rect -41064 -30652 -34849 -30588
rect -34785 -30652 -34765 -30588
rect -41064 -30668 -34765 -30652
rect -41064 -30732 -34849 -30668
rect -34785 -30732 -34765 -30668
rect -41064 -30748 -34765 -30732
rect -41064 -30812 -34849 -30748
rect -34785 -30812 -34765 -30748
rect -41064 -30828 -34765 -30812
rect -41064 -30892 -34849 -30828
rect -34785 -30892 -34765 -30828
rect -41064 -30908 -34765 -30892
rect -41064 -30972 -34849 -30908
rect -34785 -30972 -34765 -30908
rect -41064 -30988 -34765 -30972
rect -41064 -31052 -34849 -30988
rect -34785 -31052 -34765 -30988
rect -41064 -31068 -34765 -31052
rect -41064 -31132 -34849 -31068
rect -34785 -31132 -34765 -31068
rect -41064 -31148 -34765 -31132
rect -41064 -31212 -34849 -31148
rect -34785 -31212 -34765 -31148
rect -41064 -31228 -34765 -31212
rect -41064 -31292 -34849 -31228
rect -34785 -31292 -34765 -31228
rect -41064 -31308 -34765 -31292
rect -41064 -31372 -34849 -31308
rect -34785 -31372 -34765 -31308
rect -41064 -31388 -34765 -31372
rect -41064 -31452 -34849 -31388
rect -34785 -31452 -34765 -31388
rect -41064 -31468 -34765 -31452
rect -41064 -31532 -34849 -31468
rect -34785 -31532 -34765 -31468
rect -41064 -31548 -34765 -31532
rect -41064 -31612 -34849 -31548
rect -34785 -31612 -34765 -31548
rect -41064 -31628 -34765 -31612
rect -41064 -31692 -34849 -31628
rect -34785 -31692 -34765 -31628
rect -41064 -31708 -34765 -31692
rect -41064 -31772 -34849 -31708
rect -34785 -31772 -34765 -31708
rect -41064 -31788 -34765 -31772
rect -41064 -31852 -34849 -31788
rect -34785 -31852 -34765 -31788
rect -41064 -31868 -34765 -31852
rect -41064 -31932 -34849 -31868
rect -34785 -31932 -34765 -31868
rect -41064 -31948 -34765 -31932
rect -41064 -32012 -34849 -31948
rect -34785 -32012 -34765 -31948
rect -41064 -32028 -34765 -32012
rect -41064 -32092 -34849 -32028
rect -34785 -32092 -34765 -32028
rect -41064 -32108 -34765 -32092
rect -41064 -32172 -34849 -32108
rect -34785 -32172 -34765 -32108
rect -41064 -32188 -34765 -32172
rect -41064 -32252 -34849 -32188
rect -34785 -32252 -34765 -32188
rect -41064 -32268 -34765 -32252
rect -41064 -32332 -34849 -32268
rect -34785 -32332 -34765 -32268
rect -41064 -32348 -34765 -32332
rect -41064 -32412 -34849 -32348
rect -34785 -32412 -34765 -32348
rect -41064 -32428 -34765 -32412
rect -41064 -32492 -34849 -32428
rect -34785 -32492 -34765 -32428
rect -41064 -32508 -34765 -32492
rect -41064 -32572 -34849 -32508
rect -34785 -32572 -34765 -32508
rect -41064 -32588 -34765 -32572
rect -41064 -32652 -34849 -32588
rect -34785 -32652 -34765 -32588
rect -41064 -32668 -34765 -32652
rect -41064 -32732 -34849 -32668
rect -34785 -32732 -34765 -32668
rect -41064 -32748 -34765 -32732
rect -41064 -32812 -34849 -32748
rect -34785 -32812 -34765 -32748
rect -41064 -32828 -34765 -32812
rect -41064 -32892 -34849 -32828
rect -34785 -32892 -34765 -32828
rect -41064 -32908 -34765 -32892
rect -41064 -32972 -34849 -32908
rect -34785 -32972 -34765 -32908
rect -41064 -32988 -34765 -32972
rect -41064 -33052 -34849 -32988
rect -34785 -33052 -34765 -32988
rect -41064 -33068 -34765 -33052
rect -41064 -33132 -34849 -33068
rect -34785 -33132 -34765 -33068
rect -41064 -33148 -34765 -33132
rect -41064 -33212 -34849 -33148
rect -34785 -33212 -34765 -33148
rect -41064 -33228 -34765 -33212
rect -41064 -33292 -34849 -33228
rect -34785 -33292 -34765 -33228
rect -41064 -33308 -34765 -33292
rect -41064 -33372 -34849 -33308
rect -34785 -33372 -34765 -33308
rect -41064 -33388 -34765 -33372
rect -41064 -33452 -34849 -33388
rect -34785 -33452 -34765 -33388
rect -41064 -33468 -34765 -33452
rect -41064 -33532 -34849 -33468
rect -34785 -33532 -34765 -33468
rect -41064 -33548 -34765 -33532
rect -41064 -33612 -34849 -33548
rect -34785 -33612 -34765 -33548
rect -41064 -33628 -34765 -33612
rect -41064 -33692 -34849 -33628
rect -34785 -33692 -34765 -33628
rect -41064 -33708 -34765 -33692
rect -41064 -33772 -34849 -33708
rect -34785 -33772 -34765 -33708
rect -41064 -33788 -34765 -33772
rect -41064 -33852 -34849 -33788
rect -34785 -33852 -34765 -33788
rect -41064 -33868 -34765 -33852
rect -41064 -33932 -34849 -33868
rect -34785 -33932 -34765 -33868
rect -41064 -33948 -34765 -33932
rect -41064 -34012 -34849 -33948
rect -34785 -34012 -34765 -33948
rect -41064 -34028 -34765 -34012
rect -41064 -34092 -34849 -34028
rect -34785 -34092 -34765 -34028
rect -41064 -34108 -34765 -34092
rect -41064 -34172 -34849 -34108
rect -34785 -34172 -34765 -34108
rect -41064 -34188 -34765 -34172
rect -41064 -34252 -34849 -34188
rect -34785 -34252 -34765 -34188
rect -41064 -34268 -34765 -34252
rect -41064 -34332 -34849 -34268
rect -34785 -34332 -34765 -34268
rect -41064 -34348 -34765 -34332
rect -41064 -34412 -34849 -34348
rect -34785 -34412 -34765 -34348
rect -41064 -34428 -34765 -34412
rect -41064 -34492 -34849 -34428
rect -34785 -34492 -34765 -34428
rect -41064 -34508 -34765 -34492
rect -41064 -34572 -34849 -34508
rect -34785 -34572 -34765 -34508
rect -41064 -34600 -34765 -34572
rect -34745 -28428 -28446 -28400
rect -34745 -28492 -28530 -28428
rect -28466 -28492 -28446 -28428
rect -34745 -28508 -28446 -28492
rect -34745 -28572 -28530 -28508
rect -28466 -28572 -28446 -28508
rect -34745 -28588 -28446 -28572
rect -34745 -28652 -28530 -28588
rect -28466 -28652 -28446 -28588
rect -34745 -28668 -28446 -28652
rect -34745 -28732 -28530 -28668
rect -28466 -28732 -28446 -28668
rect -34745 -28748 -28446 -28732
rect -34745 -28812 -28530 -28748
rect -28466 -28812 -28446 -28748
rect -34745 -28828 -28446 -28812
rect -34745 -28892 -28530 -28828
rect -28466 -28892 -28446 -28828
rect -34745 -28908 -28446 -28892
rect -34745 -28972 -28530 -28908
rect -28466 -28972 -28446 -28908
rect -34745 -28988 -28446 -28972
rect -34745 -29052 -28530 -28988
rect -28466 -29052 -28446 -28988
rect -34745 -29068 -28446 -29052
rect -34745 -29132 -28530 -29068
rect -28466 -29132 -28446 -29068
rect -34745 -29148 -28446 -29132
rect -34745 -29212 -28530 -29148
rect -28466 -29212 -28446 -29148
rect -34745 -29228 -28446 -29212
rect -34745 -29292 -28530 -29228
rect -28466 -29292 -28446 -29228
rect -34745 -29308 -28446 -29292
rect -34745 -29372 -28530 -29308
rect -28466 -29372 -28446 -29308
rect -34745 -29388 -28446 -29372
rect -34745 -29452 -28530 -29388
rect -28466 -29452 -28446 -29388
rect -34745 -29468 -28446 -29452
rect -34745 -29532 -28530 -29468
rect -28466 -29532 -28446 -29468
rect -34745 -29548 -28446 -29532
rect -34745 -29612 -28530 -29548
rect -28466 -29612 -28446 -29548
rect -34745 -29628 -28446 -29612
rect -34745 -29692 -28530 -29628
rect -28466 -29692 -28446 -29628
rect -34745 -29708 -28446 -29692
rect -34745 -29772 -28530 -29708
rect -28466 -29772 -28446 -29708
rect -34745 -29788 -28446 -29772
rect -34745 -29852 -28530 -29788
rect -28466 -29852 -28446 -29788
rect -34745 -29868 -28446 -29852
rect -34745 -29932 -28530 -29868
rect -28466 -29932 -28446 -29868
rect -34745 -29948 -28446 -29932
rect -34745 -30012 -28530 -29948
rect -28466 -30012 -28446 -29948
rect -34745 -30028 -28446 -30012
rect -34745 -30092 -28530 -30028
rect -28466 -30092 -28446 -30028
rect -34745 -30108 -28446 -30092
rect -34745 -30172 -28530 -30108
rect -28466 -30172 -28446 -30108
rect -34745 -30188 -28446 -30172
rect -34745 -30252 -28530 -30188
rect -28466 -30252 -28446 -30188
rect -34745 -30268 -28446 -30252
rect -34745 -30332 -28530 -30268
rect -28466 -30332 -28446 -30268
rect -34745 -30348 -28446 -30332
rect -34745 -30412 -28530 -30348
rect -28466 -30412 -28446 -30348
rect -34745 -30428 -28446 -30412
rect -34745 -30492 -28530 -30428
rect -28466 -30492 -28446 -30428
rect -34745 -30508 -28446 -30492
rect -34745 -30572 -28530 -30508
rect -28466 -30572 -28446 -30508
rect -34745 -30588 -28446 -30572
rect -34745 -30652 -28530 -30588
rect -28466 -30652 -28446 -30588
rect -34745 -30668 -28446 -30652
rect -34745 -30732 -28530 -30668
rect -28466 -30732 -28446 -30668
rect -34745 -30748 -28446 -30732
rect -34745 -30812 -28530 -30748
rect -28466 -30812 -28446 -30748
rect -34745 -30828 -28446 -30812
rect -34745 -30892 -28530 -30828
rect -28466 -30892 -28446 -30828
rect -34745 -30908 -28446 -30892
rect -34745 -30972 -28530 -30908
rect -28466 -30972 -28446 -30908
rect -34745 -30988 -28446 -30972
rect -34745 -31052 -28530 -30988
rect -28466 -31052 -28446 -30988
rect -34745 -31068 -28446 -31052
rect -34745 -31132 -28530 -31068
rect -28466 -31132 -28446 -31068
rect -34745 -31148 -28446 -31132
rect -34745 -31212 -28530 -31148
rect -28466 -31212 -28446 -31148
rect -34745 -31228 -28446 -31212
rect -34745 -31292 -28530 -31228
rect -28466 -31292 -28446 -31228
rect -34745 -31308 -28446 -31292
rect -34745 -31372 -28530 -31308
rect -28466 -31372 -28446 -31308
rect -34745 -31388 -28446 -31372
rect -34745 -31452 -28530 -31388
rect -28466 -31452 -28446 -31388
rect -34745 -31468 -28446 -31452
rect -34745 -31532 -28530 -31468
rect -28466 -31532 -28446 -31468
rect -34745 -31548 -28446 -31532
rect -34745 -31612 -28530 -31548
rect -28466 -31612 -28446 -31548
rect -34745 -31628 -28446 -31612
rect -34745 -31692 -28530 -31628
rect -28466 -31692 -28446 -31628
rect -34745 -31708 -28446 -31692
rect -34745 -31772 -28530 -31708
rect -28466 -31772 -28446 -31708
rect -34745 -31788 -28446 -31772
rect -34745 -31852 -28530 -31788
rect -28466 -31852 -28446 -31788
rect -34745 -31868 -28446 -31852
rect -34745 -31932 -28530 -31868
rect -28466 -31932 -28446 -31868
rect -34745 -31948 -28446 -31932
rect -34745 -32012 -28530 -31948
rect -28466 -32012 -28446 -31948
rect -34745 -32028 -28446 -32012
rect -34745 -32092 -28530 -32028
rect -28466 -32092 -28446 -32028
rect -34745 -32108 -28446 -32092
rect -34745 -32172 -28530 -32108
rect -28466 -32172 -28446 -32108
rect -34745 -32188 -28446 -32172
rect -34745 -32252 -28530 -32188
rect -28466 -32252 -28446 -32188
rect -34745 -32268 -28446 -32252
rect -34745 -32332 -28530 -32268
rect -28466 -32332 -28446 -32268
rect -34745 -32348 -28446 -32332
rect -34745 -32412 -28530 -32348
rect -28466 -32412 -28446 -32348
rect -34745 -32428 -28446 -32412
rect -34745 -32492 -28530 -32428
rect -28466 -32492 -28446 -32428
rect -34745 -32508 -28446 -32492
rect -34745 -32572 -28530 -32508
rect -28466 -32572 -28446 -32508
rect -34745 -32588 -28446 -32572
rect -34745 -32652 -28530 -32588
rect -28466 -32652 -28446 -32588
rect -34745 -32668 -28446 -32652
rect -34745 -32732 -28530 -32668
rect -28466 -32732 -28446 -32668
rect -34745 -32748 -28446 -32732
rect -34745 -32812 -28530 -32748
rect -28466 -32812 -28446 -32748
rect -34745 -32828 -28446 -32812
rect -34745 -32892 -28530 -32828
rect -28466 -32892 -28446 -32828
rect -34745 -32908 -28446 -32892
rect -34745 -32972 -28530 -32908
rect -28466 -32972 -28446 -32908
rect -34745 -32988 -28446 -32972
rect -34745 -33052 -28530 -32988
rect -28466 -33052 -28446 -32988
rect -34745 -33068 -28446 -33052
rect -34745 -33132 -28530 -33068
rect -28466 -33132 -28446 -33068
rect -34745 -33148 -28446 -33132
rect -34745 -33212 -28530 -33148
rect -28466 -33212 -28446 -33148
rect -34745 -33228 -28446 -33212
rect -34745 -33292 -28530 -33228
rect -28466 -33292 -28446 -33228
rect -34745 -33308 -28446 -33292
rect -34745 -33372 -28530 -33308
rect -28466 -33372 -28446 -33308
rect -34745 -33388 -28446 -33372
rect -34745 -33452 -28530 -33388
rect -28466 -33452 -28446 -33388
rect -34745 -33468 -28446 -33452
rect -34745 -33532 -28530 -33468
rect -28466 -33532 -28446 -33468
rect -34745 -33548 -28446 -33532
rect -34745 -33612 -28530 -33548
rect -28466 -33612 -28446 -33548
rect -34745 -33628 -28446 -33612
rect -34745 -33692 -28530 -33628
rect -28466 -33692 -28446 -33628
rect -34745 -33708 -28446 -33692
rect -34745 -33772 -28530 -33708
rect -28466 -33772 -28446 -33708
rect -34745 -33788 -28446 -33772
rect -34745 -33852 -28530 -33788
rect -28466 -33852 -28446 -33788
rect -34745 -33868 -28446 -33852
rect -34745 -33932 -28530 -33868
rect -28466 -33932 -28446 -33868
rect -34745 -33948 -28446 -33932
rect -34745 -34012 -28530 -33948
rect -28466 -34012 -28446 -33948
rect -34745 -34028 -28446 -34012
rect -34745 -34092 -28530 -34028
rect -28466 -34092 -28446 -34028
rect -34745 -34108 -28446 -34092
rect -34745 -34172 -28530 -34108
rect -28466 -34172 -28446 -34108
rect -34745 -34188 -28446 -34172
rect -34745 -34252 -28530 -34188
rect -28466 -34252 -28446 -34188
rect -34745 -34268 -28446 -34252
rect -34745 -34332 -28530 -34268
rect -28466 -34332 -28446 -34268
rect -34745 -34348 -28446 -34332
rect -34745 -34412 -28530 -34348
rect -28466 -34412 -28446 -34348
rect -34745 -34428 -28446 -34412
rect -34745 -34492 -28530 -34428
rect -28466 -34492 -28446 -34428
rect -34745 -34508 -28446 -34492
rect -34745 -34572 -28530 -34508
rect -28466 -34572 -28446 -34508
rect -34745 -34600 -28446 -34572
rect -28426 -28428 -22127 -28400
rect -28426 -28492 -22211 -28428
rect -22147 -28492 -22127 -28428
rect -28426 -28508 -22127 -28492
rect -28426 -28572 -22211 -28508
rect -22147 -28572 -22127 -28508
rect -28426 -28588 -22127 -28572
rect -28426 -28652 -22211 -28588
rect -22147 -28652 -22127 -28588
rect -28426 -28668 -22127 -28652
rect -28426 -28732 -22211 -28668
rect -22147 -28732 -22127 -28668
rect -28426 -28748 -22127 -28732
rect -28426 -28812 -22211 -28748
rect -22147 -28812 -22127 -28748
rect -28426 -28828 -22127 -28812
rect -28426 -28892 -22211 -28828
rect -22147 -28892 -22127 -28828
rect -28426 -28908 -22127 -28892
rect -28426 -28972 -22211 -28908
rect -22147 -28972 -22127 -28908
rect -28426 -28988 -22127 -28972
rect -28426 -29052 -22211 -28988
rect -22147 -29052 -22127 -28988
rect -28426 -29068 -22127 -29052
rect -28426 -29132 -22211 -29068
rect -22147 -29132 -22127 -29068
rect -28426 -29148 -22127 -29132
rect -28426 -29212 -22211 -29148
rect -22147 -29212 -22127 -29148
rect -28426 -29228 -22127 -29212
rect -28426 -29292 -22211 -29228
rect -22147 -29292 -22127 -29228
rect -28426 -29308 -22127 -29292
rect -28426 -29372 -22211 -29308
rect -22147 -29372 -22127 -29308
rect -28426 -29388 -22127 -29372
rect -28426 -29452 -22211 -29388
rect -22147 -29452 -22127 -29388
rect -28426 -29468 -22127 -29452
rect -28426 -29532 -22211 -29468
rect -22147 -29532 -22127 -29468
rect -28426 -29548 -22127 -29532
rect -28426 -29612 -22211 -29548
rect -22147 -29612 -22127 -29548
rect -28426 -29628 -22127 -29612
rect -28426 -29692 -22211 -29628
rect -22147 -29692 -22127 -29628
rect -28426 -29708 -22127 -29692
rect -28426 -29772 -22211 -29708
rect -22147 -29772 -22127 -29708
rect -28426 -29788 -22127 -29772
rect -28426 -29852 -22211 -29788
rect -22147 -29852 -22127 -29788
rect -28426 -29868 -22127 -29852
rect -28426 -29932 -22211 -29868
rect -22147 -29932 -22127 -29868
rect -28426 -29948 -22127 -29932
rect -28426 -30012 -22211 -29948
rect -22147 -30012 -22127 -29948
rect -28426 -30028 -22127 -30012
rect -28426 -30092 -22211 -30028
rect -22147 -30092 -22127 -30028
rect -28426 -30108 -22127 -30092
rect -28426 -30172 -22211 -30108
rect -22147 -30172 -22127 -30108
rect -28426 -30188 -22127 -30172
rect -28426 -30252 -22211 -30188
rect -22147 -30252 -22127 -30188
rect -28426 -30268 -22127 -30252
rect -28426 -30332 -22211 -30268
rect -22147 -30332 -22127 -30268
rect -28426 -30348 -22127 -30332
rect -28426 -30412 -22211 -30348
rect -22147 -30412 -22127 -30348
rect -28426 -30428 -22127 -30412
rect -28426 -30492 -22211 -30428
rect -22147 -30492 -22127 -30428
rect -28426 -30508 -22127 -30492
rect -28426 -30572 -22211 -30508
rect -22147 -30572 -22127 -30508
rect -28426 -30588 -22127 -30572
rect -28426 -30652 -22211 -30588
rect -22147 -30652 -22127 -30588
rect -28426 -30668 -22127 -30652
rect -28426 -30732 -22211 -30668
rect -22147 -30732 -22127 -30668
rect -28426 -30748 -22127 -30732
rect -28426 -30812 -22211 -30748
rect -22147 -30812 -22127 -30748
rect -28426 -30828 -22127 -30812
rect -28426 -30892 -22211 -30828
rect -22147 -30892 -22127 -30828
rect -28426 -30908 -22127 -30892
rect -28426 -30972 -22211 -30908
rect -22147 -30972 -22127 -30908
rect -28426 -30988 -22127 -30972
rect -28426 -31052 -22211 -30988
rect -22147 -31052 -22127 -30988
rect -28426 -31068 -22127 -31052
rect -28426 -31132 -22211 -31068
rect -22147 -31132 -22127 -31068
rect -28426 -31148 -22127 -31132
rect -28426 -31212 -22211 -31148
rect -22147 -31212 -22127 -31148
rect -28426 -31228 -22127 -31212
rect -28426 -31292 -22211 -31228
rect -22147 -31292 -22127 -31228
rect -28426 -31308 -22127 -31292
rect -28426 -31372 -22211 -31308
rect -22147 -31372 -22127 -31308
rect -28426 -31388 -22127 -31372
rect -28426 -31452 -22211 -31388
rect -22147 -31452 -22127 -31388
rect -28426 -31468 -22127 -31452
rect -28426 -31532 -22211 -31468
rect -22147 -31532 -22127 -31468
rect -28426 -31548 -22127 -31532
rect -28426 -31612 -22211 -31548
rect -22147 -31612 -22127 -31548
rect -28426 -31628 -22127 -31612
rect -28426 -31692 -22211 -31628
rect -22147 -31692 -22127 -31628
rect -28426 -31708 -22127 -31692
rect -28426 -31772 -22211 -31708
rect -22147 -31772 -22127 -31708
rect -28426 -31788 -22127 -31772
rect -28426 -31852 -22211 -31788
rect -22147 -31852 -22127 -31788
rect -28426 -31868 -22127 -31852
rect -28426 -31932 -22211 -31868
rect -22147 -31932 -22127 -31868
rect -28426 -31948 -22127 -31932
rect -28426 -32012 -22211 -31948
rect -22147 -32012 -22127 -31948
rect -28426 -32028 -22127 -32012
rect -28426 -32092 -22211 -32028
rect -22147 -32092 -22127 -32028
rect -28426 -32108 -22127 -32092
rect -28426 -32172 -22211 -32108
rect -22147 -32172 -22127 -32108
rect -28426 -32188 -22127 -32172
rect -28426 -32252 -22211 -32188
rect -22147 -32252 -22127 -32188
rect -28426 -32268 -22127 -32252
rect -28426 -32332 -22211 -32268
rect -22147 -32332 -22127 -32268
rect -28426 -32348 -22127 -32332
rect -28426 -32412 -22211 -32348
rect -22147 -32412 -22127 -32348
rect -28426 -32428 -22127 -32412
rect -28426 -32492 -22211 -32428
rect -22147 -32492 -22127 -32428
rect -28426 -32508 -22127 -32492
rect -28426 -32572 -22211 -32508
rect -22147 -32572 -22127 -32508
rect -28426 -32588 -22127 -32572
rect -28426 -32652 -22211 -32588
rect -22147 -32652 -22127 -32588
rect -28426 -32668 -22127 -32652
rect -28426 -32732 -22211 -32668
rect -22147 -32732 -22127 -32668
rect -28426 -32748 -22127 -32732
rect -28426 -32812 -22211 -32748
rect -22147 -32812 -22127 -32748
rect -28426 -32828 -22127 -32812
rect -28426 -32892 -22211 -32828
rect -22147 -32892 -22127 -32828
rect -28426 -32908 -22127 -32892
rect -28426 -32972 -22211 -32908
rect -22147 -32972 -22127 -32908
rect -28426 -32988 -22127 -32972
rect -28426 -33052 -22211 -32988
rect -22147 -33052 -22127 -32988
rect -28426 -33068 -22127 -33052
rect -28426 -33132 -22211 -33068
rect -22147 -33132 -22127 -33068
rect -28426 -33148 -22127 -33132
rect -28426 -33212 -22211 -33148
rect -22147 -33212 -22127 -33148
rect -28426 -33228 -22127 -33212
rect -28426 -33292 -22211 -33228
rect -22147 -33292 -22127 -33228
rect -28426 -33308 -22127 -33292
rect -28426 -33372 -22211 -33308
rect -22147 -33372 -22127 -33308
rect -28426 -33388 -22127 -33372
rect -28426 -33452 -22211 -33388
rect -22147 -33452 -22127 -33388
rect -28426 -33468 -22127 -33452
rect -28426 -33532 -22211 -33468
rect -22147 -33532 -22127 -33468
rect -28426 -33548 -22127 -33532
rect -28426 -33612 -22211 -33548
rect -22147 -33612 -22127 -33548
rect -28426 -33628 -22127 -33612
rect -28426 -33692 -22211 -33628
rect -22147 -33692 -22127 -33628
rect -28426 -33708 -22127 -33692
rect -28426 -33772 -22211 -33708
rect -22147 -33772 -22127 -33708
rect -28426 -33788 -22127 -33772
rect -28426 -33852 -22211 -33788
rect -22147 -33852 -22127 -33788
rect -28426 -33868 -22127 -33852
rect -28426 -33932 -22211 -33868
rect -22147 -33932 -22127 -33868
rect -28426 -33948 -22127 -33932
rect -28426 -34012 -22211 -33948
rect -22147 -34012 -22127 -33948
rect -28426 -34028 -22127 -34012
rect -28426 -34092 -22211 -34028
rect -22147 -34092 -22127 -34028
rect -28426 -34108 -22127 -34092
rect -28426 -34172 -22211 -34108
rect -22147 -34172 -22127 -34108
rect -28426 -34188 -22127 -34172
rect -28426 -34252 -22211 -34188
rect -22147 -34252 -22127 -34188
rect -28426 -34268 -22127 -34252
rect -28426 -34332 -22211 -34268
rect -22147 -34332 -22127 -34268
rect -28426 -34348 -22127 -34332
rect -28426 -34412 -22211 -34348
rect -22147 -34412 -22127 -34348
rect -28426 -34428 -22127 -34412
rect -28426 -34492 -22211 -34428
rect -22147 -34492 -22127 -34428
rect -28426 -34508 -22127 -34492
rect -28426 -34572 -22211 -34508
rect -22147 -34572 -22127 -34508
rect -28426 -34600 -22127 -34572
rect -22107 -28428 -15808 -28400
rect -22107 -28492 -15892 -28428
rect -15828 -28492 -15808 -28428
rect -22107 -28508 -15808 -28492
rect -22107 -28572 -15892 -28508
rect -15828 -28572 -15808 -28508
rect -22107 -28588 -15808 -28572
rect -22107 -28652 -15892 -28588
rect -15828 -28652 -15808 -28588
rect -22107 -28668 -15808 -28652
rect -22107 -28732 -15892 -28668
rect -15828 -28732 -15808 -28668
rect -22107 -28748 -15808 -28732
rect -22107 -28812 -15892 -28748
rect -15828 -28812 -15808 -28748
rect -22107 -28828 -15808 -28812
rect -22107 -28892 -15892 -28828
rect -15828 -28892 -15808 -28828
rect -22107 -28908 -15808 -28892
rect -22107 -28972 -15892 -28908
rect -15828 -28972 -15808 -28908
rect -22107 -28988 -15808 -28972
rect -22107 -29052 -15892 -28988
rect -15828 -29052 -15808 -28988
rect -22107 -29068 -15808 -29052
rect -22107 -29132 -15892 -29068
rect -15828 -29132 -15808 -29068
rect -22107 -29148 -15808 -29132
rect -22107 -29212 -15892 -29148
rect -15828 -29212 -15808 -29148
rect -22107 -29228 -15808 -29212
rect -22107 -29292 -15892 -29228
rect -15828 -29292 -15808 -29228
rect -22107 -29308 -15808 -29292
rect -22107 -29372 -15892 -29308
rect -15828 -29372 -15808 -29308
rect -22107 -29388 -15808 -29372
rect -22107 -29452 -15892 -29388
rect -15828 -29452 -15808 -29388
rect -22107 -29468 -15808 -29452
rect -22107 -29532 -15892 -29468
rect -15828 -29532 -15808 -29468
rect -22107 -29548 -15808 -29532
rect -22107 -29612 -15892 -29548
rect -15828 -29612 -15808 -29548
rect -22107 -29628 -15808 -29612
rect -22107 -29692 -15892 -29628
rect -15828 -29692 -15808 -29628
rect -22107 -29708 -15808 -29692
rect -22107 -29772 -15892 -29708
rect -15828 -29772 -15808 -29708
rect -22107 -29788 -15808 -29772
rect -22107 -29852 -15892 -29788
rect -15828 -29852 -15808 -29788
rect -22107 -29868 -15808 -29852
rect -22107 -29932 -15892 -29868
rect -15828 -29932 -15808 -29868
rect -22107 -29948 -15808 -29932
rect -22107 -30012 -15892 -29948
rect -15828 -30012 -15808 -29948
rect -22107 -30028 -15808 -30012
rect -22107 -30092 -15892 -30028
rect -15828 -30092 -15808 -30028
rect -22107 -30108 -15808 -30092
rect -22107 -30172 -15892 -30108
rect -15828 -30172 -15808 -30108
rect -22107 -30188 -15808 -30172
rect -22107 -30252 -15892 -30188
rect -15828 -30252 -15808 -30188
rect -22107 -30268 -15808 -30252
rect -22107 -30332 -15892 -30268
rect -15828 -30332 -15808 -30268
rect -22107 -30348 -15808 -30332
rect -22107 -30412 -15892 -30348
rect -15828 -30412 -15808 -30348
rect -22107 -30428 -15808 -30412
rect -22107 -30492 -15892 -30428
rect -15828 -30492 -15808 -30428
rect -22107 -30508 -15808 -30492
rect -22107 -30572 -15892 -30508
rect -15828 -30572 -15808 -30508
rect -22107 -30588 -15808 -30572
rect -22107 -30652 -15892 -30588
rect -15828 -30652 -15808 -30588
rect -22107 -30668 -15808 -30652
rect -22107 -30732 -15892 -30668
rect -15828 -30732 -15808 -30668
rect -22107 -30748 -15808 -30732
rect -22107 -30812 -15892 -30748
rect -15828 -30812 -15808 -30748
rect -22107 -30828 -15808 -30812
rect -22107 -30892 -15892 -30828
rect -15828 -30892 -15808 -30828
rect -22107 -30908 -15808 -30892
rect -22107 -30972 -15892 -30908
rect -15828 -30972 -15808 -30908
rect -22107 -30988 -15808 -30972
rect -22107 -31052 -15892 -30988
rect -15828 -31052 -15808 -30988
rect -22107 -31068 -15808 -31052
rect -22107 -31132 -15892 -31068
rect -15828 -31132 -15808 -31068
rect -22107 -31148 -15808 -31132
rect -22107 -31212 -15892 -31148
rect -15828 -31212 -15808 -31148
rect -22107 -31228 -15808 -31212
rect -22107 -31292 -15892 -31228
rect -15828 -31292 -15808 -31228
rect -22107 -31308 -15808 -31292
rect -22107 -31372 -15892 -31308
rect -15828 -31372 -15808 -31308
rect -22107 -31388 -15808 -31372
rect -22107 -31452 -15892 -31388
rect -15828 -31452 -15808 -31388
rect -22107 -31468 -15808 -31452
rect -22107 -31532 -15892 -31468
rect -15828 -31532 -15808 -31468
rect -22107 -31548 -15808 -31532
rect -22107 -31612 -15892 -31548
rect -15828 -31612 -15808 -31548
rect -22107 -31628 -15808 -31612
rect -22107 -31692 -15892 -31628
rect -15828 -31692 -15808 -31628
rect -22107 -31708 -15808 -31692
rect -22107 -31772 -15892 -31708
rect -15828 -31772 -15808 -31708
rect -22107 -31788 -15808 -31772
rect -22107 -31852 -15892 -31788
rect -15828 -31852 -15808 -31788
rect -22107 -31868 -15808 -31852
rect -22107 -31932 -15892 -31868
rect -15828 -31932 -15808 -31868
rect -22107 -31948 -15808 -31932
rect -22107 -32012 -15892 -31948
rect -15828 -32012 -15808 -31948
rect -22107 -32028 -15808 -32012
rect -22107 -32092 -15892 -32028
rect -15828 -32092 -15808 -32028
rect -22107 -32108 -15808 -32092
rect -22107 -32172 -15892 -32108
rect -15828 -32172 -15808 -32108
rect -22107 -32188 -15808 -32172
rect -22107 -32252 -15892 -32188
rect -15828 -32252 -15808 -32188
rect -22107 -32268 -15808 -32252
rect -22107 -32332 -15892 -32268
rect -15828 -32332 -15808 -32268
rect -22107 -32348 -15808 -32332
rect -22107 -32412 -15892 -32348
rect -15828 -32412 -15808 -32348
rect -22107 -32428 -15808 -32412
rect -22107 -32492 -15892 -32428
rect -15828 -32492 -15808 -32428
rect -22107 -32508 -15808 -32492
rect -22107 -32572 -15892 -32508
rect -15828 -32572 -15808 -32508
rect -22107 -32588 -15808 -32572
rect -22107 -32652 -15892 -32588
rect -15828 -32652 -15808 -32588
rect -22107 -32668 -15808 -32652
rect -22107 -32732 -15892 -32668
rect -15828 -32732 -15808 -32668
rect -22107 -32748 -15808 -32732
rect -22107 -32812 -15892 -32748
rect -15828 -32812 -15808 -32748
rect -22107 -32828 -15808 -32812
rect -22107 -32892 -15892 -32828
rect -15828 -32892 -15808 -32828
rect -22107 -32908 -15808 -32892
rect -22107 -32972 -15892 -32908
rect -15828 -32972 -15808 -32908
rect -22107 -32988 -15808 -32972
rect -22107 -33052 -15892 -32988
rect -15828 -33052 -15808 -32988
rect -22107 -33068 -15808 -33052
rect -22107 -33132 -15892 -33068
rect -15828 -33132 -15808 -33068
rect -22107 -33148 -15808 -33132
rect -22107 -33212 -15892 -33148
rect -15828 -33212 -15808 -33148
rect -22107 -33228 -15808 -33212
rect -22107 -33292 -15892 -33228
rect -15828 -33292 -15808 -33228
rect -22107 -33308 -15808 -33292
rect -22107 -33372 -15892 -33308
rect -15828 -33372 -15808 -33308
rect -22107 -33388 -15808 -33372
rect -22107 -33452 -15892 -33388
rect -15828 -33452 -15808 -33388
rect -22107 -33468 -15808 -33452
rect -22107 -33532 -15892 -33468
rect -15828 -33532 -15808 -33468
rect -22107 -33548 -15808 -33532
rect -22107 -33612 -15892 -33548
rect -15828 -33612 -15808 -33548
rect -22107 -33628 -15808 -33612
rect -22107 -33692 -15892 -33628
rect -15828 -33692 -15808 -33628
rect -22107 -33708 -15808 -33692
rect -22107 -33772 -15892 -33708
rect -15828 -33772 -15808 -33708
rect -22107 -33788 -15808 -33772
rect -22107 -33852 -15892 -33788
rect -15828 -33852 -15808 -33788
rect -22107 -33868 -15808 -33852
rect -22107 -33932 -15892 -33868
rect -15828 -33932 -15808 -33868
rect -22107 -33948 -15808 -33932
rect -22107 -34012 -15892 -33948
rect -15828 -34012 -15808 -33948
rect -22107 -34028 -15808 -34012
rect -22107 -34092 -15892 -34028
rect -15828 -34092 -15808 -34028
rect -22107 -34108 -15808 -34092
rect -22107 -34172 -15892 -34108
rect -15828 -34172 -15808 -34108
rect -22107 -34188 -15808 -34172
rect -22107 -34252 -15892 -34188
rect -15828 -34252 -15808 -34188
rect -22107 -34268 -15808 -34252
rect -22107 -34332 -15892 -34268
rect -15828 -34332 -15808 -34268
rect -22107 -34348 -15808 -34332
rect -22107 -34412 -15892 -34348
rect -15828 -34412 -15808 -34348
rect -22107 -34428 -15808 -34412
rect -22107 -34492 -15892 -34428
rect -15828 -34492 -15808 -34428
rect -22107 -34508 -15808 -34492
rect -22107 -34572 -15892 -34508
rect -15828 -34572 -15808 -34508
rect -22107 -34600 -15808 -34572
rect -15788 -28428 -9489 -28400
rect -15788 -28492 -9573 -28428
rect -9509 -28492 -9489 -28428
rect -15788 -28508 -9489 -28492
rect -15788 -28572 -9573 -28508
rect -9509 -28572 -9489 -28508
rect -15788 -28588 -9489 -28572
rect -15788 -28652 -9573 -28588
rect -9509 -28652 -9489 -28588
rect -15788 -28668 -9489 -28652
rect -15788 -28732 -9573 -28668
rect -9509 -28732 -9489 -28668
rect -15788 -28748 -9489 -28732
rect -15788 -28812 -9573 -28748
rect -9509 -28812 -9489 -28748
rect -15788 -28828 -9489 -28812
rect -15788 -28892 -9573 -28828
rect -9509 -28892 -9489 -28828
rect -15788 -28908 -9489 -28892
rect -15788 -28972 -9573 -28908
rect -9509 -28972 -9489 -28908
rect -15788 -28988 -9489 -28972
rect -15788 -29052 -9573 -28988
rect -9509 -29052 -9489 -28988
rect -15788 -29068 -9489 -29052
rect -15788 -29132 -9573 -29068
rect -9509 -29132 -9489 -29068
rect -15788 -29148 -9489 -29132
rect -15788 -29212 -9573 -29148
rect -9509 -29212 -9489 -29148
rect -15788 -29228 -9489 -29212
rect -15788 -29292 -9573 -29228
rect -9509 -29292 -9489 -29228
rect -15788 -29308 -9489 -29292
rect -15788 -29372 -9573 -29308
rect -9509 -29372 -9489 -29308
rect -15788 -29388 -9489 -29372
rect -15788 -29452 -9573 -29388
rect -9509 -29452 -9489 -29388
rect -15788 -29468 -9489 -29452
rect -15788 -29532 -9573 -29468
rect -9509 -29532 -9489 -29468
rect -15788 -29548 -9489 -29532
rect -15788 -29612 -9573 -29548
rect -9509 -29612 -9489 -29548
rect -15788 -29628 -9489 -29612
rect -15788 -29692 -9573 -29628
rect -9509 -29692 -9489 -29628
rect -15788 -29708 -9489 -29692
rect -15788 -29772 -9573 -29708
rect -9509 -29772 -9489 -29708
rect -15788 -29788 -9489 -29772
rect -15788 -29852 -9573 -29788
rect -9509 -29852 -9489 -29788
rect -15788 -29868 -9489 -29852
rect -15788 -29932 -9573 -29868
rect -9509 -29932 -9489 -29868
rect -15788 -29948 -9489 -29932
rect -15788 -30012 -9573 -29948
rect -9509 -30012 -9489 -29948
rect -15788 -30028 -9489 -30012
rect -15788 -30092 -9573 -30028
rect -9509 -30092 -9489 -30028
rect -15788 -30108 -9489 -30092
rect -15788 -30172 -9573 -30108
rect -9509 -30172 -9489 -30108
rect -15788 -30188 -9489 -30172
rect -15788 -30252 -9573 -30188
rect -9509 -30252 -9489 -30188
rect -15788 -30268 -9489 -30252
rect -15788 -30332 -9573 -30268
rect -9509 -30332 -9489 -30268
rect -15788 -30348 -9489 -30332
rect -15788 -30412 -9573 -30348
rect -9509 -30412 -9489 -30348
rect -15788 -30428 -9489 -30412
rect -15788 -30492 -9573 -30428
rect -9509 -30492 -9489 -30428
rect -15788 -30508 -9489 -30492
rect -15788 -30572 -9573 -30508
rect -9509 -30572 -9489 -30508
rect -15788 -30588 -9489 -30572
rect -15788 -30652 -9573 -30588
rect -9509 -30652 -9489 -30588
rect -15788 -30668 -9489 -30652
rect -15788 -30732 -9573 -30668
rect -9509 -30732 -9489 -30668
rect -15788 -30748 -9489 -30732
rect -15788 -30812 -9573 -30748
rect -9509 -30812 -9489 -30748
rect -15788 -30828 -9489 -30812
rect -15788 -30892 -9573 -30828
rect -9509 -30892 -9489 -30828
rect -15788 -30908 -9489 -30892
rect -15788 -30972 -9573 -30908
rect -9509 -30972 -9489 -30908
rect -15788 -30988 -9489 -30972
rect -15788 -31052 -9573 -30988
rect -9509 -31052 -9489 -30988
rect -15788 -31068 -9489 -31052
rect -15788 -31132 -9573 -31068
rect -9509 -31132 -9489 -31068
rect -15788 -31148 -9489 -31132
rect -15788 -31212 -9573 -31148
rect -9509 -31212 -9489 -31148
rect -15788 -31228 -9489 -31212
rect -15788 -31292 -9573 -31228
rect -9509 -31292 -9489 -31228
rect -15788 -31308 -9489 -31292
rect -15788 -31372 -9573 -31308
rect -9509 -31372 -9489 -31308
rect -15788 -31388 -9489 -31372
rect -15788 -31452 -9573 -31388
rect -9509 -31452 -9489 -31388
rect -15788 -31468 -9489 -31452
rect -15788 -31532 -9573 -31468
rect -9509 -31532 -9489 -31468
rect -15788 -31548 -9489 -31532
rect -15788 -31612 -9573 -31548
rect -9509 -31612 -9489 -31548
rect -15788 -31628 -9489 -31612
rect -15788 -31692 -9573 -31628
rect -9509 -31692 -9489 -31628
rect -15788 -31708 -9489 -31692
rect -15788 -31772 -9573 -31708
rect -9509 -31772 -9489 -31708
rect -15788 -31788 -9489 -31772
rect -15788 -31852 -9573 -31788
rect -9509 -31852 -9489 -31788
rect -15788 -31868 -9489 -31852
rect -15788 -31932 -9573 -31868
rect -9509 -31932 -9489 -31868
rect -15788 -31948 -9489 -31932
rect -15788 -32012 -9573 -31948
rect -9509 -32012 -9489 -31948
rect -15788 -32028 -9489 -32012
rect -15788 -32092 -9573 -32028
rect -9509 -32092 -9489 -32028
rect -15788 -32108 -9489 -32092
rect -15788 -32172 -9573 -32108
rect -9509 -32172 -9489 -32108
rect -15788 -32188 -9489 -32172
rect -15788 -32252 -9573 -32188
rect -9509 -32252 -9489 -32188
rect -15788 -32268 -9489 -32252
rect -15788 -32332 -9573 -32268
rect -9509 -32332 -9489 -32268
rect -15788 -32348 -9489 -32332
rect -15788 -32412 -9573 -32348
rect -9509 -32412 -9489 -32348
rect -15788 -32428 -9489 -32412
rect -15788 -32492 -9573 -32428
rect -9509 -32492 -9489 -32428
rect -15788 -32508 -9489 -32492
rect -15788 -32572 -9573 -32508
rect -9509 -32572 -9489 -32508
rect -15788 -32588 -9489 -32572
rect -15788 -32652 -9573 -32588
rect -9509 -32652 -9489 -32588
rect -15788 -32668 -9489 -32652
rect -15788 -32732 -9573 -32668
rect -9509 -32732 -9489 -32668
rect -15788 -32748 -9489 -32732
rect -15788 -32812 -9573 -32748
rect -9509 -32812 -9489 -32748
rect -15788 -32828 -9489 -32812
rect -15788 -32892 -9573 -32828
rect -9509 -32892 -9489 -32828
rect -15788 -32908 -9489 -32892
rect -15788 -32972 -9573 -32908
rect -9509 -32972 -9489 -32908
rect -15788 -32988 -9489 -32972
rect -15788 -33052 -9573 -32988
rect -9509 -33052 -9489 -32988
rect -15788 -33068 -9489 -33052
rect -15788 -33132 -9573 -33068
rect -9509 -33132 -9489 -33068
rect -15788 -33148 -9489 -33132
rect -15788 -33212 -9573 -33148
rect -9509 -33212 -9489 -33148
rect -15788 -33228 -9489 -33212
rect -15788 -33292 -9573 -33228
rect -9509 -33292 -9489 -33228
rect -15788 -33308 -9489 -33292
rect -15788 -33372 -9573 -33308
rect -9509 -33372 -9489 -33308
rect -15788 -33388 -9489 -33372
rect -15788 -33452 -9573 -33388
rect -9509 -33452 -9489 -33388
rect -15788 -33468 -9489 -33452
rect -15788 -33532 -9573 -33468
rect -9509 -33532 -9489 -33468
rect -15788 -33548 -9489 -33532
rect -15788 -33612 -9573 -33548
rect -9509 -33612 -9489 -33548
rect -15788 -33628 -9489 -33612
rect -15788 -33692 -9573 -33628
rect -9509 -33692 -9489 -33628
rect -15788 -33708 -9489 -33692
rect -15788 -33772 -9573 -33708
rect -9509 -33772 -9489 -33708
rect -15788 -33788 -9489 -33772
rect -15788 -33852 -9573 -33788
rect -9509 -33852 -9489 -33788
rect -15788 -33868 -9489 -33852
rect -15788 -33932 -9573 -33868
rect -9509 -33932 -9489 -33868
rect -15788 -33948 -9489 -33932
rect -15788 -34012 -9573 -33948
rect -9509 -34012 -9489 -33948
rect -15788 -34028 -9489 -34012
rect -15788 -34092 -9573 -34028
rect -9509 -34092 -9489 -34028
rect -15788 -34108 -9489 -34092
rect -15788 -34172 -9573 -34108
rect -9509 -34172 -9489 -34108
rect -15788 -34188 -9489 -34172
rect -15788 -34252 -9573 -34188
rect -9509 -34252 -9489 -34188
rect -15788 -34268 -9489 -34252
rect -15788 -34332 -9573 -34268
rect -9509 -34332 -9489 -34268
rect -15788 -34348 -9489 -34332
rect -15788 -34412 -9573 -34348
rect -9509 -34412 -9489 -34348
rect -15788 -34428 -9489 -34412
rect -15788 -34492 -9573 -34428
rect -9509 -34492 -9489 -34428
rect -15788 -34508 -9489 -34492
rect -15788 -34572 -9573 -34508
rect -9509 -34572 -9489 -34508
rect -15788 -34600 -9489 -34572
rect -9469 -28428 -3170 -28400
rect -9469 -28492 -3254 -28428
rect -3190 -28492 -3170 -28428
rect -9469 -28508 -3170 -28492
rect -9469 -28572 -3254 -28508
rect -3190 -28572 -3170 -28508
rect -9469 -28588 -3170 -28572
rect -9469 -28652 -3254 -28588
rect -3190 -28652 -3170 -28588
rect -9469 -28668 -3170 -28652
rect -9469 -28732 -3254 -28668
rect -3190 -28732 -3170 -28668
rect -9469 -28748 -3170 -28732
rect -9469 -28812 -3254 -28748
rect -3190 -28812 -3170 -28748
rect -9469 -28828 -3170 -28812
rect -9469 -28892 -3254 -28828
rect -3190 -28892 -3170 -28828
rect -9469 -28908 -3170 -28892
rect -9469 -28972 -3254 -28908
rect -3190 -28972 -3170 -28908
rect -9469 -28988 -3170 -28972
rect -9469 -29052 -3254 -28988
rect -3190 -29052 -3170 -28988
rect -9469 -29068 -3170 -29052
rect -9469 -29132 -3254 -29068
rect -3190 -29132 -3170 -29068
rect -9469 -29148 -3170 -29132
rect -9469 -29212 -3254 -29148
rect -3190 -29212 -3170 -29148
rect -9469 -29228 -3170 -29212
rect -9469 -29292 -3254 -29228
rect -3190 -29292 -3170 -29228
rect -9469 -29308 -3170 -29292
rect -9469 -29372 -3254 -29308
rect -3190 -29372 -3170 -29308
rect -9469 -29388 -3170 -29372
rect -9469 -29452 -3254 -29388
rect -3190 -29452 -3170 -29388
rect -9469 -29468 -3170 -29452
rect -9469 -29532 -3254 -29468
rect -3190 -29532 -3170 -29468
rect -9469 -29548 -3170 -29532
rect -9469 -29612 -3254 -29548
rect -3190 -29612 -3170 -29548
rect -9469 -29628 -3170 -29612
rect -9469 -29692 -3254 -29628
rect -3190 -29692 -3170 -29628
rect -9469 -29708 -3170 -29692
rect -9469 -29772 -3254 -29708
rect -3190 -29772 -3170 -29708
rect -9469 -29788 -3170 -29772
rect -9469 -29852 -3254 -29788
rect -3190 -29852 -3170 -29788
rect -9469 -29868 -3170 -29852
rect -9469 -29932 -3254 -29868
rect -3190 -29932 -3170 -29868
rect -9469 -29948 -3170 -29932
rect -9469 -30012 -3254 -29948
rect -3190 -30012 -3170 -29948
rect -9469 -30028 -3170 -30012
rect -9469 -30092 -3254 -30028
rect -3190 -30092 -3170 -30028
rect -9469 -30108 -3170 -30092
rect -9469 -30172 -3254 -30108
rect -3190 -30172 -3170 -30108
rect -9469 -30188 -3170 -30172
rect -9469 -30252 -3254 -30188
rect -3190 -30252 -3170 -30188
rect -9469 -30268 -3170 -30252
rect -9469 -30332 -3254 -30268
rect -3190 -30332 -3170 -30268
rect -9469 -30348 -3170 -30332
rect -9469 -30412 -3254 -30348
rect -3190 -30412 -3170 -30348
rect -9469 -30428 -3170 -30412
rect -9469 -30492 -3254 -30428
rect -3190 -30492 -3170 -30428
rect -9469 -30508 -3170 -30492
rect -9469 -30572 -3254 -30508
rect -3190 -30572 -3170 -30508
rect -9469 -30588 -3170 -30572
rect -9469 -30652 -3254 -30588
rect -3190 -30652 -3170 -30588
rect -9469 -30668 -3170 -30652
rect -9469 -30732 -3254 -30668
rect -3190 -30732 -3170 -30668
rect -9469 -30748 -3170 -30732
rect -9469 -30812 -3254 -30748
rect -3190 -30812 -3170 -30748
rect -9469 -30828 -3170 -30812
rect -9469 -30892 -3254 -30828
rect -3190 -30892 -3170 -30828
rect -9469 -30908 -3170 -30892
rect -9469 -30972 -3254 -30908
rect -3190 -30972 -3170 -30908
rect -9469 -30988 -3170 -30972
rect -9469 -31052 -3254 -30988
rect -3190 -31052 -3170 -30988
rect -9469 -31068 -3170 -31052
rect -9469 -31132 -3254 -31068
rect -3190 -31132 -3170 -31068
rect -9469 -31148 -3170 -31132
rect -9469 -31212 -3254 -31148
rect -3190 -31212 -3170 -31148
rect -9469 -31228 -3170 -31212
rect -9469 -31292 -3254 -31228
rect -3190 -31292 -3170 -31228
rect -9469 -31308 -3170 -31292
rect -9469 -31372 -3254 -31308
rect -3190 -31372 -3170 -31308
rect -9469 -31388 -3170 -31372
rect -9469 -31452 -3254 -31388
rect -3190 -31452 -3170 -31388
rect -9469 -31468 -3170 -31452
rect -9469 -31532 -3254 -31468
rect -3190 -31532 -3170 -31468
rect -9469 -31548 -3170 -31532
rect -9469 -31612 -3254 -31548
rect -3190 -31612 -3170 -31548
rect -9469 -31628 -3170 -31612
rect -9469 -31692 -3254 -31628
rect -3190 -31692 -3170 -31628
rect -9469 -31708 -3170 -31692
rect -9469 -31772 -3254 -31708
rect -3190 -31772 -3170 -31708
rect -9469 -31788 -3170 -31772
rect -9469 -31852 -3254 -31788
rect -3190 -31852 -3170 -31788
rect -9469 -31868 -3170 -31852
rect -9469 -31932 -3254 -31868
rect -3190 -31932 -3170 -31868
rect -9469 -31948 -3170 -31932
rect -9469 -32012 -3254 -31948
rect -3190 -32012 -3170 -31948
rect -9469 -32028 -3170 -32012
rect -9469 -32092 -3254 -32028
rect -3190 -32092 -3170 -32028
rect -9469 -32108 -3170 -32092
rect -9469 -32172 -3254 -32108
rect -3190 -32172 -3170 -32108
rect -9469 -32188 -3170 -32172
rect -9469 -32252 -3254 -32188
rect -3190 -32252 -3170 -32188
rect -9469 -32268 -3170 -32252
rect -9469 -32332 -3254 -32268
rect -3190 -32332 -3170 -32268
rect -9469 -32348 -3170 -32332
rect -9469 -32412 -3254 -32348
rect -3190 -32412 -3170 -32348
rect -9469 -32428 -3170 -32412
rect -9469 -32492 -3254 -32428
rect -3190 -32492 -3170 -32428
rect -9469 -32508 -3170 -32492
rect -9469 -32572 -3254 -32508
rect -3190 -32572 -3170 -32508
rect -9469 -32588 -3170 -32572
rect -9469 -32652 -3254 -32588
rect -3190 -32652 -3170 -32588
rect -9469 -32668 -3170 -32652
rect -9469 -32732 -3254 -32668
rect -3190 -32732 -3170 -32668
rect -9469 -32748 -3170 -32732
rect -9469 -32812 -3254 -32748
rect -3190 -32812 -3170 -32748
rect -9469 -32828 -3170 -32812
rect -9469 -32892 -3254 -32828
rect -3190 -32892 -3170 -32828
rect -9469 -32908 -3170 -32892
rect -9469 -32972 -3254 -32908
rect -3190 -32972 -3170 -32908
rect -9469 -32988 -3170 -32972
rect -9469 -33052 -3254 -32988
rect -3190 -33052 -3170 -32988
rect -9469 -33068 -3170 -33052
rect -9469 -33132 -3254 -33068
rect -3190 -33132 -3170 -33068
rect -9469 -33148 -3170 -33132
rect -9469 -33212 -3254 -33148
rect -3190 -33212 -3170 -33148
rect -9469 -33228 -3170 -33212
rect -9469 -33292 -3254 -33228
rect -3190 -33292 -3170 -33228
rect -9469 -33308 -3170 -33292
rect -9469 -33372 -3254 -33308
rect -3190 -33372 -3170 -33308
rect -9469 -33388 -3170 -33372
rect -9469 -33452 -3254 -33388
rect -3190 -33452 -3170 -33388
rect -9469 -33468 -3170 -33452
rect -9469 -33532 -3254 -33468
rect -3190 -33532 -3170 -33468
rect -9469 -33548 -3170 -33532
rect -9469 -33612 -3254 -33548
rect -3190 -33612 -3170 -33548
rect -9469 -33628 -3170 -33612
rect -9469 -33692 -3254 -33628
rect -3190 -33692 -3170 -33628
rect -9469 -33708 -3170 -33692
rect -9469 -33772 -3254 -33708
rect -3190 -33772 -3170 -33708
rect -9469 -33788 -3170 -33772
rect -9469 -33852 -3254 -33788
rect -3190 -33852 -3170 -33788
rect -9469 -33868 -3170 -33852
rect -9469 -33932 -3254 -33868
rect -3190 -33932 -3170 -33868
rect -9469 -33948 -3170 -33932
rect -9469 -34012 -3254 -33948
rect -3190 -34012 -3170 -33948
rect -9469 -34028 -3170 -34012
rect -9469 -34092 -3254 -34028
rect -3190 -34092 -3170 -34028
rect -9469 -34108 -3170 -34092
rect -9469 -34172 -3254 -34108
rect -3190 -34172 -3170 -34108
rect -9469 -34188 -3170 -34172
rect -9469 -34252 -3254 -34188
rect -3190 -34252 -3170 -34188
rect -9469 -34268 -3170 -34252
rect -9469 -34332 -3254 -34268
rect -3190 -34332 -3170 -34268
rect -9469 -34348 -3170 -34332
rect -9469 -34412 -3254 -34348
rect -3190 -34412 -3170 -34348
rect -9469 -34428 -3170 -34412
rect -9469 -34492 -3254 -34428
rect -3190 -34492 -3170 -34428
rect -9469 -34508 -3170 -34492
rect -9469 -34572 -3254 -34508
rect -3190 -34572 -3170 -34508
rect -9469 -34600 -3170 -34572
rect -3150 -28428 3149 -28400
rect -3150 -28492 3065 -28428
rect 3129 -28492 3149 -28428
rect -3150 -28508 3149 -28492
rect -3150 -28572 3065 -28508
rect 3129 -28572 3149 -28508
rect -3150 -28588 3149 -28572
rect -3150 -28652 3065 -28588
rect 3129 -28652 3149 -28588
rect -3150 -28668 3149 -28652
rect -3150 -28732 3065 -28668
rect 3129 -28732 3149 -28668
rect -3150 -28748 3149 -28732
rect -3150 -28812 3065 -28748
rect 3129 -28812 3149 -28748
rect -3150 -28828 3149 -28812
rect -3150 -28892 3065 -28828
rect 3129 -28892 3149 -28828
rect -3150 -28908 3149 -28892
rect -3150 -28972 3065 -28908
rect 3129 -28972 3149 -28908
rect -3150 -28988 3149 -28972
rect -3150 -29052 3065 -28988
rect 3129 -29052 3149 -28988
rect -3150 -29068 3149 -29052
rect -3150 -29132 3065 -29068
rect 3129 -29132 3149 -29068
rect -3150 -29148 3149 -29132
rect -3150 -29212 3065 -29148
rect 3129 -29212 3149 -29148
rect -3150 -29228 3149 -29212
rect -3150 -29292 3065 -29228
rect 3129 -29292 3149 -29228
rect -3150 -29308 3149 -29292
rect -3150 -29372 3065 -29308
rect 3129 -29372 3149 -29308
rect -3150 -29388 3149 -29372
rect -3150 -29452 3065 -29388
rect 3129 -29452 3149 -29388
rect -3150 -29468 3149 -29452
rect -3150 -29532 3065 -29468
rect 3129 -29532 3149 -29468
rect -3150 -29548 3149 -29532
rect -3150 -29612 3065 -29548
rect 3129 -29612 3149 -29548
rect -3150 -29628 3149 -29612
rect -3150 -29692 3065 -29628
rect 3129 -29692 3149 -29628
rect -3150 -29708 3149 -29692
rect -3150 -29772 3065 -29708
rect 3129 -29772 3149 -29708
rect -3150 -29788 3149 -29772
rect -3150 -29852 3065 -29788
rect 3129 -29852 3149 -29788
rect -3150 -29868 3149 -29852
rect -3150 -29932 3065 -29868
rect 3129 -29932 3149 -29868
rect -3150 -29948 3149 -29932
rect -3150 -30012 3065 -29948
rect 3129 -30012 3149 -29948
rect -3150 -30028 3149 -30012
rect -3150 -30092 3065 -30028
rect 3129 -30092 3149 -30028
rect -3150 -30108 3149 -30092
rect -3150 -30172 3065 -30108
rect 3129 -30172 3149 -30108
rect -3150 -30188 3149 -30172
rect -3150 -30252 3065 -30188
rect 3129 -30252 3149 -30188
rect -3150 -30268 3149 -30252
rect -3150 -30332 3065 -30268
rect 3129 -30332 3149 -30268
rect -3150 -30348 3149 -30332
rect -3150 -30412 3065 -30348
rect 3129 -30412 3149 -30348
rect -3150 -30428 3149 -30412
rect -3150 -30492 3065 -30428
rect 3129 -30492 3149 -30428
rect -3150 -30508 3149 -30492
rect -3150 -30572 3065 -30508
rect 3129 -30572 3149 -30508
rect -3150 -30588 3149 -30572
rect -3150 -30652 3065 -30588
rect 3129 -30652 3149 -30588
rect -3150 -30668 3149 -30652
rect -3150 -30732 3065 -30668
rect 3129 -30732 3149 -30668
rect -3150 -30748 3149 -30732
rect -3150 -30812 3065 -30748
rect 3129 -30812 3149 -30748
rect -3150 -30828 3149 -30812
rect -3150 -30892 3065 -30828
rect 3129 -30892 3149 -30828
rect -3150 -30908 3149 -30892
rect -3150 -30972 3065 -30908
rect 3129 -30972 3149 -30908
rect -3150 -30988 3149 -30972
rect -3150 -31052 3065 -30988
rect 3129 -31052 3149 -30988
rect -3150 -31068 3149 -31052
rect -3150 -31132 3065 -31068
rect 3129 -31132 3149 -31068
rect -3150 -31148 3149 -31132
rect -3150 -31212 3065 -31148
rect 3129 -31212 3149 -31148
rect -3150 -31228 3149 -31212
rect -3150 -31292 3065 -31228
rect 3129 -31292 3149 -31228
rect -3150 -31308 3149 -31292
rect -3150 -31372 3065 -31308
rect 3129 -31372 3149 -31308
rect -3150 -31388 3149 -31372
rect -3150 -31452 3065 -31388
rect 3129 -31452 3149 -31388
rect -3150 -31468 3149 -31452
rect -3150 -31532 3065 -31468
rect 3129 -31532 3149 -31468
rect -3150 -31548 3149 -31532
rect -3150 -31612 3065 -31548
rect 3129 -31612 3149 -31548
rect -3150 -31628 3149 -31612
rect -3150 -31692 3065 -31628
rect 3129 -31692 3149 -31628
rect -3150 -31708 3149 -31692
rect -3150 -31772 3065 -31708
rect 3129 -31772 3149 -31708
rect -3150 -31788 3149 -31772
rect -3150 -31852 3065 -31788
rect 3129 -31852 3149 -31788
rect -3150 -31868 3149 -31852
rect -3150 -31932 3065 -31868
rect 3129 -31932 3149 -31868
rect -3150 -31948 3149 -31932
rect -3150 -32012 3065 -31948
rect 3129 -32012 3149 -31948
rect -3150 -32028 3149 -32012
rect -3150 -32092 3065 -32028
rect 3129 -32092 3149 -32028
rect -3150 -32108 3149 -32092
rect -3150 -32172 3065 -32108
rect 3129 -32172 3149 -32108
rect -3150 -32188 3149 -32172
rect -3150 -32252 3065 -32188
rect 3129 -32252 3149 -32188
rect -3150 -32268 3149 -32252
rect -3150 -32332 3065 -32268
rect 3129 -32332 3149 -32268
rect -3150 -32348 3149 -32332
rect -3150 -32412 3065 -32348
rect 3129 -32412 3149 -32348
rect -3150 -32428 3149 -32412
rect -3150 -32492 3065 -32428
rect 3129 -32492 3149 -32428
rect -3150 -32508 3149 -32492
rect -3150 -32572 3065 -32508
rect 3129 -32572 3149 -32508
rect -3150 -32588 3149 -32572
rect -3150 -32652 3065 -32588
rect 3129 -32652 3149 -32588
rect -3150 -32668 3149 -32652
rect -3150 -32732 3065 -32668
rect 3129 -32732 3149 -32668
rect -3150 -32748 3149 -32732
rect -3150 -32812 3065 -32748
rect 3129 -32812 3149 -32748
rect -3150 -32828 3149 -32812
rect -3150 -32892 3065 -32828
rect 3129 -32892 3149 -32828
rect -3150 -32908 3149 -32892
rect -3150 -32972 3065 -32908
rect 3129 -32972 3149 -32908
rect -3150 -32988 3149 -32972
rect -3150 -33052 3065 -32988
rect 3129 -33052 3149 -32988
rect -3150 -33068 3149 -33052
rect -3150 -33132 3065 -33068
rect 3129 -33132 3149 -33068
rect -3150 -33148 3149 -33132
rect -3150 -33212 3065 -33148
rect 3129 -33212 3149 -33148
rect -3150 -33228 3149 -33212
rect -3150 -33292 3065 -33228
rect 3129 -33292 3149 -33228
rect -3150 -33308 3149 -33292
rect -3150 -33372 3065 -33308
rect 3129 -33372 3149 -33308
rect -3150 -33388 3149 -33372
rect -3150 -33452 3065 -33388
rect 3129 -33452 3149 -33388
rect -3150 -33468 3149 -33452
rect -3150 -33532 3065 -33468
rect 3129 -33532 3149 -33468
rect -3150 -33548 3149 -33532
rect -3150 -33612 3065 -33548
rect 3129 -33612 3149 -33548
rect -3150 -33628 3149 -33612
rect -3150 -33692 3065 -33628
rect 3129 -33692 3149 -33628
rect -3150 -33708 3149 -33692
rect -3150 -33772 3065 -33708
rect 3129 -33772 3149 -33708
rect -3150 -33788 3149 -33772
rect -3150 -33852 3065 -33788
rect 3129 -33852 3149 -33788
rect -3150 -33868 3149 -33852
rect -3150 -33932 3065 -33868
rect 3129 -33932 3149 -33868
rect -3150 -33948 3149 -33932
rect -3150 -34012 3065 -33948
rect 3129 -34012 3149 -33948
rect -3150 -34028 3149 -34012
rect -3150 -34092 3065 -34028
rect 3129 -34092 3149 -34028
rect -3150 -34108 3149 -34092
rect -3150 -34172 3065 -34108
rect 3129 -34172 3149 -34108
rect -3150 -34188 3149 -34172
rect -3150 -34252 3065 -34188
rect 3129 -34252 3149 -34188
rect -3150 -34268 3149 -34252
rect -3150 -34332 3065 -34268
rect 3129 -34332 3149 -34268
rect -3150 -34348 3149 -34332
rect -3150 -34412 3065 -34348
rect 3129 -34412 3149 -34348
rect -3150 -34428 3149 -34412
rect -3150 -34492 3065 -34428
rect 3129 -34492 3149 -34428
rect -3150 -34508 3149 -34492
rect -3150 -34572 3065 -34508
rect 3129 -34572 3149 -34508
rect -3150 -34600 3149 -34572
rect 3169 -28428 9468 -28400
rect 3169 -28492 9384 -28428
rect 9448 -28492 9468 -28428
rect 3169 -28508 9468 -28492
rect 3169 -28572 9384 -28508
rect 9448 -28572 9468 -28508
rect 3169 -28588 9468 -28572
rect 3169 -28652 9384 -28588
rect 9448 -28652 9468 -28588
rect 3169 -28668 9468 -28652
rect 3169 -28732 9384 -28668
rect 9448 -28732 9468 -28668
rect 3169 -28748 9468 -28732
rect 3169 -28812 9384 -28748
rect 9448 -28812 9468 -28748
rect 3169 -28828 9468 -28812
rect 3169 -28892 9384 -28828
rect 9448 -28892 9468 -28828
rect 3169 -28908 9468 -28892
rect 3169 -28972 9384 -28908
rect 9448 -28972 9468 -28908
rect 3169 -28988 9468 -28972
rect 3169 -29052 9384 -28988
rect 9448 -29052 9468 -28988
rect 3169 -29068 9468 -29052
rect 3169 -29132 9384 -29068
rect 9448 -29132 9468 -29068
rect 3169 -29148 9468 -29132
rect 3169 -29212 9384 -29148
rect 9448 -29212 9468 -29148
rect 3169 -29228 9468 -29212
rect 3169 -29292 9384 -29228
rect 9448 -29292 9468 -29228
rect 3169 -29308 9468 -29292
rect 3169 -29372 9384 -29308
rect 9448 -29372 9468 -29308
rect 3169 -29388 9468 -29372
rect 3169 -29452 9384 -29388
rect 9448 -29452 9468 -29388
rect 3169 -29468 9468 -29452
rect 3169 -29532 9384 -29468
rect 9448 -29532 9468 -29468
rect 3169 -29548 9468 -29532
rect 3169 -29612 9384 -29548
rect 9448 -29612 9468 -29548
rect 3169 -29628 9468 -29612
rect 3169 -29692 9384 -29628
rect 9448 -29692 9468 -29628
rect 3169 -29708 9468 -29692
rect 3169 -29772 9384 -29708
rect 9448 -29772 9468 -29708
rect 3169 -29788 9468 -29772
rect 3169 -29852 9384 -29788
rect 9448 -29852 9468 -29788
rect 3169 -29868 9468 -29852
rect 3169 -29932 9384 -29868
rect 9448 -29932 9468 -29868
rect 3169 -29948 9468 -29932
rect 3169 -30012 9384 -29948
rect 9448 -30012 9468 -29948
rect 3169 -30028 9468 -30012
rect 3169 -30092 9384 -30028
rect 9448 -30092 9468 -30028
rect 3169 -30108 9468 -30092
rect 3169 -30172 9384 -30108
rect 9448 -30172 9468 -30108
rect 3169 -30188 9468 -30172
rect 3169 -30252 9384 -30188
rect 9448 -30252 9468 -30188
rect 3169 -30268 9468 -30252
rect 3169 -30332 9384 -30268
rect 9448 -30332 9468 -30268
rect 3169 -30348 9468 -30332
rect 3169 -30412 9384 -30348
rect 9448 -30412 9468 -30348
rect 3169 -30428 9468 -30412
rect 3169 -30492 9384 -30428
rect 9448 -30492 9468 -30428
rect 3169 -30508 9468 -30492
rect 3169 -30572 9384 -30508
rect 9448 -30572 9468 -30508
rect 3169 -30588 9468 -30572
rect 3169 -30652 9384 -30588
rect 9448 -30652 9468 -30588
rect 3169 -30668 9468 -30652
rect 3169 -30732 9384 -30668
rect 9448 -30732 9468 -30668
rect 3169 -30748 9468 -30732
rect 3169 -30812 9384 -30748
rect 9448 -30812 9468 -30748
rect 3169 -30828 9468 -30812
rect 3169 -30892 9384 -30828
rect 9448 -30892 9468 -30828
rect 3169 -30908 9468 -30892
rect 3169 -30972 9384 -30908
rect 9448 -30972 9468 -30908
rect 3169 -30988 9468 -30972
rect 3169 -31052 9384 -30988
rect 9448 -31052 9468 -30988
rect 3169 -31068 9468 -31052
rect 3169 -31132 9384 -31068
rect 9448 -31132 9468 -31068
rect 3169 -31148 9468 -31132
rect 3169 -31212 9384 -31148
rect 9448 -31212 9468 -31148
rect 3169 -31228 9468 -31212
rect 3169 -31292 9384 -31228
rect 9448 -31292 9468 -31228
rect 3169 -31308 9468 -31292
rect 3169 -31372 9384 -31308
rect 9448 -31372 9468 -31308
rect 3169 -31388 9468 -31372
rect 3169 -31452 9384 -31388
rect 9448 -31452 9468 -31388
rect 3169 -31468 9468 -31452
rect 3169 -31532 9384 -31468
rect 9448 -31532 9468 -31468
rect 3169 -31548 9468 -31532
rect 3169 -31612 9384 -31548
rect 9448 -31612 9468 -31548
rect 3169 -31628 9468 -31612
rect 3169 -31692 9384 -31628
rect 9448 -31692 9468 -31628
rect 3169 -31708 9468 -31692
rect 3169 -31772 9384 -31708
rect 9448 -31772 9468 -31708
rect 3169 -31788 9468 -31772
rect 3169 -31852 9384 -31788
rect 9448 -31852 9468 -31788
rect 3169 -31868 9468 -31852
rect 3169 -31932 9384 -31868
rect 9448 -31932 9468 -31868
rect 3169 -31948 9468 -31932
rect 3169 -32012 9384 -31948
rect 9448 -32012 9468 -31948
rect 3169 -32028 9468 -32012
rect 3169 -32092 9384 -32028
rect 9448 -32092 9468 -32028
rect 3169 -32108 9468 -32092
rect 3169 -32172 9384 -32108
rect 9448 -32172 9468 -32108
rect 3169 -32188 9468 -32172
rect 3169 -32252 9384 -32188
rect 9448 -32252 9468 -32188
rect 3169 -32268 9468 -32252
rect 3169 -32332 9384 -32268
rect 9448 -32332 9468 -32268
rect 3169 -32348 9468 -32332
rect 3169 -32412 9384 -32348
rect 9448 -32412 9468 -32348
rect 3169 -32428 9468 -32412
rect 3169 -32492 9384 -32428
rect 9448 -32492 9468 -32428
rect 3169 -32508 9468 -32492
rect 3169 -32572 9384 -32508
rect 9448 -32572 9468 -32508
rect 3169 -32588 9468 -32572
rect 3169 -32652 9384 -32588
rect 9448 -32652 9468 -32588
rect 3169 -32668 9468 -32652
rect 3169 -32732 9384 -32668
rect 9448 -32732 9468 -32668
rect 3169 -32748 9468 -32732
rect 3169 -32812 9384 -32748
rect 9448 -32812 9468 -32748
rect 3169 -32828 9468 -32812
rect 3169 -32892 9384 -32828
rect 9448 -32892 9468 -32828
rect 3169 -32908 9468 -32892
rect 3169 -32972 9384 -32908
rect 9448 -32972 9468 -32908
rect 3169 -32988 9468 -32972
rect 3169 -33052 9384 -32988
rect 9448 -33052 9468 -32988
rect 3169 -33068 9468 -33052
rect 3169 -33132 9384 -33068
rect 9448 -33132 9468 -33068
rect 3169 -33148 9468 -33132
rect 3169 -33212 9384 -33148
rect 9448 -33212 9468 -33148
rect 3169 -33228 9468 -33212
rect 3169 -33292 9384 -33228
rect 9448 -33292 9468 -33228
rect 3169 -33308 9468 -33292
rect 3169 -33372 9384 -33308
rect 9448 -33372 9468 -33308
rect 3169 -33388 9468 -33372
rect 3169 -33452 9384 -33388
rect 9448 -33452 9468 -33388
rect 3169 -33468 9468 -33452
rect 3169 -33532 9384 -33468
rect 9448 -33532 9468 -33468
rect 3169 -33548 9468 -33532
rect 3169 -33612 9384 -33548
rect 9448 -33612 9468 -33548
rect 3169 -33628 9468 -33612
rect 3169 -33692 9384 -33628
rect 9448 -33692 9468 -33628
rect 3169 -33708 9468 -33692
rect 3169 -33772 9384 -33708
rect 9448 -33772 9468 -33708
rect 3169 -33788 9468 -33772
rect 3169 -33852 9384 -33788
rect 9448 -33852 9468 -33788
rect 3169 -33868 9468 -33852
rect 3169 -33932 9384 -33868
rect 9448 -33932 9468 -33868
rect 3169 -33948 9468 -33932
rect 3169 -34012 9384 -33948
rect 9448 -34012 9468 -33948
rect 3169 -34028 9468 -34012
rect 3169 -34092 9384 -34028
rect 9448 -34092 9468 -34028
rect 3169 -34108 9468 -34092
rect 3169 -34172 9384 -34108
rect 9448 -34172 9468 -34108
rect 3169 -34188 9468 -34172
rect 3169 -34252 9384 -34188
rect 9448 -34252 9468 -34188
rect 3169 -34268 9468 -34252
rect 3169 -34332 9384 -34268
rect 9448 -34332 9468 -34268
rect 3169 -34348 9468 -34332
rect 3169 -34412 9384 -34348
rect 9448 -34412 9468 -34348
rect 3169 -34428 9468 -34412
rect 3169 -34492 9384 -34428
rect 9448 -34492 9468 -34428
rect 3169 -34508 9468 -34492
rect 3169 -34572 9384 -34508
rect 9448 -34572 9468 -34508
rect 3169 -34600 9468 -34572
rect 9488 -28428 15787 -28400
rect 9488 -28492 15703 -28428
rect 15767 -28492 15787 -28428
rect 9488 -28508 15787 -28492
rect 9488 -28572 15703 -28508
rect 15767 -28572 15787 -28508
rect 9488 -28588 15787 -28572
rect 9488 -28652 15703 -28588
rect 15767 -28652 15787 -28588
rect 9488 -28668 15787 -28652
rect 9488 -28732 15703 -28668
rect 15767 -28732 15787 -28668
rect 9488 -28748 15787 -28732
rect 9488 -28812 15703 -28748
rect 15767 -28812 15787 -28748
rect 9488 -28828 15787 -28812
rect 9488 -28892 15703 -28828
rect 15767 -28892 15787 -28828
rect 9488 -28908 15787 -28892
rect 9488 -28972 15703 -28908
rect 15767 -28972 15787 -28908
rect 9488 -28988 15787 -28972
rect 9488 -29052 15703 -28988
rect 15767 -29052 15787 -28988
rect 9488 -29068 15787 -29052
rect 9488 -29132 15703 -29068
rect 15767 -29132 15787 -29068
rect 9488 -29148 15787 -29132
rect 9488 -29212 15703 -29148
rect 15767 -29212 15787 -29148
rect 9488 -29228 15787 -29212
rect 9488 -29292 15703 -29228
rect 15767 -29292 15787 -29228
rect 9488 -29308 15787 -29292
rect 9488 -29372 15703 -29308
rect 15767 -29372 15787 -29308
rect 9488 -29388 15787 -29372
rect 9488 -29452 15703 -29388
rect 15767 -29452 15787 -29388
rect 9488 -29468 15787 -29452
rect 9488 -29532 15703 -29468
rect 15767 -29532 15787 -29468
rect 9488 -29548 15787 -29532
rect 9488 -29612 15703 -29548
rect 15767 -29612 15787 -29548
rect 9488 -29628 15787 -29612
rect 9488 -29692 15703 -29628
rect 15767 -29692 15787 -29628
rect 9488 -29708 15787 -29692
rect 9488 -29772 15703 -29708
rect 15767 -29772 15787 -29708
rect 9488 -29788 15787 -29772
rect 9488 -29852 15703 -29788
rect 15767 -29852 15787 -29788
rect 9488 -29868 15787 -29852
rect 9488 -29932 15703 -29868
rect 15767 -29932 15787 -29868
rect 9488 -29948 15787 -29932
rect 9488 -30012 15703 -29948
rect 15767 -30012 15787 -29948
rect 9488 -30028 15787 -30012
rect 9488 -30092 15703 -30028
rect 15767 -30092 15787 -30028
rect 9488 -30108 15787 -30092
rect 9488 -30172 15703 -30108
rect 15767 -30172 15787 -30108
rect 9488 -30188 15787 -30172
rect 9488 -30252 15703 -30188
rect 15767 -30252 15787 -30188
rect 9488 -30268 15787 -30252
rect 9488 -30332 15703 -30268
rect 15767 -30332 15787 -30268
rect 9488 -30348 15787 -30332
rect 9488 -30412 15703 -30348
rect 15767 -30412 15787 -30348
rect 9488 -30428 15787 -30412
rect 9488 -30492 15703 -30428
rect 15767 -30492 15787 -30428
rect 9488 -30508 15787 -30492
rect 9488 -30572 15703 -30508
rect 15767 -30572 15787 -30508
rect 9488 -30588 15787 -30572
rect 9488 -30652 15703 -30588
rect 15767 -30652 15787 -30588
rect 9488 -30668 15787 -30652
rect 9488 -30732 15703 -30668
rect 15767 -30732 15787 -30668
rect 9488 -30748 15787 -30732
rect 9488 -30812 15703 -30748
rect 15767 -30812 15787 -30748
rect 9488 -30828 15787 -30812
rect 9488 -30892 15703 -30828
rect 15767 -30892 15787 -30828
rect 9488 -30908 15787 -30892
rect 9488 -30972 15703 -30908
rect 15767 -30972 15787 -30908
rect 9488 -30988 15787 -30972
rect 9488 -31052 15703 -30988
rect 15767 -31052 15787 -30988
rect 9488 -31068 15787 -31052
rect 9488 -31132 15703 -31068
rect 15767 -31132 15787 -31068
rect 9488 -31148 15787 -31132
rect 9488 -31212 15703 -31148
rect 15767 -31212 15787 -31148
rect 9488 -31228 15787 -31212
rect 9488 -31292 15703 -31228
rect 15767 -31292 15787 -31228
rect 9488 -31308 15787 -31292
rect 9488 -31372 15703 -31308
rect 15767 -31372 15787 -31308
rect 9488 -31388 15787 -31372
rect 9488 -31452 15703 -31388
rect 15767 -31452 15787 -31388
rect 9488 -31468 15787 -31452
rect 9488 -31532 15703 -31468
rect 15767 -31532 15787 -31468
rect 9488 -31548 15787 -31532
rect 9488 -31612 15703 -31548
rect 15767 -31612 15787 -31548
rect 9488 -31628 15787 -31612
rect 9488 -31692 15703 -31628
rect 15767 -31692 15787 -31628
rect 9488 -31708 15787 -31692
rect 9488 -31772 15703 -31708
rect 15767 -31772 15787 -31708
rect 9488 -31788 15787 -31772
rect 9488 -31852 15703 -31788
rect 15767 -31852 15787 -31788
rect 9488 -31868 15787 -31852
rect 9488 -31932 15703 -31868
rect 15767 -31932 15787 -31868
rect 9488 -31948 15787 -31932
rect 9488 -32012 15703 -31948
rect 15767 -32012 15787 -31948
rect 9488 -32028 15787 -32012
rect 9488 -32092 15703 -32028
rect 15767 -32092 15787 -32028
rect 9488 -32108 15787 -32092
rect 9488 -32172 15703 -32108
rect 15767 -32172 15787 -32108
rect 9488 -32188 15787 -32172
rect 9488 -32252 15703 -32188
rect 15767 -32252 15787 -32188
rect 9488 -32268 15787 -32252
rect 9488 -32332 15703 -32268
rect 15767 -32332 15787 -32268
rect 9488 -32348 15787 -32332
rect 9488 -32412 15703 -32348
rect 15767 -32412 15787 -32348
rect 9488 -32428 15787 -32412
rect 9488 -32492 15703 -32428
rect 15767 -32492 15787 -32428
rect 9488 -32508 15787 -32492
rect 9488 -32572 15703 -32508
rect 15767 -32572 15787 -32508
rect 9488 -32588 15787 -32572
rect 9488 -32652 15703 -32588
rect 15767 -32652 15787 -32588
rect 9488 -32668 15787 -32652
rect 9488 -32732 15703 -32668
rect 15767 -32732 15787 -32668
rect 9488 -32748 15787 -32732
rect 9488 -32812 15703 -32748
rect 15767 -32812 15787 -32748
rect 9488 -32828 15787 -32812
rect 9488 -32892 15703 -32828
rect 15767 -32892 15787 -32828
rect 9488 -32908 15787 -32892
rect 9488 -32972 15703 -32908
rect 15767 -32972 15787 -32908
rect 9488 -32988 15787 -32972
rect 9488 -33052 15703 -32988
rect 15767 -33052 15787 -32988
rect 9488 -33068 15787 -33052
rect 9488 -33132 15703 -33068
rect 15767 -33132 15787 -33068
rect 9488 -33148 15787 -33132
rect 9488 -33212 15703 -33148
rect 15767 -33212 15787 -33148
rect 9488 -33228 15787 -33212
rect 9488 -33292 15703 -33228
rect 15767 -33292 15787 -33228
rect 9488 -33308 15787 -33292
rect 9488 -33372 15703 -33308
rect 15767 -33372 15787 -33308
rect 9488 -33388 15787 -33372
rect 9488 -33452 15703 -33388
rect 15767 -33452 15787 -33388
rect 9488 -33468 15787 -33452
rect 9488 -33532 15703 -33468
rect 15767 -33532 15787 -33468
rect 9488 -33548 15787 -33532
rect 9488 -33612 15703 -33548
rect 15767 -33612 15787 -33548
rect 9488 -33628 15787 -33612
rect 9488 -33692 15703 -33628
rect 15767 -33692 15787 -33628
rect 9488 -33708 15787 -33692
rect 9488 -33772 15703 -33708
rect 15767 -33772 15787 -33708
rect 9488 -33788 15787 -33772
rect 9488 -33852 15703 -33788
rect 15767 -33852 15787 -33788
rect 9488 -33868 15787 -33852
rect 9488 -33932 15703 -33868
rect 15767 -33932 15787 -33868
rect 9488 -33948 15787 -33932
rect 9488 -34012 15703 -33948
rect 15767 -34012 15787 -33948
rect 9488 -34028 15787 -34012
rect 9488 -34092 15703 -34028
rect 15767 -34092 15787 -34028
rect 9488 -34108 15787 -34092
rect 9488 -34172 15703 -34108
rect 15767 -34172 15787 -34108
rect 9488 -34188 15787 -34172
rect 9488 -34252 15703 -34188
rect 15767 -34252 15787 -34188
rect 9488 -34268 15787 -34252
rect 9488 -34332 15703 -34268
rect 15767 -34332 15787 -34268
rect 9488 -34348 15787 -34332
rect 9488 -34412 15703 -34348
rect 15767 -34412 15787 -34348
rect 9488 -34428 15787 -34412
rect 9488 -34492 15703 -34428
rect 15767 -34492 15787 -34428
rect 9488 -34508 15787 -34492
rect 9488 -34572 15703 -34508
rect 15767 -34572 15787 -34508
rect 9488 -34600 15787 -34572
rect 15807 -28428 22106 -28400
rect 15807 -28492 22022 -28428
rect 22086 -28492 22106 -28428
rect 15807 -28508 22106 -28492
rect 15807 -28572 22022 -28508
rect 22086 -28572 22106 -28508
rect 15807 -28588 22106 -28572
rect 15807 -28652 22022 -28588
rect 22086 -28652 22106 -28588
rect 15807 -28668 22106 -28652
rect 15807 -28732 22022 -28668
rect 22086 -28732 22106 -28668
rect 15807 -28748 22106 -28732
rect 15807 -28812 22022 -28748
rect 22086 -28812 22106 -28748
rect 15807 -28828 22106 -28812
rect 15807 -28892 22022 -28828
rect 22086 -28892 22106 -28828
rect 15807 -28908 22106 -28892
rect 15807 -28972 22022 -28908
rect 22086 -28972 22106 -28908
rect 15807 -28988 22106 -28972
rect 15807 -29052 22022 -28988
rect 22086 -29052 22106 -28988
rect 15807 -29068 22106 -29052
rect 15807 -29132 22022 -29068
rect 22086 -29132 22106 -29068
rect 15807 -29148 22106 -29132
rect 15807 -29212 22022 -29148
rect 22086 -29212 22106 -29148
rect 15807 -29228 22106 -29212
rect 15807 -29292 22022 -29228
rect 22086 -29292 22106 -29228
rect 15807 -29308 22106 -29292
rect 15807 -29372 22022 -29308
rect 22086 -29372 22106 -29308
rect 15807 -29388 22106 -29372
rect 15807 -29452 22022 -29388
rect 22086 -29452 22106 -29388
rect 15807 -29468 22106 -29452
rect 15807 -29532 22022 -29468
rect 22086 -29532 22106 -29468
rect 15807 -29548 22106 -29532
rect 15807 -29612 22022 -29548
rect 22086 -29612 22106 -29548
rect 15807 -29628 22106 -29612
rect 15807 -29692 22022 -29628
rect 22086 -29692 22106 -29628
rect 15807 -29708 22106 -29692
rect 15807 -29772 22022 -29708
rect 22086 -29772 22106 -29708
rect 15807 -29788 22106 -29772
rect 15807 -29852 22022 -29788
rect 22086 -29852 22106 -29788
rect 15807 -29868 22106 -29852
rect 15807 -29932 22022 -29868
rect 22086 -29932 22106 -29868
rect 15807 -29948 22106 -29932
rect 15807 -30012 22022 -29948
rect 22086 -30012 22106 -29948
rect 15807 -30028 22106 -30012
rect 15807 -30092 22022 -30028
rect 22086 -30092 22106 -30028
rect 15807 -30108 22106 -30092
rect 15807 -30172 22022 -30108
rect 22086 -30172 22106 -30108
rect 15807 -30188 22106 -30172
rect 15807 -30252 22022 -30188
rect 22086 -30252 22106 -30188
rect 15807 -30268 22106 -30252
rect 15807 -30332 22022 -30268
rect 22086 -30332 22106 -30268
rect 15807 -30348 22106 -30332
rect 15807 -30412 22022 -30348
rect 22086 -30412 22106 -30348
rect 15807 -30428 22106 -30412
rect 15807 -30492 22022 -30428
rect 22086 -30492 22106 -30428
rect 15807 -30508 22106 -30492
rect 15807 -30572 22022 -30508
rect 22086 -30572 22106 -30508
rect 15807 -30588 22106 -30572
rect 15807 -30652 22022 -30588
rect 22086 -30652 22106 -30588
rect 15807 -30668 22106 -30652
rect 15807 -30732 22022 -30668
rect 22086 -30732 22106 -30668
rect 15807 -30748 22106 -30732
rect 15807 -30812 22022 -30748
rect 22086 -30812 22106 -30748
rect 15807 -30828 22106 -30812
rect 15807 -30892 22022 -30828
rect 22086 -30892 22106 -30828
rect 15807 -30908 22106 -30892
rect 15807 -30972 22022 -30908
rect 22086 -30972 22106 -30908
rect 15807 -30988 22106 -30972
rect 15807 -31052 22022 -30988
rect 22086 -31052 22106 -30988
rect 15807 -31068 22106 -31052
rect 15807 -31132 22022 -31068
rect 22086 -31132 22106 -31068
rect 15807 -31148 22106 -31132
rect 15807 -31212 22022 -31148
rect 22086 -31212 22106 -31148
rect 15807 -31228 22106 -31212
rect 15807 -31292 22022 -31228
rect 22086 -31292 22106 -31228
rect 15807 -31308 22106 -31292
rect 15807 -31372 22022 -31308
rect 22086 -31372 22106 -31308
rect 15807 -31388 22106 -31372
rect 15807 -31452 22022 -31388
rect 22086 -31452 22106 -31388
rect 15807 -31468 22106 -31452
rect 15807 -31532 22022 -31468
rect 22086 -31532 22106 -31468
rect 15807 -31548 22106 -31532
rect 15807 -31612 22022 -31548
rect 22086 -31612 22106 -31548
rect 15807 -31628 22106 -31612
rect 15807 -31692 22022 -31628
rect 22086 -31692 22106 -31628
rect 15807 -31708 22106 -31692
rect 15807 -31772 22022 -31708
rect 22086 -31772 22106 -31708
rect 15807 -31788 22106 -31772
rect 15807 -31852 22022 -31788
rect 22086 -31852 22106 -31788
rect 15807 -31868 22106 -31852
rect 15807 -31932 22022 -31868
rect 22086 -31932 22106 -31868
rect 15807 -31948 22106 -31932
rect 15807 -32012 22022 -31948
rect 22086 -32012 22106 -31948
rect 15807 -32028 22106 -32012
rect 15807 -32092 22022 -32028
rect 22086 -32092 22106 -32028
rect 15807 -32108 22106 -32092
rect 15807 -32172 22022 -32108
rect 22086 -32172 22106 -32108
rect 15807 -32188 22106 -32172
rect 15807 -32252 22022 -32188
rect 22086 -32252 22106 -32188
rect 15807 -32268 22106 -32252
rect 15807 -32332 22022 -32268
rect 22086 -32332 22106 -32268
rect 15807 -32348 22106 -32332
rect 15807 -32412 22022 -32348
rect 22086 -32412 22106 -32348
rect 15807 -32428 22106 -32412
rect 15807 -32492 22022 -32428
rect 22086 -32492 22106 -32428
rect 15807 -32508 22106 -32492
rect 15807 -32572 22022 -32508
rect 22086 -32572 22106 -32508
rect 15807 -32588 22106 -32572
rect 15807 -32652 22022 -32588
rect 22086 -32652 22106 -32588
rect 15807 -32668 22106 -32652
rect 15807 -32732 22022 -32668
rect 22086 -32732 22106 -32668
rect 15807 -32748 22106 -32732
rect 15807 -32812 22022 -32748
rect 22086 -32812 22106 -32748
rect 15807 -32828 22106 -32812
rect 15807 -32892 22022 -32828
rect 22086 -32892 22106 -32828
rect 15807 -32908 22106 -32892
rect 15807 -32972 22022 -32908
rect 22086 -32972 22106 -32908
rect 15807 -32988 22106 -32972
rect 15807 -33052 22022 -32988
rect 22086 -33052 22106 -32988
rect 15807 -33068 22106 -33052
rect 15807 -33132 22022 -33068
rect 22086 -33132 22106 -33068
rect 15807 -33148 22106 -33132
rect 15807 -33212 22022 -33148
rect 22086 -33212 22106 -33148
rect 15807 -33228 22106 -33212
rect 15807 -33292 22022 -33228
rect 22086 -33292 22106 -33228
rect 15807 -33308 22106 -33292
rect 15807 -33372 22022 -33308
rect 22086 -33372 22106 -33308
rect 15807 -33388 22106 -33372
rect 15807 -33452 22022 -33388
rect 22086 -33452 22106 -33388
rect 15807 -33468 22106 -33452
rect 15807 -33532 22022 -33468
rect 22086 -33532 22106 -33468
rect 15807 -33548 22106 -33532
rect 15807 -33612 22022 -33548
rect 22086 -33612 22106 -33548
rect 15807 -33628 22106 -33612
rect 15807 -33692 22022 -33628
rect 22086 -33692 22106 -33628
rect 15807 -33708 22106 -33692
rect 15807 -33772 22022 -33708
rect 22086 -33772 22106 -33708
rect 15807 -33788 22106 -33772
rect 15807 -33852 22022 -33788
rect 22086 -33852 22106 -33788
rect 15807 -33868 22106 -33852
rect 15807 -33932 22022 -33868
rect 22086 -33932 22106 -33868
rect 15807 -33948 22106 -33932
rect 15807 -34012 22022 -33948
rect 22086 -34012 22106 -33948
rect 15807 -34028 22106 -34012
rect 15807 -34092 22022 -34028
rect 22086 -34092 22106 -34028
rect 15807 -34108 22106 -34092
rect 15807 -34172 22022 -34108
rect 22086 -34172 22106 -34108
rect 15807 -34188 22106 -34172
rect 15807 -34252 22022 -34188
rect 22086 -34252 22106 -34188
rect 15807 -34268 22106 -34252
rect 15807 -34332 22022 -34268
rect 22086 -34332 22106 -34268
rect 15807 -34348 22106 -34332
rect 15807 -34412 22022 -34348
rect 22086 -34412 22106 -34348
rect 15807 -34428 22106 -34412
rect 15807 -34492 22022 -34428
rect 22086 -34492 22106 -34428
rect 15807 -34508 22106 -34492
rect 15807 -34572 22022 -34508
rect 22086 -34572 22106 -34508
rect 15807 -34600 22106 -34572
rect 22126 -28428 28425 -28400
rect 22126 -28492 28341 -28428
rect 28405 -28492 28425 -28428
rect 22126 -28508 28425 -28492
rect 22126 -28572 28341 -28508
rect 28405 -28572 28425 -28508
rect 22126 -28588 28425 -28572
rect 22126 -28652 28341 -28588
rect 28405 -28652 28425 -28588
rect 22126 -28668 28425 -28652
rect 22126 -28732 28341 -28668
rect 28405 -28732 28425 -28668
rect 22126 -28748 28425 -28732
rect 22126 -28812 28341 -28748
rect 28405 -28812 28425 -28748
rect 22126 -28828 28425 -28812
rect 22126 -28892 28341 -28828
rect 28405 -28892 28425 -28828
rect 22126 -28908 28425 -28892
rect 22126 -28972 28341 -28908
rect 28405 -28972 28425 -28908
rect 22126 -28988 28425 -28972
rect 22126 -29052 28341 -28988
rect 28405 -29052 28425 -28988
rect 22126 -29068 28425 -29052
rect 22126 -29132 28341 -29068
rect 28405 -29132 28425 -29068
rect 22126 -29148 28425 -29132
rect 22126 -29212 28341 -29148
rect 28405 -29212 28425 -29148
rect 22126 -29228 28425 -29212
rect 22126 -29292 28341 -29228
rect 28405 -29292 28425 -29228
rect 22126 -29308 28425 -29292
rect 22126 -29372 28341 -29308
rect 28405 -29372 28425 -29308
rect 22126 -29388 28425 -29372
rect 22126 -29452 28341 -29388
rect 28405 -29452 28425 -29388
rect 22126 -29468 28425 -29452
rect 22126 -29532 28341 -29468
rect 28405 -29532 28425 -29468
rect 22126 -29548 28425 -29532
rect 22126 -29612 28341 -29548
rect 28405 -29612 28425 -29548
rect 22126 -29628 28425 -29612
rect 22126 -29692 28341 -29628
rect 28405 -29692 28425 -29628
rect 22126 -29708 28425 -29692
rect 22126 -29772 28341 -29708
rect 28405 -29772 28425 -29708
rect 22126 -29788 28425 -29772
rect 22126 -29852 28341 -29788
rect 28405 -29852 28425 -29788
rect 22126 -29868 28425 -29852
rect 22126 -29932 28341 -29868
rect 28405 -29932 28425 -29868
rect 22126 -29948 28425 -29932
rect 22126 -30012 28341 -29948
rect 28405 -30012 28425 -29948
rect 22126 -30028 28425 -30012
rect 22126 -30092 28341 -30028
rect 28405 -30092 28425 -30028
rect 22126 -30108 28425 -30092
rect 22126 -30172 28341 -30108
rect 28405 -30172 28425 -30108
rect 22126 -30188 28425 -30172
rect 22126 -30252 28341 -30188
rect 28405 -30252 28425 -30188
rect 22126 -30268 28425 -30252
rect 22126 -30332 28341 -30268
rect 28405 -30332 28425 -30268
rect 22126 -30348 28425 -30332
rect 22126 -30412 28341 -30348
rect 28405 -30412 28425 -30348
rect 22126 -30428 28425 -30412
rect 22126 -30492 28341 -30428
rect 28405 -30492 28425 -30428
rect 22126 -30508 28425 -30492
rect 22126 -30572 28341 -30508
rect 28405 -30572 28425 -30508
rect 22126 -30588 28425 -30572
rect 22126 -30652 28341 -30588
rect 28405 -30652 28425 -30588
rect 22126 -30668 28425 -30652
rect 22126 -30732 28341 -30668
rect 28405 -30732 28425 -30668
rect 22126 -30748 28425 -30732
rect 22126 -30812 28341 -30748
rect 28405 -30812 28425 -30748
rect 22126 -30828 28425 -30812
rect 22126 -30892 28341 -30828
rect 28405 -30892 28425 -30828
rect 22126 -30908 28425 -30892
rect 22126 -30972 28341 -30908
rect 28405 -30972 28425 -30908
rect 22126 -30988 28425 -30972
rect 22126 -31052 28341 -30988
rect 28405 -31052 28425 -30988
rect 22126 -31068 28425 -31052
rect 22126 -31132 28341 -31068
rect 28405 -31132 28425 -31068
rect 22126 -31148 28425 -31132
rect 22126 -31212 28341 -31148
rect 28405 -31212 28425 -31148
rect 22126 -31228 28425 -31212
rect 22126 -31292 28341 -31228
rect 28405 -31292 28425 -31228
rect 22126 -31308 28425 -31292
rect 22126 -31372 28341 -31308
rect 28405 -31372 28425 -31308
rect 22126 -31388 28425 -31372
rect 22126 -31452 28341 -31388
rect 28405 -31452 28425 -31388
rect 22126 -31468 28425 -31452
rect 22126 -31532 28341 -31468
rect 28405 -31532 28425 -31468
rect 22126 -31548 28425 -31532
rect 22126 -31612 28341 -31548
rect 28405 -31612 28425 -31548
rect 22126 -31628 28425 -31612
rect 22126 -31692 28341 -31628
rect 28405 -31692 28425 -31628
rect 22126 -31708 28425 -31692
rect 22126 -31772 28341 -31708
rect 28405 -31772 28425 -31708
rect 22126 -31788 28425 -31772
rect 22126 -31852 28341 -31788
rect 28405 -31852 28425 -31788
rect 22126 -31868 28425 -31852
rect 22126 -31932 28341 -31868
rect 28405 -31932 28425 -31868
rect 22126 -31948 28425 -31932
rect 22126 -32012 28341 -31948
rect 28405 -32012 28425 -31948
rect 22126 -32028 28425 -32012
rect 22126 -32092 28341 -32028
rect 28405 -32092 28425 -32028
rect 22126 -32108 28425 -32092
rect 22126 -32172 28341 -32108
rect 28405 -32172 28425 -32108
rect 22126 -32188 28425 -32172
rect 22126 -32252 28341 -32188
rect 28405 -32252 28425 -32188
rect 22126 -32268 28425 -32252
rect 22126 -32332 28341 -32268
rect 28405 -32332 28425 -32268
rect 22126 -32348 28425 -32332
rect 22126 -32412 28341 -32348
rect 28405 -32412 28425 -32348
rect 22126 -32428 28425 -32412
rect 22126 -32492 28341 -32428
rect 28405 -32492 28425 -32428
rect 22126 -32508 28425 -32492
rect 22126 -32572 28341 -32508
rect 28405 -32572 28425 -32508
rect 22126 -32588 28425 -32572
rect 22126 -32652 28341 -32588
rect 28405 -32652 28425 -32588
rect 22126 -32668 28425 -32652
rect 22126 -32732 28341 -32668
rect 28405 -32732 28425 -32668
rect 22126 -32748 28425 -32732
rect 22126 -32812 28341 -32748
rect 28405 -32812 28425 -32748
rect 22126 -32828 28425 -32812
rect 22126 -32892 28341 -32828
rect 28405 -32892 28425 -32828
rect 22126 -32908 28425 -32892
rect 22126 -32972 28341 -32908
rect 28405 -32972 28425 -32908
rect 22126 -32988 28425 -32972
rect 22126 -33052 28341 -32988
rect 28405 -33052 28425 -32988
rect 22126 -33068 28425 -33052
rect 22126 -33132 28341 -33068
rect 28405 -33132 28425 -33068
rect 22126 -33148 28425 -33132
rect 22126 -33212 28341 -33148
rect 28405 -33212 28425 -33148
rect 22126 -33228 28425 -33212
rect 22126 -33292 28341 -33228
rect 28405 -33292 28425 -33228
rect 22126 -33308 28425 -33292
rect 22126 -33372 28341 -33308
rect 28405 -33372 28425 -33308
rect 22126 -33388 28425 -33372
rect 22126 -33452 28341 -33388
rect 28405 -33452 28425 -33388
rect 22126 -33468 28425 -33452
rect 22126 -33532 28341 -33468
rect 28405 -33532 28425 -33468
rect 22126 -33548 28425 -33532
rect 22126 -33612 28341 -33548
rect 28405 -33612 28425 -33548
rect 22126 -33628 28425 -33612
rect 22126 -33692 28341 -33628
rect 28405 -33692 28425 -33628
rect 22126 -33708 28425 -33692
rect 22126 -33772 28341 -33708
rect 28405 -33772 28425 -33708
rect 22126 -33788 28425 -33772
rect 22126 -33852 28341 -33788
rect 28405 -33852 28425 -33788
rect 22126 -33868 28425 -33852
rect 22126 -33932 28341 -33868
rect 28405 -33932 28425 -33868
rect 22126 -33948 28425 -33932
rect 22126 -34012 28341 -33948
rect 28405 -34012 28425 -33948
rect 22126 -34028 28425 -34012
rect 22126 -34092 28341 -34028
rect 28405 -34092 28425 -34028
rect 22126 -34108 28425 -34092
rect 22126 -34172 28341 -34108
rect 28405 -34172 28425 -34108
rect 22126 -34188 28425 -34172
rect 22126 -34252 28341 -34188
rect 28405 -34252 28425 -34188
rect 22126 -34268 28425 -34252
rect 22126 -34332 28341 -34268
rect 28405 -34332 28425 -34268
rect 22126 -34348 28425 -34332
rect 22126 -34412 28341 -34348
rect 28405 -34412 28425 -34348
rect 22126 -34428 28425 -34412
rect 22126 -34492 28341 -34428
rect 28405 -34492 28425 -34428
rect 22126 -34508 28425 -34492
rect 22126 -34572 28341 -34508
rect 28405 -34572 28425 -34508
rect 22126 -34600 28425 -34572
rect 28445 -28428 34744 -28400
rect 28445 -28492 34660 -28428
rect 34724 -28492 34744 -28428
rect 28445 -28508 34744 -28492
rect 28445 -28572 34660 -28508
rect 34724 -28572 34744 -28508
rect 28445 -28588 34744 -28572
rect 28445 -28652 34660 -28588
rect 34724 -28652 34744 -28588
rect 28445 -28668 34744 -28652
rect 28445 -28732 34660 -28668
rect 34724 -28732 34744 -28668
rect 28445 -28748 34744 -28732
rect 28445 -28812 34660 -28748
rect 34724 -28812 34744 -28748
rect 28445 -28828 34744 -28812
rect 28445 -28892 34660 -28828
rect 34724 -28892 34744 -28828
rect 28445 -28908 34744 -28892
rect 28445 -28972 34660 -28908
rect 34724 -28972 34744 -28908
rect 28445 -28988 34744 -28972
rect 28445 -29052 34660 -28988
rect 34724 -29052 34744 -28988
rect 28445 -29068 34744 -29052
rect 28445 -29132 34660 -29068
rect 34724 -29132 34744 -29068
rect 28445 -29148 34744 -29132
rect 28445 -29212 34660 -29148
rect 34724 -29212 34744 -29148
rect 28445 -29228 34744 -29212
rect 28445 -29292 34660 -29228
rect 34724 -29292 34744 -29228
rect 28445 -29308 34744 -29292
rect 28445 -29372 34660 -29308
rect 34724 -29372 34744 -29308
rect 28445 -29388 34744 -29372
rect 28445 -29452 34660 -29388
rect 34724 -29452 34744 -29388
rect 28445 -29468 34744 -29452
rect 28445 -29532 34660 -29468
rect 34724 -29532 34744 -29468
rect 28445 -29548 34744 -29532
rect 28445 -29612 34660 -29548
rect 34724 -29612 34744 -29548
rect 28445 -29628 34744 -29612
rect 28445 -29692 34660 -29628
rect 34724 -29692 34744 -29628
rect 28445 -29708 34744 -29692
rect 28445 -29772 34660 -29708
rect 34724 -29772 34744 -29708
rect 28445 -29788 34744 -29772
rect 28445 -29852 34660 -29788
rect 34724 -29852 34744 -29788
rect 28445 -29868 34744 -29852
rect 28445 -29932 34660 -29868
rect 34724 -29932 34744 -29868
rect 28445 -29948 34744 -29932
rect 28445 -30012 34660 -29948
rect 34724 -30012 34744 -29948
rect 28445 -30028 34744 -30012
rect 28445 -30092 34660 -30028
rect 34724 -30092 34744 -30028
rect 28445 -30108 34744 -30092
rect 28445 -30172 34660 -30108
rect 34724 -30172 34744 -30108
rect 28445 -30188 34744 -30172
rect 28445 -30252 34660 -30188
rect 34724 -30252 34744 -30188
rect 28445 -30268 34744 -30252
rect 28445 -30332 34660 -30268
rect 34724 -30332 34744 -30268
rect 28445 -30348 34744 -30332
rect 28445 -30412 34660 -30348
rect 34724 -30412 34744 -30348
rect 28445 -30428 34744 -30412
rect 28445 -30492 34660 -30428
rect 34724 -30492 34744 -30428
rect 28445 -30508 34744 -30492
rect 28445 -30572 34660 -30508
rect 34724 -30572 34744 -30508
rect 28445 -30588 34744 -30572
rect 28445 -30652 34660 -30588
rect 34724 -30652 34744 -30588
rect 28445 -30668 34744 -30652
rect 28445 -30732 34660 -30668
rect 34724 -30732 34744 -30668
rect 28445 -30748 34744 -30732
rect 28445 -30812 34660 -30748
rect 34724 -30812 34744 -30748
rect 28445 -30828 34744 -30812
rect 28445 -30892 34660 -30828
rect 34724 -30892 34744 -30828
rect 28445 -30908 34744 -30892
rect 28445 -30972 34660 -30908
rect 34724 -30972 34744 -30908
rect 28445 -30988 34744 -30972
rect 28445 -31052 34660 -30988
rect 34724 -31052 34744 -30988
rect 28445 -31068 34744 -31052
rect 28445 -31132 34660 -31068
rect 34724 -31132 34744 -31068
rect 28445 -31148 34744 -31132
rect 28445 -31212 34660 -31148
rect 34724 -31212 34744 -31148
rect 28445 -31228 34744 -31212
rect 28445 -31292 34660 -31228
rect 34724 -31292 34744 -31228
rect 28445 -31308 34744 -31292
rect 28445 -31372 34660 -31308
rect 34724 -31372 34744 -31308
rect 28445 -31388 34744 -31372
rect 28445 -31452 34660 -31388
rect 34724 -31452 34744 -31388
rect 28445 -31468 34744 -31452
rect 28445 -31532 34660 -31468
rect 34724 -31532 34744 -31468
rect 28445 -31548 34744 -31532
rect 28445 -31612 34660 -31548
rect 34724 -31612 34744 -31548
rect 28445 -31628 34744 -31612
rect 28445 -31692 34660 -31628
rect 34724 -31692 34744 -31628
rect 28445 -31708 34744 -31692
rect 28445 -31772 34660 -31708
rect 34724 -31772 34744 -31708
rect 28445 -31788 34744 -31772
rect 28445 -31852 34660 -31788
rect 34724 -31852 34744 -31788
rect 28445 -31868 34744 -31852
rect 28445 -31932 34660 -31868
rect 34724 -31932 34744 -31868
rect 28445 -31948 34744 -31932
rect 28445 -32012 34660 -31948
rect 34724 -32012 34744 -31948
rect 28445 -32028 34744 -32012
rect 28445 -32092 34660 -32028
rect 34724 -32092 34744 -32028
rect 28445 -32108 34744 -32092
rect 28445 -32172 34660 -32108
rect 34724 -32172 34744 -32108
rect 28445 -32188 34744 -32172
rect 28445 -32252 34660 -32188
rect 34724 -32252 34744 -32188
rect 28445 -32268 34744 -32252
rect 28445 -32332 34660 -32268
rect 34724 -32332 34744 -32268
rect 28445 -32348 34744 -32332
rect 28445 -32412 34660 -32348
rect 34724 -32412 34744 -32348
rect 28445 -32428 34744 -32412
rect 28445 -32492 34660 -32428
rect 34724 -32492 34744 -32428
rect 28445 -32508 34744 -32492
rect 28445 -32572 34660 -32508
rect 34724 -32572 34744 -32508
rect 28445 -32588 34744 -32572
rect 28445 -32652 34660 -32588
rect 34724 -32652 34744 -32588
rect 28445 -32668 34744 -32652
rect 28445 -32732 34660 -32668
rect 34724 -32732 34744 -32668
rect 28445 -32748 34744 -32732
rect 28445 -32812 34660 -32748
rect 34724 -32812 34744 -32748
rect 28445 -32828 34744 -32812
rect 28445 -32892 34660 -32828
rect 34724 -32892 34744 -32828
rect 28445 -32908 34744 -32892
rect 28445 -32972 34660 -32908
rect 34724 -32972 34744 -32908
rect 28445 -32988 34744 -32972
rect 28445 -33052 34660 -32988
rect 34724 -33052 34744 -32988
rect 28445 -33068 34744 -33052
rect 28445 -33132 34660 -33068
rect 34724 -33132 34744 -33068
rect 28445 -33148 34744 -33132
rect 28445 -33212 34660 -33148
rect 34724 -33212 34744 -33148
rect 28445 -33228 34744 -33212
rect 28445 -33292 34660 -33228
rect 34724 -33292 34744 -33228
rect 28445 -33308 34744 -33292
rect 28445 -33372 34660 -33308
rect 34724 -33372 34744 -33308
rect 28445 -33388 34744 -33372
rect 28445 -33452 34660 -33388
rect 34724 -33452 34744 -33388
rect 28445 -33468 34744 -33452
rect 28445 -33532 34660 -33468
rect 34724 -33532 34744 -33468
rect 28445 -33548 34744 -33532
rect 28445 -33612 34660 -33548
rect 34724 -33612 34744 -33548
rect 28445 -33628 34744 -33612
rect 28445 -33692 34660 -33628
rect 34724 -33692 34744 -33628
rect 28445 -33708 34744 -33692
rect 28445 -33772 34660 -33708
rect 34724 -33772 34744 -33708
rect 28445 -33788 34744 -33772
rect 28445 -33852 34660 -33788
rect 34724 -33852 34744 -33788
rect 28445 -33868 34744 -33852
rect 28445 -33932 34660 -33868
rect 34724 -33932 34744 -33868
rect 28445 -33948 34744 -33932
rect 28445 -34012 34660 -33948
rect 34724 -34012 34744 -33948
rect 28445 -34028 34744 -34012
rect 28445 -34092 34660 -34028
rect 34724 -34092 34744 -34028
rect 28445 -34108 34744 -34092
rect 28445 -34172 34660 -34108
rect 34724 -34172 34744 -34108
rect 28445 -34188 34744 -34172
rect 28445 -34252 34660 -34188
rect 34724 -34252 34744 -34188
rect 28445 -34268 34744 -34252
rect 28445 -34332 34660 -34268
rect 34724 -34332 34744 -34268
rect 28445 -34348 34744 -34332
rect 28445 -34412 34660 -34348
rect 34724 -34412 34744 -34348
rect 28445 -34428 34744 -34412
rect 28445 -34492 34660 -34428
rect 34724 -34492 34744 -34428
rect 28445 -34508 34744 -34492
rect 28445 -34572 34660 -34508
rect 34724 -34572 34744 -34508
rect 28445 -34600 34744 -34572
rect 34764 -28428 41063 -28400
rect 34764 -28492 40979 -28428
rect 41043 -28492 41063 -28428
rect 34764 -28508 41063 -28492
rect 34764 -28572 40979 -28508
rect 41043 -28572 41063 -28508
rect 34764 -28588 41063 -28572
rect 34764 -28652 40979 -28588
rect 41043 -28652 41063 -28588
rect 34764 -28668 41063 -28652
rect 34764 -28732 40979 -28668
rect 41043 -28732 41063 -28668
rect 34764 -28748 41063 -28732
rect 34764 -28812 40979 -28748
rect 41043 -28812 41063 -28748
rect 34764 -28828 41063 -28812
rect 34764 -28892 40979 -28828
rect 41043 -28892 41063 -28828
rect 34764 -28908 41063 -28892
rect 34764 -28972 40979 -28908
rect 41043 -28972 41063 -28908
rect 34764 -28988 41063 -28972
rect 34764 -29052 40979 -28988
rect 41043 -29052 41063 -28988
rect 34764 -29068 41063 -29052
rect 34764 -29132 40979 -29068
rect 41043 -29132 41063 -29068
rect 34764 -29148 41063 -29132
rect 34764 -29212 40979 -29148
rect 41043 -29212 41063 -29148
rect 34764 -29228 41063 -29212
rect 34764 -29292 40979 -29228
rect 41043 -29292 41063 -29228
rect 34764 -29308 41063 -29292
rect 34764 -29372 40979 -29308
rect 41043 -29372 41063 -29308
rect 34764 -29388 41063 -29372
rect 34764 -29452 40979 -29388
rect 41043 -29452 41063 -29388
rect 34764 -29468 41063 -29452
rect 34764 -29532 40979 -29468
rect 41043 -29532 41063 -29468
rect 34764 -29548 41063 -29532
rect 34764 -29612 40979 -29548
rect 41043 -29612 41063 -29548
rect 34764 -29628 41063 -29612
rect 34764 -29692 40979 -29628
rect 41043 -29692 41063 -29628
rect 34764 -29708 41063 -29692
rect 34764 -29772 40979 -29708
rect 41043 -29772 41063 -29708
rect 34764 -29788 41063 -29772
rect 34764 -29852 40979 -29788
rect 41043 -29852 41063 -29788
rect 34764 -29868 41063 -29852
rect 34764 -29932 40979 -29868
rect 41043 -29932 41063 -29868
rect 34764 -29948 41063 -29932
rect 34764 -30012 40979 -29948
rect 41043 -30012 41063 -29948
rect 34764 -30028 41063 -30012
rect 34764 -30092 40979 -30028
rect 41043 -30092 41063 -30028
rect 34764 -30108 41063 -30092
rect 34764 -30172 40979 -30108
rect 41043 -30172 41063 -30108
rect 34764 -30188 41063 -30172
rect 34764 -30252 40979 -30188
rect 41043 -30252 41063 -30188
rect 34764 -30268 41063 -30252
rect 34764 -30332 40979 -30268
rect 41043 -30332 41063 -30268
rect 34764 -30348 41063 -30332
rect 34764 -30412 40979 -30348
rect 41043 -30412 41063 -30348
rect 34764 -30428 41063 -30412
rect 34764 -30492 40979 -30428
rect 41043 -30492 41063 -30428
rect 34764 -30508 41063 -30492
rect 34764 -30572 40979 -30508
rect 41043 -30572 41063 -30508
rect 34764 -30588 41063 -30572
rect 34764 -30652 40979 -30588
rect 41043 -30652 41063 -30588
rect 34764 -30668 41063 -30652
rect 34764 -30732 40979 -30668
rect 41043 -30732 41063 -30668
rect 34764 -30748 41063 -30732
rect 34764 -30812 40979 -30748
rect 41043 -30812 41063 -30748
rect 34764 -30828 41063 -30812
rect 34764 -30892 40979 -30828
rect 41043 -30892 41063 -30828
rect 34764 -30908 41063 -30892
rect 34764 -30972 40979 -30908
rect 41043 -30972 41063 -30908
rect 34764 -30988 41063 -30972
rect 34764 -31052 40979 -30988
rect 41043 -31052 41063 -30988
rect 34764 -31068 41063 -31052
rect 34764 -31132 40979 -31068
rect 41043 -31132 41063 -31068
rect 34764 -31148 41063 -31132
rect 34764 -31212 40979 -31148
rect 41043 -31212 41063 -31148
rect 34764 -31228 41063 -31212
rect 34764 -31292 40979 -31228
rect 41043 -31292 41063 -31228
rect 34764 -31308 41063 -31292
rect 34764 -31372 40979 -31308
rect 41043 -31372 41063 -31308
rect 34764 -31388 41063 -31372
rect 34764 -31452 40979 -31388
rect 41043 -31452 41063 -31388
rect 34764 -31468 41063 -31452
rect 34764 -31532 40979 -31468
rect 41043 -31532 41063 -31468
rect 34764 -31548 41063 -31532
rect 34764 -31612 40979 -31548
rect 41043 -31612 41063 -31548
rect 34764 -31628 41063 -31612
rect 34764 -31692 40979 -31628
rect 41043 -31692 41063 -31628
rect 34764 -31708 41063 -31692
rect 34764 -31772 40979 -31708
rect 41043 -31772 41063 -31708
rect 34764 -31788 41063 -31772
rect 34764 -31852 40979 -31788
rect 41043 -31852 41063 -31788
rect 34764 -31868 41063 -31852
rect 34764 -31932 40979 -31868
rect 41043 -31932 41063 -31868
rect 34764 -31948 41063 -31932
rect 34764 -32012 40979 -31948
rect 41043 -32012 41063 -31948
rect 34764 -32028 41063 -32012
rect 34764 -32092 40979 -32028
rect 41043 -32092 41063 -32028
rect 34764 -32108 41063 -32092
rect 34764 -32172 40979 -32108
rect 41043 -32172 41063 -32108
rect 34764 -32188 41063 -32172
rect 34764 -32252 40979 -32188
rect 41043 -32252 41063 -32188
rect 34764 -32268 41063 -32252
rect 34764 -32332 40979 -32268
rect 41043 -32332 41063 -32268
rect 34764 -32348 41063 -32332
rect 34764 -32412 40979 -32348
rect 41043 -32412 41063 -32348
rect 34764 -32428 41063 -32412
rect 34764 -32492 40979 -32428
rect 41043 -32492 41063 -32428
rect 34764 -32508 41063 -32492
rect 34764 -32572 40979 -32508
rect 41043 -32572 41063 -32508
rect 34764 -32588 41063 -32572
rect 34764 -32652 40979 -32588
rect 41043 -32652 41063 -32588
rect 34764 -32668 41063 -32652
rect 34764 -32732 40979 -32668
rect 41043 -32732 41063 -32668
rect 34764 -32748 41063 -32732
rect 34764 -32812 40979 -32748
rect 41043 -32812 41063 -32748
rect 34764 -32828 41063 -32812
rect 34764 -32892 40979 -32828
rect 41043 -32892 41063 -32828
rect 34764 -32908 41063 -32892
rect 34764 -32972 40979 -32908
rect 41043 -32972 41063 -32908
rect 34764 -32988 41063 -32972
rect 34764 -33052 40979 -32988
rect 41043 -33052 41063 -32988
rect 34764 -33068 41063 -33052
rect 34764 -33132 40979 -33068
rect 41043 -33132 41063 -33068
rect 34764 -33148 41063 -33132
rect 34764 -33212 40979 -33148
rect 41043 -33212 41063 -33148
rect 34764 -33228 41063 -33212
rect 34764 -33292 40979 -33228
rect 41043 -33292 41063 -33228
rect 34764 -33308 41063 -33292
rect 34764 -33372 40979 -33308
rect 41043 -33372 41063 -33308
rect 34764 -33388 41063 -33372
rect 34764 -33452 40979 -33388
rect 41043 -33452 41063 -33388
rect 34764 -33468 41063 -33452
rect 34764 -33532 40979 -33468
rect 41043 -33532 41063 -33468
rect 34764 -33548 41063 -33532
rect 34764 -33612 40979 -33548
rect 41043 -33612 41063 -33548
rect 34764 -33628 41063 -33612
rect 34764 -33692 40979 -33628
rect 41043 -33692 41063 -33628
rect 34764 -33708 41063 -33692
rect 34764 -33772 40979 -33708
rect 41043 -33772 41063 -33708
rect 34764 -33788 41063 -33772
rect 34764 -33852 40979 -33788
rect 41043 -33852 41063 -33788
rect 34764 -33868 41063 -33852
rect 34764 -33932 40979 -33868
rect 41043 -33932 41063 -33868
rect 34764 -33948 41063 -33932
rect 34764 -34012 40979 -33948
rect 41043 -34012 41063 -33948
rect 34764 -34028 41063 -34012
rect 34764 -34092 40979 -34028
rect 41043 -34092 41063 -34028
rect 34764 -34108 41063 -34092
rect 34764 -34172 40979 -34108
rect 41043 -34172 41063 -34108
rect 34764 -34188 41063 -34172
rect 34764 -34252 40979 -34188
rect 41043 -34252 41063 -34188
rect 34764 -34268 41063 -34252
rect 34764 -34332 40979 -34268
rect 41043 -34332 41063 -34268
rect 34764 -34348 41063 -34332
rect 34764 -34412 40979 -34348
rect 41043 -34412 41063 -34348
rect 34764 -34428 41063 -34412
rect 34764 -34492 40979 -34428
rect 41043 -34492 41063 -34428
rect 34764 -34508 41063 -34492
rect 34764 -34572 40979 -34508
rect 41043 -34572 41063 -34508
rect 34764 -34600 41063 -34572
rect 41083 -28428 47382 -28400
rect 41083 -28492 47298 -28428
rect 47362 -28492 47382 -28428
rect 41083 -28508 47382 -28492
rect 41083 -28572 47298 -28508
rect 47362 -28572 47382 -28508
rect 41083 -28588 47382 -28572
rect 41083 -28652 47298 -28588
rect 47362 -28652 47382 -28588
rect 41083 -28668 47382 -28652
rect 41083 -28732 47298 -28668
rect 47362 -28732 47382 -28668
rect 41083 -28748 47382 -28732
rect 41083 -28812 47298 -28748
rect 47362 -28812 47382 -28748
rect 41083 -28828 47382 -28812
rect 41083 -28892 47298 -28828
rect 47362 -28892 47382 -28828
rect 41083 -28908 47382 -28892
rect 41083 -28972 47298 -28908
rect 47362 -28972 47382 -28908
rect 41083 -28988 47382 -28972
rect 41083 -29052 47298 -28988
rect 47362 -29052 47382 -28988
rect 41083 -29068 47382 -29052
rect 41083 -29132 47298 -29068
rect 47362 -29132 47382 -29068
rect 41083 -29148 47382 -29132
rect 41083 -29212 47298 -29148
rect 47362 -29212 47382 -29148
rect 41083 -29228 47382 -29212
rect 41083 -29292 47298 -29228
rect 47362 -29292 47382 -29228
rect 41083 -29308 47382 -29292
rect 41083 -29372 47298 -29308
rect 47362 -29372 47382 -29308
rect 41083 -29388 47382 -29372
rect 41083 -29452 47298 -29388
rect 47362 -29452 47382 -29388
rect 41083 -29468 47382 -29452
rect 41083 -29532 47298 -29468
rect 47362 -29532 47382 -29468
rect 41083 -29548 47382 -29532
rect 41083 -29612 47298 -29548
rect 47362 -29612 47382 -29548
rect 41083 -29628 47382 -29612
rect 41083 -29692 47298 -29628
rect 47362 -29692 47382 -29628
rect 41083 -29708 47382 -29692
rect 41083 -29772 47298 -29708
rect 47362 -29772 47382 -29708
rect 41083 -29788 47382 -29772
rect 41083 -29852 47298 -29788
rect 47362 -29852 47382 -29788
rect 41083 -29868 47382 -29852
rect 41083 -29932 47298 -29868
rect 47362 -29932 47382 -29868
rect 41083 -29948 47382 -29932
rect 41083 -30012 47298 -29948
rect 47362 -30012 47382 -29948
rect 41083 -30028 47382 -30012
rect 41083 -30092 47298 -30028
rect 47362 -30092 47382 -30028
rect 41083 -30108 47382 -30092
rect 41083 -30172 47298 -30108
rect 47362 -30172 47382 -30108
rect 41083 -30188 47382 -30172
rect 41083 -30252 47298 -30188
rect 47362 -30252 47382 -30188
rect 41083 -30268 47382 -30252
rect 41083 -30332 47298 -30268
rect 47362 -30332 47382 -30268
rect 41083 -30348 47382 -30332
rect 41083 -30412 47298 -30348
rect 47362 -30412 47382 -30348
rect 41083 -30428 47382 -30412
rect 41083 -30492 47298 -30428
rect 47362 -30492 47382 -30428
rect 41083 -30508 47382 -30492
rect 41083 -30572 47298 -30508
rect 47362 -30572 47382 -30508
rect 41083 -30588 47382 -30572
rect 41083 -30652 47298 -30588
rect 47362 -30652 47382 -30588
rect 41083 -30668 47382 -30652
rect 41083 -30732 47298 -30668
rect 47362 -30732 47382 -30668
rect 41083 -30748 47382 -30732
rect 41083 -30812 47298 -30748
rect 47362 -30812 47382 -30748
rect 41083 -30828 47382 -30812
rect 41083 -30892 47298 -30828
rect 47362 -30892 47382 -30828
rect 41083 -30908 47382 -30892
rect 41083 -30972 47298 -30908
rect 47362 -30972 47382 -30908
rect 41083 -30988 47382 -30972
rect 41083 -31052 47298 -30988
rect 47362 -31052 47382 -30988
rect 41083 -31068 47382 -31052
rect 41083 -31132 47298 -31068
rect 47362 -31132 47382 -31068
rect 41083 -31148 47382 -31132
rect 41083 -31212 47298 -31148
rect 47362 -31212 47382 -31148
rect 41083 -31228 47382 -31212
rect 41083 -31292 47298 -31228
rect 47362 -31292 47382 -31228
rect 41083 -31308 47382 -31292
rect 41083 -31372 47298 -31308
rect 47362 -31372 47382 -31308
rect 41083 -31388 47382 -31372
rect 41083 -31452 47298 -31388
rect 47362 -31452 47382 -31388
rect 41083 -31468 47382 -31452
rect 41083 -31532 47298 -31468
rect 47362 -31532 47382 -31468
rect 41083 -31548 47382 -31532
rect 41083 -31612 47298 -31548
rect 47362 -31612 47382 -31548
rect 41083 -31628 47382 -31612
rect 41083 -31692 47298 -31628
rect 47362 -31692 47382 -31628
rect 41083 -31708 47382 -31692
rect 41083 -31772 47298 -31708
rect 47362 -31772 47382 -31708
rect 41083 -31788 47382 -31772
rect 41083 -31852 47298 -31788
rect 47362 -31852 47382 -31788
rect 41083 -31868 47382 -31852
rect 41083 -31932 47298 -31868
rect 47362 -31932 47382 -31868
rect 41083 -31948 47382 -31932
rect 41083 -32012 47298 -31948
rect 47362 -32012 47382 -31948
rect 41083 -32028 47382 -32012
rect 41083 -32092 47298 -32028
rect 47362 -32092 47382 -32028
rect 41083 -32108 47382 -32092
rect 41083 -32172 47298 -32108
rect 47362 -32172 47382 -32108
rect 41083 -32188 47382 -32172
rect 41083 -32252 47298 -32188
rect 47362 -32252 47382 -32188
rect 41083 -32268 47382 -32252
rect 41083 -32332 47298 -32268
rect 47362 -32332 47382 -32268
rect 41083 -32348 47382 -32332
rect 41083 -32412 47298 -32348
rect 47362 -32412 47382 -32348
rect 41083 -32428 47382 -32412
rect 41083 -32492 47298 -32428
rect 47362 -32492 47382 -32428
rect 41083 -32508 47382 -32492
rect 41083 -32572 47298 -32508
rect 47362 -32572 47382 -32508
rect 41083 -32588 47382 -32572
rect 41083 -32652 47298 -32588
rect 47362 -32652 47382 -32588
rect 41083 -32668 47382 -32652
rect 41083 -32732 47298 -32668
rect 47362 -32732 47382 -32668
rect 41083 -32748 47382 -32732
rect 41083 -32812 47298 -32748
rect 47362 -32812 47382 -32748
rect 41083 -32828 47382 -32812
rect 41083 -32892 47298 -32828
rect 47362 -32892 47382 -32828
rect 41083 -32908 47382 -32892
rect 41083 -32972 47298 -32908
rect 47362 -32972 47382 -32908
rect 41083 -32988 47382 -32972
rect 41083 -33052 47298 -32988
rect 47362 -33052 47382 -32988
rect 41083 -33068 47382 -33052
rect 41083 -33132 47298 -33068
rect 47362 -33132 47382 -33068
rect 41083 -33148 47382 -33132
rect 41083 -33212 47298 -33148
rect 47362 -33212 47382 -33148
rect 41083 -33228 47382 -33212
rect 41083 -33292 47298 -33228
rect 47362 -33292 47382 -33228
rect 41083 -33308 47382 -33292
rect 41083 -33372 47298 -33308
rect 47362 -33372 47382 -33308
rect 41083 -33388 47382 -33372
rect 41083 -33452 47298 -33388
rect 47362 -33452 47382 -33388
rect 41083 -33468 47382 -33452
rect 41083 -33532 47298 -33468
rect 47362 -33532 47382 -33468
rect 41083 -33548 47382 -33532
rect 41083 -33612 47298 -33548
rect 47362 -33612 47382 -33548
rect 41083 -33628 47382 -33612
rect 41083 -33692 47298 -33628
rect 47362 -33692 47382 -33628
rect 41083 -33708 47382 -33692
rect 41083 -33772 47298 -33708
rect 47362 -33772 47382 -33708
rect 41083 -33788 47382 -33772
rect 41083 -33852 47298 -33788
rect 47362 -33852 47382 -33788
rect 41083 -33868 47382 -33852
rect 41083 -33932 47298 -33868
rect 47362 -33932 47382 -33868
rect 41083 -33948 47382 -33932
rect 41083 -34012 47298 -33948
rect 47362 -34012 47382 -33948
rect 41083 -34028 47382 -34012
rect 41083 -34092 47298 -34028
rect 47362 -34092 47382 -34028
rect 41083 -34108 47382 -34092
rect 41083 -34172 47298 -34108
rect 47362 -34172 47382 -34108
rect 41083 -34188 47382 -34172
rect 41083 -34252 47298 -34188
rect 47362 -34252 47382 -34188
rect 41083 -34268 47382 -34252
rect 41083 -34332 47298 -34268
rect 47362 -34332 47382 -34268
rect 41083 -34348 47382 -34332
rect 41083 -34412 47298 -34348
rect 47362 -34412 47382 -34348
rect 41083 -34428 47382 -34412
rect 41083 -34492 47298 -34428
rect 47362 -34492 47382 -34428
rect 41083 -34508 47382 -34492
rect 41083 -34572 47298 -34508
rect 47362 -34572 47382 -34508
rect 41083 -34600 47382 -34572
rect -47383 -34728 -41084 -34700
rect -47383 -34792 -41168 -34728
rect -41104 -34792 -41084 -34728
rect -47383 -34808 -41084 -34792
rect -47383 -34872 -41168 -34808
rect -41104 -34872 -41084 -34808
rect -47383 -34888 -41084 -34872
rect -47383 -34952 -41168 -34888
rect -41104 -34952 -41084 -34888
rect -47383 -34968 -41084 -34952
rect -47383 -35032 -41168 -34968
rect -41104 -35032 -41084 -34968
rect -47383 -35048 -41084 -35032
rect -47383 -35112 -41168 -35048
rect -41104 -35112 -41084 -35048
rect -47383 -35128 -41084 -35112
rect -47383 -35192 -41168 -35128
rect -41104 -35192 -41084 -35128
rect -47383 -35208 -41084 -35192
rect -47383 -35272 -41168 -35208
rect -41104 -35272 -41084 -35208
rect -47383 -35288 -41084 -35272
rect -47383 -35352 -41168 -35288
rect -41104 -35352 -41084 -35288
rect -47383 -35368 -41084 -35352
rect -47383 -35432 -41168 -35368
rect -41104 -35432 -41084 -35368
rect -47383 -35448 -41084 -35432
rect -47383 -35512 -41168 -35448
rect -41104 -35512 -41084 -35448
rect -47383 -35528 -41084 -35512
rect -47383 -35592 -41168 -35528
rect -41104 -35592 -41084 -35528
rect -47383 -35608 -41084 -35592
rect -47383 -35672 -41168 -35608
rect -41104 -35672 -41084 -35608
rect -47383 -35688 -41084 -35672
rect -47383 -35752 -41168 -35688
rect -41104 -35752 -41084 -35688
rect -47383 -35768 -41084 -35752
rect -47383 -35832 -41168 -35768
rect -41104 -35832 -41084 -35768
rect -47383 -35848 -41084 -35832
rect -47383 -35912 -41168 -35848
rect -41104 -35912 -41084 -35848
rect -47383 -35928 -41084 -35912
rect -47383 -35992 -41168 -35928
rect -41104 -35992 -41084 -35928
rect -47383 -36008 -41084 -35992
rect -47383 -36072 -41168 -36008
rect -41104 -36072 -41084 -36008
rect -47383 -36088 -41084 -36072
rect -47383 -36152 -41168 -36088
rect -41104 -36152 -41084 -36088
rect -47383 -36168 -41084 -36152
rect -47383 -36232 -41168 -36168
rect -41104 -36232 -41084 -36168
rect -47383 -36248 -41084 -36232
rect -47383 -36312 -41168 -36248
rect -41104 -36312 -41084 -36248
rect -47383 -36328 -41084 -36312
rect -47383 -36392 -41168 -36328
rect -41104 -36392 -41084 -36328
rect -47383 -36408 -41084 -36392
rect -47383 -36472 -41168 -36408
rect -41104 -36472 -41084 -36408
rect -47383 -36488 -41084 -36472
rect -47383 -36552 -41168 -36488
rect -41104 -36552 -41084 -36488
rect -47383 -36568 -41084 -36552
rect -47383 -36632 -41168 -36568
rect -41104 -36632 -41084 -36568
rect -47383 -36648 -41084 -36632
rect -47383 -36712 -41168 -36648
rect -41104 -36712 -41084 -36648
rect -47383 -36728 -41084 -36712
rect -47383 -36792 -41168 -36728
rect -41104 -36792 -41084 -36728
rect -47383 -36808 -41084 -36792
rect -47383 -36872 -41168 -36808
rect -41104 -36872 -41084 -36808
rect -47383 -36888 -41084 -36872
rect -47383 -36952 -41168 -36888
rect -41104 -36952 -41084 -36888
rect -47383 -36968 -41084 -36952
rect -47383 -37032 -41168 -36968
rect -41104 -37032 -41084 -36968
rect -47383 -37048 -41084 -37032
rect -47383 -37112 -41168 -37048
rect -41104 -37112 -41084 -37048
rect -47383 -37128 -41084 -37112
rect -47383 -37192 -41168 -37128
rect -41104 -37192 -41084 -37128
rect -47383 -37208 -41084 -37192
rect -47383 -37272 -41168 -37208
rect -41104 -37272 -41084 -37208
rect -47383 -37288 -41084 -37272
rect -47383 -37352 -41168 -37288
rect -41104 -37352 -41084 -37288
rect -47383 -37368 -41084 -37352
rect -47383 -37432 -41168 -37368
rect -41104 -37432 -41084 -37368
rect -47383 -37448 -41084 -37432
rect -47383 -37512 -41168 -37448
rect -41104 -37512 -41084 -37448
rect -47383 -37528 -41084 -37512
rect -47383 -37592 -41168 -37528
rect -41104 -37592 -41084 -37528
rect -47383 -37608 -41084 -37592
rect -47383 -37672 -41168 -37608
rect -41104 -37672 -41084 -37608
rect -47383 -37688 -41084 -37672
rect -47383 -37752 -41168 -37688
rect -41104 -37752 -41084 -37688
rect -47383 -37768 -41084 -37752
rect -47383 -37832 -41168 -37768
rect -41104 -37832 -41084 -37768
rect -47383 -37848 -41084 -37832
rect -47383 -37912 -41168 -37848
rect -41104 -37912 -41084 -37848
rect -47383 -37928 -41084 -37912
rect -47383 -37992 -41168 -37928
rect -41104 -37992 -41084 -37928
rect -47383 -38008 -41084 -37992
rect -47383 -38072 -41168 -38008
rect -41104 -38072 -41084 -38008
rect -47383 -38088 -41084 -38072
rect -47383 -38152 -41168 -38088
rect -41104 -38152 -41084 -38088
rect -47383 -38168 -41084 -38152
rect -47383 -38232 -41168 -38168
rect -41104 -38232 -41084 -38168
rect -47383 -38248 -41084 -38232
rect -47383 -38312 -41168 -38248
rect -41104 -38312 -41084 -38248
rect -47383 -38328 -41084 -38312
rect -47383 -38392 -41168 -38328
rect -41104 -38392 -41084 -38328
rect -47383 -38408 -41084 -38392
rect -47383 -38472 -41168 -38408
rect -41104 -38472 -41084 -38408
rect -47383 -38488 -41084 -38472
rect -47383 -38552 -41168 -38488
rect -41104 -38552 -41084 -38488
rect -47383 -38568 -41084 -38552
rect -47383 -38632 -41168 -38568
rect -41104 -38632 -41084 -38568
rect -47383 -38648 -41084 -38632
rect -47383 -38712 -41168 -38648
rect -41104 -38712 -41084 -38648
rect -47383 -38728 -41084 -38712
rect -47383 -38792 -41168 -38728
rect -41104 -38792 -41084 -38728
rect -47383 -38808 -41084 -38792
rect -47383 -38872 -41168 -38808
rect -41104 -38872 -41084 -38808
rect -47383 -38888 -41084 -38872
rect -47383 -38952 -41168 -38888
rect -41104 -38952 -41084 -38888
rect -47383 -38968 -41084 -38952
rect -47383 -39032 -41168 -38968
rect -41104 -39032 -41084 -38968
rect -47383 -39048 -41084 -39032
rect -47383 -39112 -41168 -39048
rect -41104 -39112 -41084 -39048
rect -47383 -39128 -41084 -39112
rect -47383 -39192 -41168 -39128
rect -41104 -39192 -41084 -39128
rect -47383 -39208 -41084 -39192
rect -47383 -39272 -41168 -39208
rect -41104 -39272 -41084 -39208
rect -47383 -39288 -41084 -39272
rect -47383 -39352 -41168 -39288
rect -41104 -39352 -41084 -39288
rect -47383 -39368 -41084 -39352
rect -47383 -39432 -41168 -39368
rect -41104 -39432 -41084 -39368
rect -47383 -39448 -41084 -39432
rect -47383 -39512 -41168 -39448
rect -41104 -39512 -41084 -39448
rect -47383 -39528 -41084 -39512
rect -47383 -39592 -41168 -39528
rect -41104 -39592 -41084 -39528
rect -47383 -39608 -41084 -39592
rect -47383 -39672 -41168 -39608
rect -41104 -39672 -41084 -39608
rect -47383 -39688 -41084 -39672
rect -47383 -39752 -41168 -39688
rect -41104 -39752 -41084 -39688
rect -47383 -39768 -41084 -39752
rect -47383 -39832 -41168 -39768
rect -41104 -39832 -41084 -39768
rect -47383 -39848 -41084 -39832
rect -47383 -39912 -41168 -39848
rect -41104 -39912 -41084 -39848
rect -47383 -39928 -41084 -39912
rect -47383 -39992 -41168 -39928
rect -41104 -39992 -41084 -39928
rect -47383 -40008 -41084 -39992
rect -47383 -40072 -41168 -40008
rect -41104 -40072 -41084 -40008
rect -47383 -40088 -41084 -40072
rect -47383 -40152 -41168 -40088
rect -41104 -40152 -41084 -40088
rect -47383 -40168 -41084 -40152
rect -47383 -40232 -41168 -40168
rect -41104 -40232 -41084 -40168
rect -47383 -40248 -41084 -40232
rect -47383 -40312 -41168 -40248
rect -41104 -40312 -41084 -40248
rect -47383 -40328 -41084 -40312
rect -47383 -40392 -41168 -40328
rect -41104 -40392 -41084 -40328
rect -47383 -40408 -41084 -40392
rect -47383 -40472 -41168 -40408
rect -41104 -40472 -41084 -40408
rect -47383 -40488 -41084 -40472
rect -47383 -40552 -41168 -40488
rect -41104 -40552 -41084 -40488
rect -47383 -40568 -41084 -40552
rect -47383 -40632 -41168 -40568
rect -41104 -40632 -41084 -40568
rect -47383 -40648 -41084 -40632
rect -47383 -40712 -41168 -40648
rect -41104 -40712 -41084 -40648
rect -47383 -40728 -41084 -40712
rect -47383 -40792 -41168 -40728
rect -41104 -40792 -41084 -40728
rect -47383 -40808 -41084 -40792
rect -47383 -40872 -41168 -40808
rect -41104 -40872 -41084 -40808
rect -47383 -40900 -41084 -40872
rect -41064 -34728 -34765 -34700
rect -41064 -34792 -34849 -34728
rect -34785 -34792 -34765 -34728
rect -41064 -34808 -34765 -34792
rect -41064 -34872 -34849 -34808
rect -34785 -34872 -34765 -34808
rect -41064 -34888 -34765 -34872
rect -41064 -34952 -34849 -34888
rect -34785 -34952 -34765 -34888
rect -41064 -34968 -34765 -34952
rect -41064 -35032 -34849 -34968
rect -34785 -35032 -34765 -34968
rect -41064 -35048 -34765 -35032
rect -41064 -35112 -34849 -35048
rect -34785 -35112 -34765 -35048
rect -41064 -35128 -34765 -35112
rect -41064 -35192 -34849 -35128
rect -34785 -35192 -34765 -35128
rect -41064 -35208 -34765 -35192
rect -41064 -35272 -34849 -35208
rect -34785 -35272 -34765 -35208
rect -41064 -35288 -34765 -35272
rect -41064 -35352 -34849 -35288
rect -34785 -35352 -34765 -35288
rect -41064 -35368 -34765 -35352
rect -41064 -35432 -34849 -35368
rect -34785 -35432 -34765 -35368
rect -41064 -35448 -34765 -35432
rect -41064 -35512 -34849 -35448
rect -34785 -35512 -34765 -35448
rect -41064 -35528 -34765 -35512
rect -41064 -35592 -34849 -35528
rect -34785 -35592 -34765 -35528
rect -41064 -35608 -34765 -35592
rect -41064 -35672 -34849 -35608
rect -34785 -35672 -34765 -35608
rect -41064 -35688 -34765 -35672
rect -41064 -35752 -34849 -35688
rect -34785 -35752 -34765 -35688
rect -41064 -35768 -34765 -35752
rect -41064 -35832 -34849 -35768
rect -34785 -35832 -34765 -35768
rect -41064 -35848 -34765 -35832
rect -41064 -35912 -34849 -35848
rect -34785 -35912 -34765 -35848
rect -41064 -35928 -34765 -35912
rect -41064 -35992 -34849 -35928
rect -34785 -35992 -34765 -35928
rect -41064 -36008 -34765 -35992
rect -41064 -36072 -34849 -36008
rect -34785 -36072 -34765 -36008
rect -41064 -36088 -34765 -36072
rect -41064 -36152 -34849 -36088
rect -34785 -36152 -34765 -36088
rect -41064 -36168 -34765 -36152
rect -41064 -36232 -34849 -36168
rect -34785 -36232 -34765 -36168
rect -41064 -36248 -34765 -36232
rect -41064 -36312 -34849 -36248
rect -34785 -36312 -34765 -36248
rect -41064 -36328 -34765 -36312
rect -41064 -36392 -34849 -36328
rect -34785 -36392 -34765 -36328
rect -41064 -36408 -34765 -36392
rect -41064 -36472 -34849 -36408
rect -34785 -36472 -34765 -36408
rect -41064 -36488 -34765 -36472
rect -41064 -36552 -34849 -36488
rect -34785 -36552 -34765 -36488
rect -41064 -36568 -34765 -36552
rect -41064 -36632 -34849 -36568
rect -34785 -36632 -34765 -36568
rect -41064 -36648 -34765 -36632
rect -41064 -36712 -34849 -36648
rect -34785 -36712 -34765 -36648
rect -41064 -36728 -34765 -36712
rect -41064 -36792 -34849 -36728
rect -34785 -36792 -34765 -36728
rect -41064 -36808 -34765 -36792
rect -41064 -36872 -34849 -36808
rect -34785 -36872 -34765 -36808
rect -41064 -36888 -34765 -36872
rect -41064 -36952 -34849 -36888
rect -34785 -36952 -34765 -36888
rect -41064 -36968 -34765 -36952
rect -41064 -37032 -34849 -36968
rect -34785 -37032 -34765 -36968
rect -41064 -37048 -34765 -37032
rect -41064 -37112 -34849 -37048
rect -34785 -37112 -34765 -37048
rect -41064 -37128 -34765 -37112
rect -41064 -37192 -34849 -37128
rect -34785 -37192 -34765 -37128
rect -41064 -37208 -34765 -37192
rect -41064 -37272 -34849 -37208
rect -34785 -37272 -34765 -37208
rect -41064 -37288 -34765 -37272
rect -41064 -37352 -34849 -37288
rect -34785 -37352 -34765 -37288
rect -41064 -37368 -34765 -37352
rect -41064 -37432 -34849 -37368
rect -34785 -37432 -34765 -37368
rect -41064 -37448 -34765 -37432
rect -41064 -37512 -34849 -37448
rect -34785 -37512 -34765 -37448
rect -41064 -37528 -34765 -37512
rect -41064 -37592 -34849 -37528
rect -34785 -37592 -34765 -37528
rect -41064 -37608 -34765 -37592
rect -41064 -37672 -34849 -37608
rect -34785 -37672 -34765 -37608
rect -41064 -37688 -34765 -37672
rect -41064 -37752 -34849 -37688
rect -34785 -37752 -34765 -37688
rect -41064 -37768 -34765 -37752
rect -41064 -37832 -34849 -37768
rect -34785 -37832 -34765 -37768
rect -41064 -37848 -34765 -37832
rect -41064 -37912 -34849 -37848
rect -34785 -37912 -34765 -37848
rect -41064 -37928 -34765 -37912
rect -41064 -37992 -34849 -37928
rect -34785 -37992 -34765 -37928
rect -41064 -38008 -34765 -37992
rect -41064 -38072 -34849 -38008
rect -34785 -38072 -34765 -38008
rect -41064 -38088 -34765 -38072
rect -41064 -38152 -34849 -38088
rect -34785 -38152 -34765 -38088
rect -41064 -38168 -34765 -38152
rect -41064 -38232 -34849 -38168
rect -34785 -38232 -34765 -38168
rect -41064 -38248 -34765 -38232
rect -41064 -38312 -34849 -38248
rect -34785 -38312 -34765 -38248
rect -41064 -38328 -34765 -38312
rect -41064 -38392 -34849 -38328
rect -34785 -38392 -34765 -38328
rect -41064 -38408 -34765 -38392
rect -41064 -38472 -34849 -38408
rect -34785 -38472 -34765 -38408
rect -41064 -38488 -34765 -38472
rect -41064 -38552 -34849 -38488
rect -34785 -38552 -34765 -38488
rect -41064 -38568 -34765 -38552
rect -41064 -38632 -34849 -38568
rect -34785 -38632 -34765 -38568
rect -41064 -38648 -34765 -38632
rect -41064 -38712 -34849 -38648
rect -34785 -38712 -34765 -38648
rect -41064 -38728 -34765 -38712
rect -41064 -38792 -34849 -38728
rect -34785 -38792 -34765 -38728
rect -41064 -38808 -34765 -38792
rect -41064 -38872 -34849 -38808
rect -34785 -38872 -34765 -38808
rect -41064 -38888 -34765 -38872
rect -41064 -38952 -34849 -38888
rect -34785 -38952 -34765 -38888
rect -41064 -38968 -34765 -38952
rect -41064 -39032 -34849 -38968
rect -34785 -39032 -34765 -38968
rect -41064 -39048 -34765 -39032
rect -41064 -39112 -34849 -39048
rect -34785 -39112 -34765 -39048
rect -41064 -39128 -34765 -39112
rect -41064 -39192 -34849 -39128
rect -34785 -39192 -34765 -39128
rect -41064 -39208 -34765 -39192
rect -41064 -39272 -34849 -39208
rect -34785 -39272 -34765 -39208
rect -41064 -39288 -34765 -39272
rect -41064 -39352 -34849 -39288
rect -34785 -39352 -34765 -39288
rect -41064 -39368 -34765 -39352
rect -41064 -39432 -34849 -39368
rect -34785 -39432 -34765 -39368
rect -41064 -39448 -34765 -39432
rect -41064 -39512 -34849 -39448
rect -34785 -39512 -34765 -39448
rect -41064 -39528 -34765 -39512
rect -41064 -39592 -34849 -39528
rect -34785 -39592 -34765 -39528
rect -41064 -39608 -34765 -39592
rect -41064 -39672 -34849 -39608
rect -34785 -39672 -34765 -39608
rect -41064 -39688 -34765 -39672
rect -41064 -39752 -34849 -39688
rect -34785 -39752 -34765 -39688
rect -41064 -39768 -34765 -39752
rect -41064 -39832 -34849 -39768
rect -34785 -39832 -34765 -39768
rect -41064 -39848 -34765 -39832
rect -41064 -39912 -34849 -39848
rect -34785 -39912 -34765 -39848
rect -41064 -39928 -34765 -39912
rect -41064 -39992 -34849 -39928
rect -34785 -39992 -34765 -39928
rect -41064 -40008 -34765 -39992
rect -41064 -40072 -34849 -40008
rect -34785 -40072 -34765 -40008
rect -41064 -40088 -34765 -40072
rect -41064 -40152 -34849 -40088
rect -34785 -40152 -34765 -40088
rect -41064 -40168 -34765 -40152
rect -41064 -40232 -34849 -40168
rect -34785 -40232 -34765 -40168
rect -41064 -40248 -34765 -40232
rect -41064 -40312 -34849 -40248
rect -34785 -40312 -34765 -40248
rect -41064 -40328 -34765 -40312
rect -41064 -40392 -34849 -40328
rect -34785 -40392 -34765 -40328
rect -41064 -40408 -34765 -40392
rect -41064 -40472 -34849 -40408
rect -34785 -40472 -34765 -40408
rect -41064 -40488 -34765 -40472
rect -41064 -40552 -34849 -40488
rect -34785 -40552 -34765 -40488
rect -41064 -40568 -34765 -40552
rect -41064 -40632 -34849 -40568
rect -34785 -40632 -34765 -40568
rect -41064 -40648 -34765 -40632
rect -41064 -40712 -34849 -40648
rect -34785 -40712 -34765 -40648
rect -41064 -40728 -34765 -40712
rect -41064 -40792 -34849 -40728
rect -34785 -40792 -34765 -40728
rect -41064 -40808 -34765 -40792
rect -41064 -40872 -34849 -40808
rect -34785 -40872 -34765 -40808
rect -41064 -40900 -34765 -40872
rect -34745 -34728 -28446 -34700
rect -34745 -34792 -28530 -34728
rect -28466 -34792 -28446 -34728
rect -34745 -34808 -28446 -34792
rect -34745 -34872 -28530 -34808
rect -28466 -34872 -28446 -34808
rect -34745 -34888 -28446 -34872
rect -34745 -34952 -28530 -34888
rect -28466 -34952 -28446 -34888
rect -34745 -34968 -28446 -34952
rect -34745 -35032 -28530 -34968
rect -28466 -35032 -28446 -34968
rect -34745 -35048 -28446 -35032
rect -34745 -35112 -28530 -35048
rect -28466 -35112 -28446 -35048
rect -34745 -35128 -28446 -35112
rect -34745 -35192 -28530 -35128
rect -28466 -35192 -28446 -35128
rect -34745 -35208 -28446 -35192
rect -34745 -35272 -28530 -35208
rect -28466 -35272 -28446 -35208
rect -34745 -35288 -28446 -35272
rect -34745 -35352 -28530 -35288
rect -28466 -35352 -28446 -35288
rect -34745 -35368 -28446 -35352
rect -34745 -35432 -28530 -35368
rect -28466 -35432 -28446 -35368
rect -34745 -35448 -28446 -35432
rect -34745 -35512 -28530 -35448
rect -28466 -35512 -28446 -35448
rect -34745 -35528 -28446 -35512
rect -34745 -35592 -28530 -35528
rect -28466 -35592 -28446 -35528
rect -34745 -35608 -28446 -35592
rect -34745 -35672 -28530 -35608
rect -28466 -35672 -28446 -35608
rect -34745 -35688 -28446 -35672
rect -34745 -35752 -28530 -35688
rect -28466 -35752 -28446 -35688
rect -34745 -35768 -28446 -35752
rect -34745 -35832 -28530 -35768
rect -28466 -35832 -28446 -35768
rect -34745 -35848 -28446 -35832
rect -34745 -35912 -28530 -35848
rect -28466 -35912 -28446 -35848
rect -34745 -35928 -28446 -35912
rect -34745 -35992 -28530 -35928
rect -28466 -35992 -28446 -35928
rect -34745 -36008 -28446 -35992
rect -34745 -36072 -28530 -36008
rect -28466 -36072 -28446 -36008
rect -34745 -36088 -28446 -36072
rect -34745 -36152 -28530 -36088
rect -28466 -36152 -28446 -36088
rect -34745 -36168 -28446 -36152
rect -34745 -36232 -28530 -36168
rect -28466 -36232 -28446 -36168
rect -34745 -36248 -28446 -36232
rect -34745 -36312 -28530 -36248
rect -28466 -36312 -28446 -36248
rect -34745 -36328 -28446 -36312
rect -34745 -36392 -28530 -36328
rect -28466 -36392 -28446 -36328
rect -34745 -36408 -28446 -36392
rect -34745 -36472 -28530 -36408
rect -28466 -36472 -28446 -36408
rect -34745 -36488 -28446 -36472
rect -34745 -36552 -28530 -36488
rect -28466 -36552 -28446 -36488
rect -34745 -36568 -28446 -36552
rect -34745 -36632 -28530 -36568
rect -28466 -36632 -28446 -36568
rect -34745 -36648 -28446 -36632
rect -34745 -36712 -28530 -36648
rect -28466 -36712 -28446 -36648
rect -34745 -36728 -28446 -36712
rect -34745 -36792 -28530 -36728
rect -28466 -36792 -28446 -36728
rect -34745 -36808 -28446 -36792
rect -34745 -36872 -28530 -36808
rect -28466 -36872 -28446 -36808
rect -34745 -36888 -28446 -36872
rect -34745 -36952 -28530 -36888
rect -28466 -36952 -28446 -36888
rect -34745 -36968 -28446 -36952
rect -34745 -37032 -28530 -36968
rect -28466 -37032 -28446 -36968
rect -34745 -37048 -28446 -37032
rect -34745 -37112 -28530 -37048
rect -28466 -37112 -28446 -37048
rect -34745 -37128 -28446 -37112
rect -34745 -37192 -28530 -37128
rect -28466 -37192 -28446 -37128
rect -34745 -37208 -28446 -37192
rect -34745 -37272 -28530 -37208
rect -28466 -37272 -28446 -37208
rect -34745 -37288 -28446 -37272
rect -34745 -37352 -28530 -37288
rect -28466 -37352 -28446 -37288
rect -34745 -37368 -28446 -37352
rect -34745 -37432 -28530 -37368
rect -28466 -37432 -28446 -37368
rect -34745 -37448 -28446 -37432
rect -34745 -37512 -28530 -37448
rect -28466 -37512 -28446 -37448
rect -34745 -37528 -28446 -37512
rect -34745 -37592 -28530 -37528
rect -28466 -37592 -28446 -37528
rect -34745 -37608 -28446 -37592
rect -34745 -37672 -28530 -37608
rect -28466 -37672 -28446 -37608
rect -34745 -37688 -28446 -37672
rect -34745 -37752 -28530 -37688
rect -28466 -37752 -28446 -37688
rect -34745 -37768 -28446 -37752
rect -34745 -37832 -28530 -37768
rect -28466 -37832 -28446 -37768
rect -34745 -37848 -28446 -37832
rect -34745 -37912 -28530 -37848
rect -28466 -37912 -28446 -37848
rect -34745 -37928 -28446 -37912
rect -34745 -37992 -28530 -37928
rect -28466 -37992 -28446 -37928
rect -34745 -38008 -28446 -37992
rect -34745 -38072 -28530 -38008
rect -28466 -38072 -28446 -38008
rect -34745 -38088 -28446 -38072
rect -34745 -38152 -28530 -38088
rect -28466 -38152 -28446 -38088
rect -34745 -38168 -28446 -38152
rect -34745 -38232 -28530 -38168
rect -28466 -38232 -28446 -38168
rect -34745 -38248 -28446 -38232
rect -34745 -38312 -28530 -38248
rect -28466 -38312 -28446 -38248
rect -34745 -38328 -28446 -38312
rect -34745 -38392 -28530 -38328
rect -28466 -38392 -28446 -38328
rect -34745 -38408 -28446 -38392
rect -34745 -38472 -28530 -38408
rect -28466 -38472 -28446 -38408
rect -34745 -38488 -28446 -38472
rect -34745 -38552 -28530 -38488
rect -28466 -38552 -28446 -38488
rect -34745 -38568 -28446 -38552
rect -34745 -38632 -28530 -38568
rect -28466 -38632 -28446 -38568
rect -34745 -38648 -28446 -38632
rect -34745 -38712 -28530 -38648
rect -28466 -38712 -28446 -38648
rect -34745 -38728 -28446 -38712
rect -34745 -38792 -28530 -38728
rect -28466 -38792 -28446 -38728
rect -34745 -38808 -28446 -38792
rect -34745 -38872 -28530 -38808
rect -28466 -38872 -28446 -38808
rect -34745 -38888 -28446 -38872
rect -34745 -38952 -28530 -38888
rect -28466 -38952 -28446 -38888
rect -34745 -38968 -28446 -38952
rect -34745 -39032 -28530 -38968
rect -28466 -39032 -28446 -38968
rect -34745 -39048 -28446 -39032
rect -34745 -39112 -28530 -39048
rect -28466 -39112 -28446 -39048
rect -34745 -39128 -28446 -39112
rect -34745 -39192 -28530 -39128
rect -28466 -39192 -28446 -39128
rect -34745 -39208 -28446 -39192
rect -34745 -39272 -28530 -39208
rect -28466 -39272 -28446 -39208
rect -34745 -39288 -28446 -39272
rect -34745 -39352 -28530 -39288
rect -28466 -39352 -28446 -39288
rect -34745 -39368 -28446 -39352
rect -34745 -39432 -28530 -39368
rect -28466 -39432 -28446 -39368
rect -34745 -39448 -28446 -39432
rect -34745 -39512 -28530 -39448
rect -28466 -39512 -28446 -39448
rect -34745 -39528 -28446 -39512
rect -34745 -39592 -28530 -39528
rect -28466 -39592 -28446 -39528
rect -34745 -39608 -28446 -39592
rect -34745 -39672 -28530 -39608
rect -28466 -39672 -28446 -39608
rect -34745 -39688 -28446 -39672
rect -34745 -39752 -28530 -39688
rect -28466 -39752 -28446 -39688
rect -34745 -39768 -28446 -39752
rect -34745 -39832 -28530 -39768
rect -28466 -39832 -28446 -39768
rect -34745 -39848 -28446 -39832
rect -34745 -39912 -28530 -39848
rect -28466 -39912 -28446 -39848
rect -34745 -39928 -28446 -39912
rect -34745 -39992 -28530 -39928
rect -28466 -39992 -28446 -39928
rect -34745 -40008 -28446 -39992
rect -34745 -40072 -28530 -40008
rect -28466 -40072 -28446 -40008
rect -34745 -40088 -28446 -40072
rect -34745 -40152 -28530 -40088
rect -28466 -40152 -28446 -40088
rect -34745 -40168 -28446 -40152
rect -34745 -40232 -28530 -40168
rect -28466 -40232 -28446 -40168
rect -34745 -40248 -28446 -40232
rect -34745 -40312 -28530 -40248
rect -28466 -40312 -28446 -40248
rect -34745 -40328 -28446 -40312
rect -34745 -40392 -28530 -40328
rect -28466 -40392 -28446 -40328
rect -34745 -40408 -28446 -40392
rect -34745 -40472 -28530 -40408
rect -28466 -40472 -28446 -40408
rect -34745 -40488 -28446 -40472
rect -34745 -40552 -28530 -40488
rect -28466 -40552 -28446 -40488
rect -34745 -40568 -28446 -40552
rect -34745 -40632 -28530 -40568
rect -28466 -40632 -28446 -40568
rect -34745 -40648 -28446 -40632
rect -34745 -40712 -28530 -40648
rect -28466 -40712 -28446 -40648
rect -34745 -40728 -28446 -40712
rect -34745 -40792 -28530 -40728
rect -28466 -40792 -28446 -40728
rect -34745 -40808 -28446 -40792
rect -34745 -40872 -28530 -40808
rect -28466 -40872 -28446 -40808
rect -34745 -40900 -28446 -40872
rect -28426 -34728 -22127 -34700
rect -28426 -34792 -22211 -34728
rect -22147 -34792 -22127 -34728
rect -28426 -34808 -22127 -34792
rect -28426 -34872 -22211 -34808
rect -22147 -34872 -22127 -34808
rect -28426 -34888 -22127 -34872
rect -28426 -34952 -22211 -34888
rect -22147 -34952 -22127 -34888
rect -28426 -34968 -22127 -34952
rect -28426 -35032 -22211 -34968
rect -22147 -35032 -22127 -34968
rect -28426 -35048 -22127 -35032
rect -28426 -35112 -22211 -35048
rect -22147 -35112 -22127 -35048
rect -28426 -35128 -22127 -35112
rect -28426 -35192 -22211 -35128
rect -22147 -35192 -22127 -35128
rect -28426 -35208 -22127 -35192
rect -28426 -35272 -22211 -35208
rect -22147 -35272 -22127 -35208
rect -28426 -35288 -22127 -35272
rect -28426 -35352 -22211 -35288
rect -22147 -35352 -22127 -35288
rect -28426 -35368 -22127 -35352
rect -28426 -35432 -22211 -35368
rect -22147 -35432 -22127 -35368
rect -28426 -35448 -22127 -35432
rect -28426 -35512 -22211 -35448
rect -22147 -35512 -22127 -35448
rect -28426 -35528 -22127 -35512
rect -28426 -35592 -22211 -35528
rect -22147 -35592 -22127 -35528
rect -28426 -35608 -22127 -35592
rect -28426 -35672 -22211 -35608
rect -22147 -35672 -22127 -35608
rect -28426 -35688 -22127 -35672
rect -28426 -35752 -22211 -35688
rect -22147 -35752 -22127 -35688
rect -28426 -35768 -22127 -35752
rect -28426 -35832 -22211 -35768
rect -22147 -35832 -22127 -35768
rect -28426 -35848 -22127 -35832
rect -28426 -35912 -22211 -35848
rect -22147 -35912 -22127 -35848
rect -28426 -35928 -22127 -35912
rect -28426 -35992 -22211 -35928
rect -22147 -35992 -22127 -35928
rect -28426 -36008 -22127 -35992
rect -28426 -36072 -22211 -36008
rect -22147 -36072 -22127 -36008
rect -28426 -36088 -22127 -36072
rect -28426 -36152 -22211 -36088
rect -22147 -36152 -22127 -36088
rect -28426 -36168 -22127 -36152
rect -28426 -36232 -22211 -36168
rect -22147 -36232 -22127 -36168
rect -28426 -36248 -22127 -36232
rect -28426 -36312 -22211 -36248
rect -22147 -36312 -22127 -36248
rect -28426 -36328 -22127 -36312
rect -28426 -36392 -22211 -36328
rect -22147 -36392 -22127 -36328
rect -28426 -36408 -22127 -36392
rect -28426 -36472 -22211 -36408
rect -22147 -36472 -22127 -36408
rect -28426 -36488 -22127 -36472
rect -28426 -36552 -22211 -36488
rect -22147 -36552 -22127 -36488
rect -28426 -36568 -22127 -36552
rect -28426 -36632 -22211 -36568
rect -22147 -36632 -22127 -36568
rect -28426 -36648 -22127 -36632
rect -28426 -36712 -22211 -36648
rect -22147 -36712 -22127 -36648
rect -28426 -36728 -22127 -36712
rect -28426 -36792 -22211 -36728
rect -22147 -36792 -22127 -36728
rect -28426 -36808 -22127 -36792
rect -28426 -36872 -22211 -36808
rect -22147 -36872 -22127 -36808
rect -28426 -36888 -22127 -36872
rect -28426 -36952 -22211 -36888
rect -22147 -36952 -22127 -36888
rect -28426 -36968 -22127 -36952
rect -28426 -37032 -22211 -36968
rect -22147 -37032 -22127 -36968
rect -28426 -37048 -22127 -37032
rect -28426 -37112 -22211 -37048
rect -22147 -37112 -22127 -37048
rect -28426 -37128 -22127 -37112
rect -28426 -37192 -22211 -37128
rect -22147 -37192 -22127 -37128
rect -28426 -37208 -22127 -37192
rect -28426 -37272 -22211 -37208
rect -22147 -37272 -22127 -37208
rect -28426 -37288 -22127 -37272
rect -28426 -37352 -22211 -37288
rect -22147 -37352 -22127 -37288
rect -28426 -37368 -22127 -37352
rect -28426 -37432 -22211 -37368
rect -22147 -37432 -22127 -37368
rect -28426 -37448 -22127 -37432
rect -28426 -37512 -22211 -37448
rect -22147 -37512 -22127 -37448
rect -28426 -37528 -22127 -37512
rect -28426 -37592 -22211 -37528
rect -22147 -37592 -22127 -37528
rect -28426 -37608 -22127 -37592
rect -28426 -37672 -22211 -37608
rect -22147 -37672 -22127 -37608
rect -28426 -37688 -22127 -37672
rect -28426 -37752 -22211 -37688
rect -22147 -37752 -22127 -37688
rect -28426 -37768 -22127 -37752
rect -28426 -37832 -22211 -37768
rect -22147 -37832 -22127 -37768
rect -28426 -37848 -22127 -37832
rect -28426 -37912 -22211 -37848
rect -22147 -37912 -22127 -37848
rect -28426 -37928 -22127 -37912
rect -28426 -37992 -22211 -37928
rect -22147 -37992 -22127 -37928
rect -28426 -38008 -22127 -37992
rect -28426 -38072 -22211 -38008
rect -22147 -38072 -22127 -38008
rect -28426 -38088 -22127 -38072
rect -28426 -38152 -22211 -38088
rect -22147 -38152 -22127 -38088
rect -28426 -38168 -22127 -38152
rect -28426 -38232 -22211 -38168
rect -22147 -38232 -22127 -38168
rect -28426 -38248 -22127 -38232
rect -28426 -38312 -22211 -38248
rect -22147 -38312 -22127 -38248
rect -28426 -38328 -22127 -38312
rect -28426 -38392 -22211 -38328
rect -22147 -38392 -22127 -38328
rect -28426 -38408 -22127 -38392
rect -28426 -38472 -22211 -38408
rect -22147 -38472 -22127 -38408
rect -28426 -38488 -22127 -38472
rect -28426 -38552 -22211 -38488
rect -22147 -38552 -22127 -38488
rect -28426 -38568 -22127 -38552
rect -28426 -38632 -22211 -38568
rect -22147 -38632 -22127 -38568
rect -28426 -38648 -22127 -38632
rect -28426 -38712 -22211 -38648
rect -22147 -38712 -22127 -38648
rect -28426 -38728 -22127 -38712
rect -28426 -38792 -22211 -38728
rect -22147 -38792 -22127 -38728
rect -28426 -38808 -22127 -38792
rect -28426 -38872 -22211 -38808
rect -22147 -38872 -22127 -38808
rect -28426 -38888 -22127 -38872
rect -28426 -38952 -22211 -38888
rect -22147 -38952 -22127 -38888
rect -28426 -38968 -22127 -38952
rect -28426 -39032 -22211 -38968
rect -22147 -39032 -22127 -38968
rect -28426 -39048 -22127 -39032
rect -28426 -39112 -22211 -39048
rect -22147 -39112 -22127 -39048
rect -28426 -39128 -22127 -39112
rect -28426 -39192 -22211 -39128
rect -22147 -39192 -22127 -39128
rect -28426 -39208 -22127 -39192
rect -28426 -39272 -22211 -39208
rect -22147 -39272 -22127 -39208
rect -28426 -39288 -22127 -39272
rect -28426 -39352 -22211 -39288
rect -22147 -39352 -22127 -39288
rect -28426 -39368 -22127 -39352
rect -28426 -39432 -22211 -39368
rect -22147 -39432 -22127 -39368
rect -28426 -39448 -22127 -39432
rect -28426 -39512 -22211 -39448
rect -22147 -39512 -22127 -39448
rect -28426 -39528 -22127 -39512
rect -28426 -39592 -22211 -39528
rect -22147 -39592 -22127 -39528
rect -28426 -39608 -22127 -39592
rect -28426 -39672 -22211 -39608
rect -22147 -39672 -22127 -39608
rect -28426 -39688 -22127 -39672
rect -28426 -39752 -22211 -39688
rect -22147 -39752 -22127 -39688
rect -28426 -39768 -22127 -39752
rect -28426 -39832 -22211 -39768
rect -22147 -39832 -22127 -39768
rect -28426 -39848 -22127 -39832
rect -28426 -39912 -22211 -39848
rect -22147 -39912 -22127 -39848
rect -28426 -39928 -22127 -39912
rect -28426 -39992 -22211 -39928
rect -22147 -39992 -22127 -39928
rect -28426 -40008 -22127 -39992
rect -28426 -40072 -22211 -40008
rect -22147 -40072 -22127 -40008
rect -28426 -40088 -22127 -40072
rect -28426 -40152 -22211 -40088
rect -22147 -40152 -22127 -40088
rect -28426 -40168 -22127 -40152
rect -28426 -40232 -22211 -40168
rect -22147 -40232 -22127 -40168
rect -28426 -40248 -22127 -40232
rect -28426 -40312 -22211 -40248
rect -22147 -40312 -22127 -40248
rect -28426 -40328 -22127 -40312
rect -28426 -40392 -22211 -40328
rect -22147 -40392 -22127 -40328
rect -28426 -40408 -22127 -40392
rect -28426 -40472 -22211 -40408
rect -22147 -40472 -22127 -40408
rect -28426 -40488 -22127 -40472
rect -28426 -40552 -22211 -40488
rect -22147 -40552 -22127 -40488
rect -28426 -40568 -22127 -40552
rect -28426 -40632 -22211 -40568
rect -22147 -40632 -22127 -40568
rect -28426 -40648 -22127 -40632
rect -28426 -40712 -22211 -40648
rect -22147 -40712 -22127 -40648
rect -28426 -40728 -22127 -40712
rect -28426 -40792 -22211 -40728
rect -22147 -40792 -22127 -40728
rect -28426 -40808 -22127 -40792
rect -28426 -40872 -22211 -40808
rect -22147 -40872 -22127 -40808
rect -28426 -40900 -22127 -40872
rect -22107 -34728 -15808 -34700
rect -22107 -34792 -15892 -34728
rect -15828 -34792 -15808 -34728
rect -22107 -34808 -15808 -34792
rect -22107 -34872 -15892 -34808
rect -15828 -34872 -15808 -34808
rect -22107 -34888 -15808 -34872
rect -22107 -34952 -15892 -34888
rect -15828 -34952 -15808 -34888
rect -22107 -34968 -15808 -34952
rect -22107 -35032 -15892 -34968
rect -15828 -35032 -15808 -34968
rect -22107 -35048 -15808 -35032
rect -22107 -35112 -15892 -35048
rect -15828 -35112 -15808 -35048
rect -22107 -35128 -15808 -35112
rect -22107 -35192 -15892 -35128
rect -15828 -35192 -15808 -35128
rect -22107 -35208 -15808 -35192
rect -22107 -35272 -15892 -35208
rect -15828 -35272 -15808 -35208
rect -22107 -35288 -15808 -35272
rect -22107 -35352 -15892 -35288
rect -15828 -35352 -15808 -35288
rect -22107 -35368 -15808 -35352
rect -22107 -35432 -15892 -35368
rect -15828 -35432 -15808 -35368
rect -22107 -35448 -15808 -35432
rect -22107 -35512 -15892 -35448
rect -15828 -35512 -15808 -35448
rect -22107 -35528 -15808 -35512
rect -22107 -35592 -15892 -35528
rect -15828 -35592 -15808 -35528
rect -22107 -35608 -15808 -35592
rect -22107 -35672 -15892 -35608
rect -15828 -35672 -15808 -35608
rect -22107 -35688 -15808 -35672
rect -22107 -35752 -15892 -35688
rect -15828 -35752 -15808 -35688
rect -22107 -35768 -15808 -35752
rect -22107 -35832 -15892 -35768
rect -15828 -35832 -15808 -35768
rect -22107 -35848 -15808 -35832
rect -22107 -35912 -15892 -35848
rect -15828 -35912 -15808 -35848
rect -22107 -35928 -15808 -35912
rect -22107 -35992 -15892 -35928
rect -15828 -35992 -15808 -35928
rect -22107 -36008 -15808 -35992
rect -22107 -36072 -15892 -36008
rect -15828 -36072 -15808 -36008
rect -22107 -36088 -15808 -36072
rect -22107 -36152 -15892 -36088
rect -15828 -36152 -15808 -36088
rect -22107 -36168 -15808 -36152
rect -22107 -36232 -15892 -36168
rect -15828 -36232 -15808 -36168
rect -22107 -36248 -15808 -36232
rect -22107 -36312 -15892 -36248
rect -15828 -36312 -15808 -36248
rect -22107 -36328 -15808 -36312
rect -22107 -36392 -15892 -36328
rect -15828 -36392 -15808 -36328
rect -22107 -36408 -15808 -36392
rect -22107 -36472 -15892 -36408
rect -15828 -36472 -15808 -36408
rect -22107 -36488 -15808 -36472
rect -22107 -36552 -15892 -36488
rect -15828 -36552 -15808 -36488
rect -22107 -36568 -15808 -36552
rect -22107 -36632 -15892 -36568
rect -15828 -36632 -15808 -36568
rect -22107 -36648 -15808 -36632
rect -22107 -36712 -15892 -36648
rect -15828 -36712 -15808 -36648
rect -22107 -36728 -15808 -36712
rect -22107 -36792 -15892 -36728
rect -15828 -36792 -15808 -36728
rect -22107 -36808 -15808 -36792
rect -22107 -36872 -15892 -36808
rect -15828 -36872 -15808 -36808
rect -22107 -36888 -15808 -36872
rect -22107 -36952 -15892 -36888
rect -15828 -36952 -15808 -36888
rect -22107 -36968 -15808 -36952
rect -22107 -37032 -15892 -36968
rect -15828 -37032 -15808 -36968
rect -22107 -37048 -15808 -37032
rect -22107 -37112 -15892 -37048
rect -15828 -37112 -15808 -37048
rect -22107 -37128 -15808 -37112
rect -22107 -37192 -15892 -37128
rect -15828 -37192 -15808 -37128
rect -22107 -37208 -15808 -37192
rect -22107 -37272 -15892 -37208
rect -15828 -37272 -15808 -37208
rect -22107 -37288 -15808 -37272
rect -22107 -37352 -15892 -37288
rect -15828 -37352 -15808 -37288
rect -22107 -37368 -15808 -37352
rect -22107 -37432 -15892 -37368
rect -15828 -37432 -15808 -37368
rect -22107 -37448 -15808 -37432
rect -22107 -37512 -15892 -37448
rect -15828 -37512 -15808 -37448
rect -22107 -37528 -15808 -37512
rect -22107 -37592 -15892 -37528
rect -15828 -37592 -15808 -37528
rect -22107 -37608 -15808 -37592
rect -22107 -37672 -15892 -37608
rect -15828 -37672 -15808 -37608
rect -22107 -37688 -15808 -37672
rect -22107 -37752 -15892 -37688
rect -15828 -37752 -15808 -37688
rect -22107 -37768 -15808 -37752
rect -22107 -37832 -15892 -37768
rect -15828 -37832 -15808 -37768
rect -22107 -37848 -15808 -37832
rect -22107 -37912 -15892 -37848
rect -15828 -37912 -15808 -37848
rect -22107 -37928 -15808 -37912
rect -22107 -37992 -15892 -37928
rect -15828 -37992 -15808 -37928
rect -22107 -38008 -15808 -37992
rect -22107 -38072 -15892 -38008
rect -15828 -38072 -15808 -38008
rect -22107 -38088 -15808 -38072
rect -22107 -38152 -15892 -38088
rect -15828 -38152 -15808 -38088
rect -22107 -38168 -15808 -38152
rect -22107 -38232 -15892 -38168
rect -15828 -38232 -15808 -38168
rect -22107 -38248 -15808 -38232
rect -22107 -38312 -15892 -38248
rect -15828 -38312 -15808 -38248
rect -22107 -38328 -15808 -38312
rect -22107 -38392 -15892 -38328
rect -15828 -38392 -15808 -38328
rect -22107 -38408 -15808 -38392
rect -22107 -38472 -15892 -38408
rect -15828 -38472 -15808 -38408
rect -22107 -38488 -15808 -38472
rect -22107 -38552 -15892 -38488
rect -15828 -38552 -15808 -38488
rect -22107 -38568 -15808 -38552
rect -22107 -38632 -15892 -38568
rect -15828 -38632 -15808 -38568
rect -22107 -38648 -15808 -38632
rect -22107 -38712 -15892 -38648
rect -15828 -38712 -15808 -38648
rect -22107 -38728 -15808 -38712
rect -22107 -38792 -15892 -38728
rect -15828 -38792 -15808 -38728
rect -22107 -38808 -15808 -38792
rect -22107 -38872 -15892 -38808
rect -15828 -38872 -15808 -38808
rect -22107 -38888 -15808 -38872
rect -22107 -38952 -15892 -38888
rect -15828 -38952 -15808 -38888
rect -22107 -38968 -15808 -38952
rect -22107 -39032 -15892 -38968
rect -15828 -39032 -15808 -38968
rect -22107 -39048 -15808 -39032
rect -22107 -39112 -15892 -39048
rect -15828 -39112 -15808 -39048
rect -22107 -39128 -15808 -39112
rect -22107 -39192 -15892 -39128
rect -15828 -39192 -15808 -39128
rect -22107 -39208 -15808 -39192
rect -22107 -39272 -15892 -39208
rect -15828 -39272 -15808 -39208
rect -22107 -39288 -15808 -39272
rect -22107 -39352 -15892 -39288
rect -15828 -39352 -15808 -39288
rect -22107 -39368 -15808 -39352
rect -22107 -39432 -15892 -39368
rect -15828 -39432 -15808 -39368
rect -22107 -39448 -15808 -39432
rect -22107 -39512 -15892 -39448
rect -15828 -39512 -15808 -39448
rect -22107 -39528 -15808 -39512
rect -22107 -39592 -15892 -39528
rect -15828 -39592 -15808 -39528
rect -22107 -39608 -15808 -39592
rect -22107 -39672 -15892 -39608
rect -15828 -39672 -15808 -39608
rect -22107 -39688 -15808 -39672
rect -22107 -39752 -15892 -39688
rect -15828 -39752 -15808 -39688
rect -22107 -39768 -15808 -39752
rect -22107 -39832 -15892 -39768
rect -15828 -39832 -15808 -39768
rect -22107 -39848 -15808 -39832
rect -22107 -39912 -15892 -39848
rect -15828 -39912 -15808 -39848
rect -22107 -39928 -15808 -39912
rect -22107 -39992 -15892 -39928
rect -15828 -39992 -15808 -39928
rect -22107 -40008 -15808 -39992
rect -22107 -40072 -15892 -40008
rect -15828 -40072 -15808 -40008
rect -22107 -40088 -15808 -40072
rect -22107 -40152 -15892 -40088
rect -15828 -40152 -15808 -40088
rect -22107 -40168 -15808 -40152
rect -22107 -40232 -15892 -40168
rect -15828 -40232 -15808 -40168
rect -22107 -40248 -15808 -40232
rect -22107 -40312 -15892 -40248
rect -15828 -40312 -15808 -40248
rect -22107 -40328 -15808 -40312
rect -22107 -40392 -15892 -40328
rect -15828 -40392 -15808 -40328
rect -22107 -40408 -15808 -40392
rect -22107 -40472 -15892 -40408
rect -15828 -40472 -15808 -40408
rect -22107 -40488 -15808 -40472
rect -22107 -40552 -15892 -40488
rect -15828 -40552 -15808 -40488
rect -22107 -40568 -15808 -40552
rect -22107 -40632 -15892 -40568
rect -15828 -40632 -15808 -40568
rect -22107 -40648 -15808 -40632
rect -22107 -40712 -15892 -40648
rect -15828 -40712 -15808 -40648
rect -22107 -40728 -15808 -40712
rect -22107 -40792 -15892 -40728
rect -15828 -40792 -15808 -40728
rect -22107 -40808 -15808 -40792
rect -22107 -40872 -15892 -40808
rect -15828 -40872 -15808 -40808
rect -22107 -40900 -15808 -40872
rect -15788 -34728 -9489 -34700
rect -15788 -34792 -9573 -34728
rect -9509 -34792 -9489 -34728
rect -15788 -34808 -9489 -34792
rect -15788 -34872 -9573 -34808
rect -9509 -34872 -9489 -34808
rect -15788 -34888 -9489 -34872
rect -15788 -34952 -9573 -34888
rect -9509 -34952 -9489 -34888
rect -15788 -34968 -9489 -34952
rect -15788 -35032 -9573 -34968
rect -9509 -35032 -9489 -34968
rect -15788 -35048 -9489 -35032
rect -15788 -35112 -9573 -35048
rect -9509 -35112 -9489 -35048
rect -15788 -35128 -9489 -35112
rect -15788 -35192 -9573 -35128
rect -9509 -35192 -9489 -35128
rect -15788 -35208 -9489 -35192
rect -15788 -35272 -9573 -35208
rect -9509 -35272 -9489 -35208
rect -15788 -35288 -9489 -35272
rect -15788 -35352 -9573 -35288
rect -9509 -35352 -9489 -35288
rect -15788 -35368 -9489 -35352
rect -15788 -35432 -9573 -35368
rect -9509 -35432 -9489 -35368
rect -15788 -35448 -9489 -35432
rect -15788 -35512 -9573 -35448
rect -9509 -35512 -9489 -35448
rect -15788 -35528 -9489 -35512
rect -15788 -35592 -9573 -35528
rect -9509 -35592 -9489 -35528
rect -15788 -35608 -9489 -35592
rect -15788 -35672 -9573 -35608
rect -9509 -35672 -9489 -35608
rect -15788 -35688 -9489 -35672
rect -15788 -35752 -9573 -35688
rect -9509 -35752 -9489 -35688
rect -15788 -35768 -9489 -35752
rect -15788 -35832 -9573 -35768
rect -9509 -35832 -9489 -35768
rect -15788 -35848 -9489 -35832
rect -15788 -35912 -9573 -35848
rect -9509 -35912 -9489 -35848
rect -15788 -35928 -9489 -35912
rect -15788 -35992 -9573 -35928
rect -9509 -35992 -9489 -35928
rect -15788 -36008 -9489 -35992
rect -15788 -36072 -9573 -36008
rect -9509 -36072 -9489 -36008
rect -15788 -36088 -9489 -36072
rect -15788 -36152 -9573 -36088
rect -9509 -36152 -9489 -36088
rect -15788 -36168 -9489 -36152
rect -15788 -36232 -9573 -36168
rect -9509 -36232 -9489 -36168
rect -15788 -36248 -9489 -36232
rect -15788 -36312 -9573 -36248
rect -9509 -36312 -9489 -36248
rect -15788 -36328 -9489 -36312
rect -15788 -36392 -9573 -36328
rect -9509 -36392 -9489 -36328
rect -15788 -36408 -9489 -36392
rect -15788 -36472 -9573 -36408
rect -9509 -36472 -9489 -36408
rect -15788 -36488 -9489 -36472
rect -15788 -36552 -9573 -36488
rect -9509 -36552 -9489 -36488
rect -15788 -36568 -9489 -36552
rect -15788 -36632 -9573 -36568
rect -9509 -36632 -9489 -36568
rect -15788 -36648 -9489 -36632
rect -15788 -36712 -9573 -36648
rect -9509 -36712 -9489 -36648
rect -15788 -36728 -9489 -36712
rect -15788 -36792 -9573 -36728
rect -9509 -36792 -9489 -36728
rect -15788 -36808 -9489 -36792
rect -15788 -36872 -9573 -36808
rect -9509 -36872 -9489 -36808
rect -15788 -36888 -9489 -36872
rect -15788 -36952 -9573 -36888
rect -9509 -36952 -9489 -36888
rect -15788 -36968 -9489 -36952
rect -15788 -37032 -9573 -36968
rect -9509 -37032 -9489 -36968
rect -15788 -37048 -9489 -37032
rect -15788 -37112 -9573 -37048
rect -9509 -37112 -9489 -37048
rect -15788 -37128 -9489 -37112
rect -15788 -37192 -9573 -37128
rect -9509 -37192 -9489 -37128
rect -15788 -37208 -9489 -37192
rect -15788 -37272 -9573 -37208
rect -9509 -37272 -9489 -37208
rect -15788 -37288 -9489 -37272
rect -15788 -37352 -9573 -37288
rect -9509 -37352 -9489 -37288
rect -15788 -37368 -9489 -37352
rect -15788 -37432 -9573 -37368
rect -9509 -37432 -9489 -37368
rect -15788 -37448 -9489 -37432
rect -15788 -37512 -9573 -37448
rect -9509 -37512 -9489 -37448
rect -15788 -37528 -9489 -37512
rect -15788 -37592 -9573 -37528
rect -9509 -37592 -9489 -37528
rect -15788 -37608 -9489 -37592
rect -15788 -37672 -9573 -37608
rect -9509 -37672 -9489 -37608
rect -15788 -37688 -9489 -37672
rect -15788 -37752 -9573 -37688
rect -9509 -37752 -9489 -37688
rect -15788 -37768 -9489 -37752
rect -15788 -37832 -9573 -37768
rect -9509 -37832 -9489 -37768
rect -15788 -37848 -9489 -37832
rect -15788 -37912 -9573 -37848
rect -9509 -37912 -9489 -37848
rect -15788 -37928 -9489 -37912
rect -15788 -37992 -9573 -37928
rect -9509 -37992 -9489 -37928
rect -15788 -38008 -9489 -37992
rect -15788 -38072 -9573 -38008
rect -9509 -38072 -9489 -38008
rect -15788 -38088 -9489 -38072
rect -15788 -38152 -9573 -38088
rect -9509 -38152 -9489 -38088
rect -15788 -38168 -9489 -38152
rect -15788 -38232 -9573 -38168
rect -9509 -38232 -9489 -38168
rect -15788 -38248 -9489 -38232
rect -15788 -38312 -9573 -38248
rect -9509 -38312 -9489 -38248
rect -15788 -38328 -9489 -38312
rect -15788 -38392 -9573 -38328
rect -9509 -38392 -9489 -38328
rect -15788 -38408 -9489 -38392
rect -15788 -38472 -9573 -38408
rect -9509 -38472 -9489 -38408
rect -15788 -38488 -9489 -38472
rect -15788 -38552 -9573 -38488
rect -9509 -38552 -9489 -38488
rect -15788 -38568 -9489 -38552
rect -15788 -38632 -9573 -38568
rect -9509 -38632 -9489 -38568
rect -15788 -38648 -9489 -38632
rect -15788 -38712 -9573 -38648
rect -9509 -38712 -9489 -38648
rect -15788 -38728 -9489 -38712
rect -15788 -38792 -9573 -38728
rect -9509 -38792 -9489 -38728
rect -15788 -38808 -9489 -38792
rect -15788 -38872 -9573 -38808
rect -9509 -38872 -9489 -38808
rect -15788 -38888 -9489 -38872
rect -15788 -38952 -9573 -38888
rect -9509 -38952 -9489 -38888
rect -15788 -38968 -9489 -38952
rect -15788 -39032 -9573 -38968
rect -9509 -39032 -9489 -38968
rect -15788 -39048 -9489 -39032
rect -15788 -39112 -9573 -39048
rect -9509 -39112 -9489 -39048
rect -15788 -39128 -9489 -39112
rect -15788 -39192 -9573 -39128
rect -9509 -39192 -9489 -39128
rect -15788 -39208 -9489 -39192
rect -15788 -39272 -9573 -39208
rect -9509 -39272 -9489 -39208
rect -15788 -39288 -9489 -39272
rect -15788 -39352 -9573 -39288
rect -9509 -39352 -9489 -39288
rect -15788 -39368 -9489 -39352
rect -15788 -39432 -9573 -39368
rect -9509 -39432 -9489 -39368
rect -15788 -39448 -9489 -39432
rect -15788 -39512 -9573 -39448
rect -9509 -39512 -9489 -39448
rect -15788 -39528 -9489 -39512
rect -15788 -39592 -9573 -39528
rect -9509 -39592 -9489 -39528
rect -15788 -39608 -9489 -39592
rect -15788 -39672 -9573 -39608
rect -9509 -39672 -9489 -39608
rect -15788 -39688 -9489 -39672
rect -15788 -39752 -9573 -39688
rect -9509 -39752 -9489 -39688
rect -15788 -39768 -9489 -39752
rect -15788 -39832 -9573 -39768
rect -9509 -39832 -9489 -39768
rect -15788 -39848 -9489 -39832
rect -15788 -39912 -9573 -39848
rect -9509 -39912 -9489 -39848
rect -15788 -39928 -9489 -39912
rect -15788 -39992 -9573 -39928
rect -9509 -39992 -9489 -39928
rect -15788 -40008 -9489 -39992
rect -15788 -40072 -9573 -40008
rect -9509 -40072 -9489 -40008
rect -15788 -40088 -9489 -40072
rect -15788 -40152 -9573 -40088
rect -9509 -40152 -9489 -40088
rect -15788 -40168 -9489 -40152
rect -15788 -40232 -9573 -40168
rect -9509 -40232 -9489 -40168
rect -15788 -40248 -9489 -40232
rect -15788 -40312 -9573 -40248
rect -9509 -40312 -9489 -40248
rect -15788 -40328 -9489 -40312
rect -15788 -40392 -9573 -40328
rect -9509 -40392 -9489 -40328
rect -15788 -40408 -9489 -40392
rect -15788 -40472 -9573 -40408
rect -9509 -40472 -9489 -40408
rect -15788 -40488 -9489 -40472
rect -15788 -40552 -9573 -40488
rect -9509 -40552 -9489 -40488
rect -15788 -40568 -9489 -40552
rect -15788 -40632 -9573 -40568
rect -9509 -40632 -9489 -40568
rect -15788 -40648 -9489 -40632
rect -15788 -40712 -9573 -40648
rect -9509 -40712 -9489 -40648
rect -15788 -40728 -9489 -40712
rect -15788 -40792 -9573 -40728
rect -9509 -40792 -9489 -40728
rect -15788 -40808 -9489 -40792
rect -15788 -40872 -9573 -40808
rect -9509 -40872 -9489 -40808
rect -15788 -40900 -9489 -40872
rect -9469 -34728 -3170 -34700
rect -9469 -34792 -3254 -34728
rect -3190 -34792 -3170 -34728
rect -9469 -34808 -3170 -34792
rect -9469 -34872 -3254 -34808
rect -3190 -34872 -3170 -34808
rect -9469 -34888 -3170 -34872
rect -9469 -34952 -3254 -34888
rect -3190 -34952 -3170 -34888
rect -9469 -34968 -3170 -34952
rect -9469 -35032 -3254 -34968
rect -3190 -35032 -3170 -34968
rect -9469 -35048 -3170 -35032
rect -9469 -35112 -3254 -35048
rect -3190 -35112 -3170 -35048
rect -9469 -35128 -3170 -35112
rect -9469 -35192 -3254 -35128
rect -3190 -35192 -3170 -35128
rect -9469 -35208 -3170 -35192
rect -9469 -35272 -3254 -35208
rect -3190 -35272 -3170 -35208
rect -9469 -35288 -3170 -35272
rect -9469 -35352 -3254 -35288
rect -3190 -35352 -3170 -35288
rect -9469 -35368 -3170 -35352
rect -9469 -35432 -3254 -35368
rect -3190 -35432 -3170 -35368
rect -9469 -35448 -3170 -35432
rect -9469 -35512 -3254 -35448
rect -3190 -35512 -3170 -35448
rect -9469 -35528 -3170 -35512
rect -9469 -35592 -3254 -35528
rect -3190 -35592 -3170 -35528
rect -9469 -35608 -3170 -35592
rect -9469 -35672 -3254 -35608
rect -3190 -35672 -3170 -35608
rect -9469 -35688 -3170 -35672
rect -9469 -35752 -3254 -35688
rect -3190 -35752 -3170 -35688
rect -9469 -35768 -3170 -35752
rect -9469 -35832 -3254 -35768
rect -3190 -35832 -3170 -35768
rect -9469 -35848 -3170 -35832
rect -9469 -35912 -3254 -35848
rect -3190 -35912 -3170 -35848
rect -9469 -35928 -3170 -35912
rect -9469 -35992 -3254 -35928
rect -3190 -35992 -3170 -35928
rect -9469 -36008 -3170 -35992
rect -9469 -36072 -3254 -36008
rect -3190 -36072 -3170 -36008
rect -9469 -36088 -3170 -36072
rect -9469 -36152 -3254 -36088
rect -3190 -36152 -3170 -36088
rect -9469 -36168 -3170 -36152
rect -9469 -36232 -3254 -36168
rect -3190 -36232 -3170 -36168
rect -9469 -36248 -3170 -36232
rect -9469 -36312 -3254 -36248
rect -3190 -36312 -3170 -36248
rect -9469 -36328 -3170 -36312
rect -9469 -36392 -3254 -36328
rect -3190 -36392 -3170 -36328
rect -9469 -36408 -3170 -36392
rect -9469 -36472 -3254 -36408
rect -3190 -36472 -3170 -36408
rect -9469 -36488 -3170 -36472
rect -9469 -36552 -3254 -36488
rect -3190 -36552 -3170 -36488
rect -9469 -36568 -3170 -36552
rect -9469 -36632 -3254 -36568
rect -3190 -36632 -3170 -36568
rect -9469 -36648 -3170 -36632
rect -9469 -36712 -3254 -36648
rect -3190 -36712 -3170 -36648
rect -9469 -36728 -3170 -36712
rect -9469 -36792 -3254 -36728
rect -3190 -36792 -3170 -36728
rect -9469 -36808 -3170 -36792
rect -9469 -36872 -3254 -36808
rect -3190 -36872 -3170 -36808
rect -9469 -36888 -3170 -36872
rect -9469 -36952 -3254 -36888
rect -3190 -36952 -3170 -36888
rect -9469 -36968 -3170 -36952
rect -9469 -37032 -3254 -36968
rect -3190 -37032 -3170 -36968
rect -9469 -37048 -3170 -37032
rect -9469 -37112 -3254 -37048
rect -3190 -37112 -3170 -37048
rect -9469 -37128 -3170 -37112
rect -9469 -37192 -3254 -37128
rect -3190 -37192 -3170 -37128
rect -9469 -37208 -3170 -37192
rect -9469 -37272 -3254 -37208
rect -3190 -37272 -3170 -37208
rect -9469 -37288 -3170 -37272
rect -9469 -37352 -3254 -37288
rect -3190 -37352 -3170 -37288
rect -9469 -37368 -3170 -37352
rect -9469 -37432 -3254 -37368
rect -3190 -37432 -3170 -37368
rect -9469 -37448 -3170 -37432
rect -9469 -37512 -3254 -37448
rect -3190 -37512 -3170 -37448
rect -9469 -37528 -3170 -37512
rect -9469 -37592 -3254 -37528
rect -3190 -37592 -3170 -37528
rect -9469 -37608 -3170 -37592
rect -9469 -37672 -3254 -37608
rect -3190 -37672 -3170 -37608
rect -9469 -37688 -3170 -37672
rect -9469 -37752 -3254 -37688
rect -3190 -37752 -3170 -37688
rect -9469 -37768 -3170 -37752
rect -9469 -37832 -3254 -37768
rect -3190 -37832 -3170 -37768
rect -9469 -37848 -3170 -37832
rect -9469 -37912 -3254 -37848
rect -3190 -37912 -3170 -37848
rect -9469 -37928 -3170 -37912
rect -9469 -37992 -3254 -37928
rect -3190 -37992 -3170 -37928
rect -9469 -38008 -3170 -37992
rect -9469 -38072 -3254 -38008
rect -3190 -38072 -3170 -38008
rect -9469 -38088 -3170 -38072
rect -9469 -38152 -3254 -38088
rect -3190 -38152 -3170 -38088
rect -9469 -38168 -3170 -38152
rect -9469 -38232 -3254 -38168
rect -3190 -38232 -3170 -38168
rect -9469 -38248 -3170 -38232
rect -9469 -38312 -3254 -38248
rect -3190 -38312 -3170 -38248
rect -9469 -38328 -3170 -38312
rect -9469 -38392 -3254 -38328
rect -3190 -38392 -3170 -38328
rect -9469 -38408 -3170 -38392
rect -9469 -38472 -3254 -38408
rect -3190 -38472 -3170 -38408
rect -9469 -38488 -3170 -38472
rect -9469 -38552 -3254 -38488
rect -3190 -38552 -3170 -38488
rect -9469 -38568 -3170 -38552
rect -9469 -38632 -3254 -38568
rect -3190 -38632 -3170 -38568
rect -9469 -38648 -3170 -38632
rect -9469 -38712 -3254 -38648
rect -3190 -38712 -3170 -38648
rect -9469 -38728 -3170 -38712
rect -9469 -38792 -3254 -38728
rect -3190 -38792 -3170 -38728
rect -9469 -38808 -3170 -38792
rect -9469 -38872 -3254 -38808
rect -3190 -38872 -3170 -38808
rect -9469 -38888 -3170 -38872
rect -9469 -38952 -3254 -38888
rect -3190 -38952 -3170 -38888
rect -9469 -38968 -3170 -38952
rect -9469 -39032 -3254 -38968
rect -3190 -39032 -3170 -38968
rect -9469 -39048 -3170 -39032
rect -9469 -39112 -3254 -39048
rect -3190 -39112 -3170 -39048
rect -9469 -39128 -3170 -39112
rect -9469 -39192 -3254 -39128
rect -3190 -39192 -3170 -39128
rect -9469 -39208 -3170 -39192
rect -9469 -39272 -3254 -39208
rect -3190 -39272 -3170 -39208
rect -9469 -39288 -3170 -39272
rect -9469 -39352 -3254 -39288
rect -3190 -39352 -3170 -39288
rect -9469 -39368 -3170 -39352
rect -9469 -39432 -3254 -39368
rect -3190 -39432 -3170 -39368
rect -9469 -39448 -3170 -39432
rect -9469 -39512 -3254 -39448
rect -3190 -39512 -3170 -39448
rect -9469 -39528 -3170 -39512
rect -9469 -39592 -3254 -39528
rect -3190 -39592 -3170 -39528
rect -9469 -39608 -3170 -39592
rect -9469 -39672 -3254 -39608
rect -3190 -39672 -3170 -39608
rect -9469 -39688 -3170 -39672
rect -9469 -39752 -3254 -39688
rect -3190 -39752 -3170 -39688
rect -9469 -39768 -3170 -39752
rect -9469 -39832 -3254 -39768
rect -3190 -39832 -3170 -39768
rect -9469 -39848 -3170 -39832
rect -9469 -39912 -3254 -39848
rect -3190 -39912 -3170 -39848
rect -9469 -39928 -3170 -39912
rect -9469 -39992 -3254 -39928
rect -3190 -39992 -3170 -39928
rect -9469 -40008 -3170 -39992
rect -9469 -40072 -3254 -40008
rect -3190 -40072 -3170 -40008
rect -9469 -40088 -3170 -40072
rect -9469 -40152 -3254 -40088
rect -3190 -40152 -3170 -40088
rect -9469 -40168 -3170 -40152
rect -9469 -40232 -3254 -40168
rect -3190 -40232 -3170 -40168
rect -9469 -40248 -3170 -40232
rect -9469 -40312 -3254 -40248
rect -3190 -40312 -3170 -40248
rect -9469 -40328 -3170 -40312
rect -9469 -40392 -3254 -40328
rect -3190 -40392 -3170 -40328
rect -9469 -40408 -3170 -40392
rect -9469 -40472 -3254 -40408
rect -3190 -40472 -3170 -40408
rect -9469 -40488 -3170 -40472
rect -9469 -40552 -3254 -40488
rect -3190 -40552 -3170 -40488
rect -9469 -40568 -3170 -40552
rect -9469 -40632 -3254 -40568
rect -3190 -40632 -3170 -40568
rect -9469 -40648 -3170 -40632
rect -9469 -40712 -3254 -40648
rect -3190 -40712 -3170 -40648
rect -9469 -40728 -3170 -40712
rect -9469 -40792 -3254 -40728
rect -3190 -40792 -3170 -40728
rect -9469 -40808 -3170 -40792
rect -9469 -40872 -3254 -40808
rect -3190 -40872 -3170 -40808
rect -9469 -40900 -3170 -40872
rect -3150 -34728 3149 -34700
rect -3150 -34792 3065 -34728
rect 3129 -34792 3149 -34728
rect -3150 -34808 3149 -34792
rect -3150 -34872 3065 -34808
rect 3129 -34872 3149 -34808
rect -3150 -34888 3149 -34872
rect -3150 -34952 3065 -34888
rect 3129 -34952 3149 -34888
rect -3150 -34968 3149 -34952
rect -3150 -35032 3065 -34968
rect 3129 -35032 3149 -34968
rect -3150 -35048 3149 -35032
rect -3150 -35112 3065 -35048
rect 3129 -35112 3149 -35048
rect -3150 -35128 3149 -35112
rect -3150 -35192 3065 -35128
rect 3129 -35192 3149 -35128
rect -3150 -35208 3149 -35192
rect -3150 -35272 3065 -35208
rect 3129 -35272 3149 -35208
rect -3150 -35288 3149 -35272
rect -3150 -35352 3065 -35288
rect 3129 -35352 3149 -35288
rect -3150 -35368 3149 -35352
rect -3150 -35432 3065 -35368
rect 3129 -35432 3149 -35368
rect -3150 -35448 3149 -35432
rect -3150 -35512 3065 -35448
rect 3129 -35512 3149 -35448
rect -3150 -35528 3149 -35512
rect -3150 -35592 3065 -35528
rect 3129 -35592 3149 -35528
rect -3150 -35608 3149 -35592
rect -3150 -35672 3065 -35608
rect 3129 -35672 3149 -35608
rect -3150 -35688 3149 -35672
rect -3150 -35752 3065 -35688
rect 3129 -35752 3149 -35688
rect -3150 -35768 3149 -35752
rect -3150 -35832 3065 -35768
rect 3129 -35832 3149 -35768
rect -3150 -35848 3149 -35832
rect -3150 -35912 3065 -35848
rect 3129 -35912 3149 -35848
rect -3150 -35928 3149 -35912
rect -3150 -35992 3065 -35928
rect 3129 -35992 3149 -35928
rect -3150 -36008 3149 -35992
rect -3150 -36072 3065 -36008
rect 3129 -36072 3149 -36008
rect -3150 -36088 3149 -36072
rect -3150 -36152 3065 -36088
rect 3129 -36152 3149 -36088
rect -3150 -36168 3149 -36152
rect -3150 -36232 3065 -36168
rect 3129 -36232 3149 -36168
rect -3150 -36248 3149 -36232
rect -3150 -36312 3065 -36248
rect 3129 -36312 3149 -36248
rect -3150 -36328 3149 -36312
rect -3150 -36392 3065 -36328
rect 3129 -36392 3149 -36328
rect -3150 -36408 3149 -36392
rect -3150 -36472 3065 -36408
rect 3129 -36472 3149 -36408
rect -3150 -36488 3149 -36472
rect -3150 -36552 3065 -36488
rect 3129 -36552 3149 -36488
rect -3150 -36568 3149 -36552
rect -3150 -36632 3065 -36568
rect 3129 -36632 3149 -36568
rect -3150 -36648 3149 -36632
rect -3150 -36712 3065 -36648
rect 3129 -36712 3149 -36648
rect -3150 -36728 3149 -36712
rect -3150 -36792 3065 -36728
rect 3129 -36792 3149 -36728
rect -3150 -36808 3149 -36792
rect -3150 -36872 3065 -36808
rect 3129 -36872 3149 -36808
rect -3150 -36888 3149 -36872
rect -3150 -36952 3065 -36888
rect 3129 -36952 3149 -36888
rect -3150 -36968 3149 -36952
rect -3150 -37032 3065 -36968
rect 3129 -37032 3149 -36968
rect -3150 -37048 3149 -37032
rect -3150 -37112 3065 -37048
rect 3129 -37112 3149 -37048
rect -3150 -37128 3149 -37112
rect -3150 -37192 3065 -37128
rect 3129 -37192 3149 -37128
rect -3150 -37208 3149 -37192
rect -3150 -37272 3065 -37208
rect 3129 -37272 3149 -37208
rect -3150 -37288 3149 -37272
rect -3150 -37352 3065 -37288
rect 3129 -37352 3149 -37288
rect -3150 -37368 3149 -37352
rect -3150 -37432 3065 -37368
rect 3129 -37432 3149 -37368
rect -3150 -37448 3149 -37432
rect -3150 -37512 3065 -37448
rect 3129 -37512 3149 -37448
rect -3150 -37528 3149 -37512
rect -3150 -37592 3065 -37528
rect 3129 -37592 3149 -37528
rect -3150 -37608 3149 -37592
rect -3150 -37672 3065 -37608
rect 3129 -37672 3149 -37608
rect -3150 -37688 3149 -37672
rect -3150 -37752 3065 -37688
rect 3129 -37752 3149 -37688
rect -3150 -37768 3149 -37752
rect -3150 -37832 3065 -37768
rect 3129 -37832 3149 -37768
rect -3150 -37848 3149 -37832
rect -3150 -37912 3065 -37848
rect 3129 -37912 3149 -37848
rect -3150 -37928 3149 -37912
rect -3150 -37992 3065 -37928
rect 3129 -37992 3149 -37928
rect -3150 -38008 3149 -37992
rect -3150 -38072 3065 -38008
rect 3129 -38072 3149 -38008
rect -3150 -38088 3149 -38072
rect -3150 -38152 3065 -38088
rect 3129 -38152 3149 -38088
rect -3150 -38168 3149 -38152
rect -3150 -38232 3065 -38168
rect 3129 -38232 3149 -38168
rect -3150 -38248 3149 -38232
rect -3150 -38312 3065 -38248
rect 3129 -38312 3149 -38248
rect -3150 -38328 3149 -38312
rect -3150 -38392 3065 -38328
rect 3129 -38392 3149 -38328
rect -3150 -38408 3149 -38392
rect -3150 -38472 3065 -38408
rect 3129 -38472 3149 -38408
rect -3150 -38488 3149 -38472
rect -3150 -38552 3065 -38488
rect 3129 -38552 3149 -38488
rect -3150 -38568 3149 -38552
rect -3150 -38632 3065 -38568
rect 3129 -38632 3149 -38568
rect -3150 -38648 3149 -38632
rect -3150 -38712 3065 -38648
rect 3129 -38712 3149 -38648
rect -3150 -38728 3149 -38712
rect -3150 -38792 3065 -38728
rect 3129 -38792 3149 -38728
rect -3150 -38808 3149 -38792
rect -3150 -38872 3065 -38808
rect 3129 -38872 3149 -38808
rect -3150 -38888 3149 -38872
rect -3150 -38952 3065 -38888
rect 3129 -38952 3149 -38888
rect -3150 -38968 3149 -38952
rect -3150 -39032 3065 -38968
rect 3129 -39032 3149 -38968
rect -3150 -39048 3149 -39032
rect -3150 -39112 3065 -39048
rect 3129 -39112 3149 -39048
rect -3150 -39128 3149 -39112
rect -3150 -39192 3065 -39128
rect 3129 -39192 3149 -39128
rect -3150 -39208 3149 -39192
rect -3150 -39272 3065 -39208
rect 3129 -39272 3149 -39208
rect -3150 -39288 3149 -39272
rect -3150 -39352 3065 -39288
rect 3129 -39352 3149 -39288
rect -3150 -39368 3149 -39352
rect -3150 -39432 3065 -39368
rect 3129 -39432 3149 -39368
rect -3150 -39448 3149 -39432
rect -3150 -39512 3065 -39448
rect 3129 -39512 3149 -39448
rect -3150 -39528 3149 -39512
rect -3150 -39592 3065 -39528
rect 3129 -39592 3149 -39528
rect -3150 -39608 3149 -39592
rect -3150 -39672 3065 -39608
rect 3129 -39672 3149 -39608
rect -3150 -39688 3149 -39672
rect -3150 -39752 3065 -39688
rect 3129 -39752 3149 -39688
rect -3150 -39768 3149 -39752
rect -3150 -39832 3065 -39768
rect 3129 -39832 3149 -39768
rect -3150 -39848 3149 -39832
rect -3150 -39912 3065 -39848
rect 3129 -39912 3149 -39848
rect -3150 -39928 3149 -39912
rect -3150 -39992 3065 -39928
rect 3129 -39992 3149 -39928
rect -3150 -40008 3149 -39992
rect -3150 -40072 3065 -40008
rect 3129 -40072 3149 -40008
rect -3150 -40088 3149 -40072
rect -3150 -40152 3065 -40088
rect 3129 -40152 3149 -40088
rect -3150 -40168 3149 -40152
rect -3150 -40232 3065 -40168
rect 3129 -40232 3149 -40168
rect -3150 -40248 3149 -40232
rect -3150 -40312 3065 -40248
rect 3129 -40312 3149 -40248
rect -3150 -40328 3149 -40312
rect -3150 -40392 3065 -40328
rect 3129 -40392 3149 -40328
rect -3150 -40408 3149 -40392
rect -3150 -40472 3065 -40408
rect 3129 -40472 3149 -40408
rect -3150 -40488 3149 -40472
rect -3150 -40552 3065 -40488
rect 3129 -40552 3149 -40488
rect -3150 -40568 3149 -40552
rect -3150 -40632 3065 -40568
rect 3129 -40632 3149 -40568
rect -3150 -40648 3149 -40632
rect -3150 -40712 3065 -40648
rect 3129 -40712 3149 -40648
rect -3150 -40728 3149 -40712
rect -3150 -40792 3065 -40728
rect 3129 -40792 3149 -40728
rect -3150 -40808 3149 -40792
rect -3150 -40872 3065 -40808
rect 3129 -40872 3149 -40808
rect -3150 -40900 3149 -40872
rect 3169 -34728 9468 -34700
rect 3169 -34792 9384 -34728
rect 9448 -34792 9468 -34728
rect 3169 -34808 9468 -34792
rect 3169 -34872 9384 -34808
rect 9448 -34872 9468 -34808
rect 3169 -34888 9468 -34872
rect 3169 -34952 9384 -34888
rect 9448 -34952 9468 -34888
rect 3169 -34968 9468 -34952
rect 3169 -35032 9384 -34968
rect 9448 -35032 9468 -34968
rect 3169 -35048 9468 -35032
rect 3169 -35112 9384 -35048
rect 9448 -35112 9468 -35048
rect 3169 -35128 9468 -35112
rect 3169 -35192 9384 -35128
rect 9448 -35192 9468 -35128
rect 3169 -35208 9468 -35192
rect 3169 -35272 9384 -35208
rect 9448 -35272 9468 -35208
rect 3169 -35288 9468 -35272
rect 3169 -35352 9384 -35288
rect 9448 -35352 9468 -35288
rect 3169 -35368 9468 -35352
rect 3169 -35432 9384 -35368
rect 9448 -35432 9468 -35368
rect 3169 -35448 9468 -35432
rect 3169 -35512 9384 -35448
rect 9448 -35512 9468 -35448
rect 3169 -35528 9468 -35512
rect 3169 -35592 9384 -35528
rect 9448 -35592 9468 -35528
rect 3169 -35608 9468 -35592
rect 3169 -35672 9384 -35608
rect 9448 -35672 9468 -35608
rect 3169 -35688 9468 -35672
rect 3169 -35752 9384 -35688
rect 9448 -35752 9468 -35688
rect 3169 -35768 9468 -35752
rect 3169 -35832 9384 -35768
rect 9448 -35832 9468 -35768
rect 3169 -35848 9468 -35832
rect 3169 -35912 9384 -35848
rect 9448 -35912 9468 -35848
rect 3169 -35928 9468 -35912
rect 3169 -35992 9384 -35928
rect 9448 -35992 9468 -35928
rect 3169 -36008 9468 -35992
rect 3169 -36072 9384 -36008
rect 9448 -36072 9468 -36008
rect 3169 -36088 9468 -36072
rect 3169 -36152 9384 -36088
rect 9448 -36152 9468 -36088
rect 3169 -36168 9468 -36152
rect 3169 -36232 9384 -36168
rect 9448 -36232 9468 -36168
rect 3169 -36248 9468 -36232
rect 3169 -36312 9384 -36248
rect 9448 -36312 9468 -36248
rect 3169 -36328 9468 -36312
rect 3169 -36392 9384 -36328
rect 9448 -36392 9468 -36328
rect 3169 -36408 9468 -36392
rect 3169 -36472 9384 -36408
rect 9448 -36472 9468 -36408
rect 3169 -36488 9468 -36472
rect 3169 -36552 9384 -36488
rect 9448 -36552 9468 -36488
rect 3169 -36568 9468 -36552
rect 3169 -36632 9384 -36568
rect 9448 -36632 9468 -36568
rect 3169 -36648 9468 -36632
rect 3169 -36712 9384 -36648
rect 9448 -36712 9468 -36648
rect 3169 -36728 9468 -36712
rect 3169 -36792 9384 -36728
rect 9448 -36792 9468 -36728
rect 3169 -36808 9468 -36792
rect 3169 -36872 9384 -36808
rect 9448 -36872 9468 -36808
rect 3169 -36888 9468 -36872
rect 3169 -36952 9384 -36888
rect 9448 -36952 9468 -36888
rect 3169 -36968 9468 -36952
rect 3169 -37032 9384 -36968
rect 9448 -37032 9468 -36968
rect 3169 -37048 9468 -37032
rect 3169 -37112 9384 -37048
rect 9448 -37112 9468 -37048
rect 3169 -37128 9468 -37112
rect 3169 -37192 9384 -37128
rect 9448 -37192 9468 -37128
rect 3169 -37208 9468 -37192
rect 3169 -37272 9384 -37208
rect 9448 -37272 9468 -37208
rect 3169 -37288 9468 -37272
rect 3169 -37352 9384 -37288
rect 9448 -37352 9468 -37288
rect 3169 -37368 9468 -37352
rect 3169 -37432 9384 -37368
rect 9448 -37432 9468 -37368
rect 3169 -37448 9468 -37432
rect 3169 -37512 9384 -37448
rect 9448 -37512 9468 -37448
rect 3169 -37528 9468 -37512
rect 3169 -37592 9384 -37528
rect 9448 -37592 9468 -37528
rect 3169 -37608 9468 -37592
rect 3169 -37672 9384 -37608
rect 9448 -37672 9468 -37608
rect 3169 -37688 9468 -37672
rect 3169 -37752 9384 -37688
rect 9448 -37752 9468 -37688
rect 3169 -37768 9468 -37752
rect 3169 -37832 9384 -37768
rect 9448 -37832 9468 -37768
rect 3169 -37848 9468 -37832
rect 3169 -37912 9384 -37848
rect 9448 -37912 9468 -37848
rect 3169 -37928 9468 -37912
rect 3169 -37992 9384 -37928
rect 9448 -37992 9468 -37928
rect 3169 -38008 9468 -37992
rect 3169 -38072 9384 -38008
rect 9448 -38072 9468 -38008
rect 3169 -38088 9468 -38072
rect 3169 -38152 9384 -38088
rect 9448 -38152 9468 -38088
rect 3169 -38168 9468 -38152
rect 3169 -38232 9384 -38168
rect 9448 -38232 9468 -38168
rect 3169 -38248 9468 -38232
rect 3169 -38312 9384 -38248
rect 9448 -38312 9468 -38248
rect 3169 -38328 9468 -38312
rect 3169 -38392 9384 -38328
rect 9448 -38392 9468 -38328
rect 3169 -38408 9468 -38392
rect 3169 -38472 9384 -38408
rect 9448 -38472 9468 -38408
rect 3169 -38488 9468 -38472
rect 3169 -38552 9384 -38488
rect 9448 -38552 9468 -38488
rect 3169 -38568 9468 -38552
rect 3169 -38632 9384 -38568
rect 9448 -38632 9468 -38568
rect 3169 -38648 9468 -38632
rect 3169 -38712 9384 -38648
rect 9448 -38712 9468 -38648
rect 3169 -38728 9468 -38712
rect 3169 -38792 9384 -38728
rect 9448 -38792 9468 -38728
rect 3169 -38808 9468 -38792
rect 3169 -38872 9384 -38808
rect 9448 -38872 9468 -38808
rect 3169 -38888 9468 -38872
rect 3169 -38952 9384 -38888
rect 9448 -38952 9468 -38888
rect 3169 -38968 9468 -38952
rect 3169 -39032 9384 -38968
rect 9448 -39032 9468 -38968
rect 3169 -39048 9468 -39032
rect 3169 -39112 9384 -39048
rect 9448 -39112 9468 -39048
rect 3169 -39128 9468 -39112
rect 3169 -39192 9384 -39128
rect 9448 -39192 9468 -39128
rect 3169 -39208 9468 -39192
rect 3169 -39272 9384 -39208
rect 9448 -39272 9468 -39208
rect 3169 -39288 9468 -39272
rect 3169 -39352 9384 -39288
rect 9448 -39352 9468 -39288
rect 3169 -39368 9468 -39352
rect 3169 -39432 9384 -39368
rect 9448 -39432 9468 -39368
rect 3169 -39448 9468 -39432
rect 3169 -39512 9384 -39448
rect 9448 -39512 9468 -39448
rect 3169 -39528 9468 -39512
rect 3169 -39592 9384 -39528
rect 9448 -39592 9468 -39528
rect 3169 -39608 9468 -39592
rect 3169 -39672 9384 -39608
rect 9448 -39672 9468 -39608
rect 3169 -39688 9468 -39672
rect 3169 -39752 9384 -39688
rect 9448 -39752 9468 -39688
rect 3169 -39768 9468 -39752
rect 3169 -39832 9384 -39768
rect 9448 -39832 9468 -39768
rect 3169 -39848 9468 -39832
rect 3169 -39912 9384 -39848
rect 9448 -39912 9468 -39848
rect 3169 -39928 9468 -39912
rect 3169 -39992 9384 -39928
rect 9448 -39992 9468 -39928
rect 3169 -40008 9468 -39992
rect 3169 -40072 9384 -40008
rect 9448 -40072 9468 -40008
rect 3169 -40088 9468 -40072
rect 3169 -40152 9384 -40088
rect 9448 -40152 9468 -40088
rect 3169 -40168 9468 -40152
rect 3169 -40232 9384 -40168
rect 9448 -40232 9468 -40168
rect 3169 -40248 9468 -40232
rect 3169 -40312 9384 -40248
rect 9448 -40312 9468 -40248
rect 3169 -40328 9468 -40312
rect 3169 -40392 9384 -40328
rect 9448 -40392 9468 -40328
rect 3169 -40408 9468 -40392
rect 3169 -40472 9384 -40408
rect 9448 -40472 9468 -40408
rect 3169 -40488 9468 -40472
rect 3169 -40552 9384 -40488
rect 9448 -40552 9468 -40488
rect 3169 -40568 9468 -40552
rect 3169 -40632 9384 -40568
rect 9448 -40632 9468 -40568
rect 3169 -40648 9468 -40632
rect 3169 -40712 9384 -40648
rect 9448 -40712 9468 -40648
rect 3169 -40728 9468 -40712
rect 3169 -40792 9384 -40728
rect 9448 -40792 9468 -40728
rect 3169 -40808 9468 -40792
rect 3169 -40872 9384 -40808
rect 9448 -40872 9468 -40808
rect 3169 -40900 9468 -40872
rect 9488 -34728 15787 -34700
rect 9488 -34792 15703 -34728
rect 15767 -34792 15787 -34728
rect 9488 -34808 15787 -34792
rect 9488 -34872 15703 -34808
rect 15767 -34872 15787 -34808
rect 9488 -34888 15787 -34872
rect 9488 -34952 15703 -34888
rect 15767 -34952 15787 -34888
rect 9488 -34968 15787 -34952
rect 9488 -35032 15703 -34968
rect 15767 -35032 15787 -34968
rect 9488 -35048 15787 -35032
rect 9488 -35112 15703 -35048
rect 15767 -35112 15787 -35048
rect 9488 -35128 15787 -35112
rect 9488 -35192 15703 -35128
rect 15767 -35192 15787 -35128
rect 9488 -35208 15787 -35192
rect 9488 -35272 15703 -35208
rect 15767 -35272 15787 -35208
rect 9488 -35288 15787 -35272
rect 9488 -35352 15703 -35288
rect 15767 -35352 15787 -35288
rect 9488 -35368 15787 -35352
rect 9488 -35432 15703 -35368
rect 15767 -35432 15787 -35368
rect 9488 -35448 15787 -35432
rect 9488 -35512 15703 -35448
rect 15767 -35512 15787 -35448
rect 9488 -35528 15787 -35512
rect 9488 -35592 15703 -35528
rect 15767 -35592 15787 -35528
rect 9488 -35608 15787 -35592
rect 9488 -35672 15703 -35608
rect 15767 -35672 15787 -35608
rect 9488 -35688 15787 -35672
rect 9488 -35752 15703 -35688
rect 15767 -35752 15787 -35688
rect 9488 -35768 15787 -35752
rect 9488 -35832 15703 -35768
rect 15767 -35832 15787 -35768
rect 9488 -35848 15787 -35832
rect 9488 -35912 15703 -35848
rect 15767 -35912 15787 -35848
rect 9488 -35928 15787 -35912
rect 9488 -35992 15703 -35928
rect 15767 -35992 15787 -35928
rect 9488 -36008 15787 -35992
rect 9488 -36072 15703 -36008
rect 15767 -36072 15787 -36008
rect 9488 -36088 15787 -36072
rect 9488 -36152 15703 -36088
rect 15767 -36152 15787 -36088
rect 9488 -36168 15787 -36152
rect 9488 -36232 15703 -36168
rect 15767 -36232 15787 -36168
rect 9488 -36248 15787 -36232
rect 9488 -36312 15703 -36248
rect 15767 -36312 15787 -36248
rect 9488 -36328 15787 -36312
rect 9488 -36392 15703 -36328
rect 15767 -36392 15787 -36328
rect 9488 -36408 15787 -36392
rect 9488 -36472 15703 -36408
rect 15767 -36472 15787 -36408
rect 9488 -36488 15787 -36472
rect 9488 -36552 15703 -36488
rect 15767 -36552 15787 -36488
rect 9488 -36568 15787 -36552
rect 9488 -36632 15703 -36568
rect 15767 -36632 15787 -36568
rect 9488 -36648 15787 -36632
rect 9488 -36712 15703 -36648
rect 15767 -36712 15787 -36648
rect 9488 -36728 15787 -36712
rect 9488 -36792 15703 -36728
rect 15767 -36792 15787 -36728
rect 9488 -36808 15787 -36792
rect 9488 -36872 15703 -36808
rect 15767 -36872 15787 -36808
rect 9488 -36888 15787 -36872
rect 9488 -36952 15703 -36888
rect 15767 -36952 15787 -36888
rect 9488 -36968 15787 -36952
rect 9488 -37032 15703 -36968
rect 15767 -37032 15787 -36968
rect 9488 -37048 15787 -37032
rect 9488 -37112 15703 -37048
rect 15767 -37112 15787 -37048
rect 9488 -37128 15787 -37112
rect 9488 -37192 15703 -37128
rect 15767 -37192 15787 -37128
rect 9488 -37208 15787 -37192
rect 9488 -37272 15703 -37208
rect 15767 -37272 15787 -37208
rect 9488 -37288 15787 -37272
rect 9488 -37352 15703 -37288
rect 15767 -37352 15787 -37288
rect 9488 -37368 15787 -37352
rect 9488 -37432 15703 -37368
rect 15767 -37432 15787 -37368
rect 9488 -37448 15787 -37432
rect 9488 -37512 15703 -37448
rect 15767 -37512 15787 -37448
rect 9488 -37528 15787 -37512
rect 9488 -37592 15703 -37528
rect 15767 -37592 15787 -37528
rect 9488 -37608 15787 -37592
rect 9488 -37672 15703 -37608
rect 15767 -37672 15787 -37608
rect 9488 -37688 15787 -37672
rect 9488 -37752 15703 -37688
rect 15767 -37752 15787 -37688
rect 9488 -37768 15787 -37752
rect 9488 -37832 15703 -37768
rect 15767 -37832 15787 -37768
rect 9488 -37848 15787 -37832
rect 9488 -37912 15703 -37848
rect 15767 -37912 15787 -37848
rect 9488 -37928 15787 -37912
rect 9488 -37992 15703 -37928
rect 15767 -37992 15787 -37928
rect 9488 -38008 15787 -37992
rect 9488 -38072 15703 -38008
rect 15767 -38072 15787 -38008
rect 9488 -38088 15787 -38072
rect 9488 -38152 15703 -38088
rect 15767 -38152 15787 -38088
rect 9488 -38168 15787 -38152
rect 9488 -38232 15703 -38168
rect 15767 -38232 15787 -38168
rect 9488 -38248 15787 -38232
rect 9488 -38312 15703 -38248
rect 15767 -38312 15787 -38248
rect 9488 -38328 15787 -38312
rect 9488 -38392 15703 -38328
rect 15767 -38392 15787 -38328
rect 9488 -38408 15787 -38392
rect 9488 -38472 15703 -38408
rect 15767 -38472 15787 -38408
rect 9488 -38488 15787 -38472
rect 9488 -38552 15703 -38488
rect 15767 -38552 15787 -38488
rect 9488 -38568 15787 -38552
rect 9488 -38632 15703 -38568
rect 15767 -38632 15787 -38568
rect 9488 -38648 15787 -38632
rect 9488 -38712 15703 -38648
rect 15767 -38712 15787 -38648
rect 9488 -38728 15787 -38712
rect 9488 -38792 15703 -38728
rect 15767 -38792 15787 -38728
rect 9488 -38808 15787 -38792
rect 9488 -38872 15703 -38808
rect 15767 -38872 15787 -38808
rect 9488 -38888 15787 -38872
rect 9488 -38952 15703 -38888
rect 15767 -38952 15787 -38888
rect 9488 -38968 15787 -38952
rect 9488 -39032 15703 -38968
rect 15767 -39032 15787 -38968
rect 9488 -39048 15787 -39032
rect 9488 -39112 15703 -39048
rect 15767 -39112 15787 -39048
rect 9488 -39128 15787 -39112
rect 9488 -39192 15703 -39128
rect 15767 -39192 15787 -39128
rect 9488 -39208 15787 -39192
rect 9488 -39272 15703 -39208
rect 15767 -39272 15787 -39208
rect 9488 -39288 15787 -39272
rect 9488 -39352 15703 -39288
rect 15767 -39352 15787 -39288
rect 9488 -39368 15787 -39352
rect 9488 -39432 15703 -39368
rect 15767 -39432 15787 -39368
rect 9488 -39448 15787 -39432
rect 9488 -39512 15703 -39448
rect 15767 -39512 15787 -39448
rect 9488 -39528 15787 -39512
rect 9488 -39592 15703 -39528
rect 15767 -39592 15787 -39528
rect 9488 -39608 15787 -39592
rect 9488 -39672 15703 -39608
rect 15767 -39672 15787 -39608
rect 9488 -39688 15787 -39672
rect 9488 -39752 15703 -39688
rect 15767 -39752 15787 -39688
rect 9488 -39768 15787 -39752
rect 9488 -39832 15703 -39768
rect 15767 -39832 15787 -39768
rect 9488 -39848 15787 -39832
rect 9488 -39912 15703 -39848
rect 15767 -39912 15787 -39848
rect 9488 -39928 15787 -39912
rect 9488 -39992 15703 -39928
rect 15767 -39992 15787 -39928
rect 9488 -40008 15787 -39992
rect 9488 -40072 15703 -40008
rect 15767 -40072 15787 -40008
rect 9488 -40088 15787 -40072
rect 9488 -40152 15703 -40088
rect 15767 -40152 15787 -40088
rect 9488 -40168 15787 -40152
rect 9488 -40232 15703 -40168
rect 15767 -40232 15787 -40168
rect 9488 -40248 15787 -40232
rect 9488 -40312 15703 -40248
rect 15767 -40312 15787 -40248
rect 9488 -40328 15787 -40312
rect 9488 -40392 15703 -40328
rect 15767 -40392 15787 -40328
rect 9488 -40408 15787 -40392
rect 9488 -40472 15703 -40408
rect 15767 -40472 15787 -40408
rect 9488 -40488 15787 -40472
rect 9488 -40552 15703 -40488
rect 15767 -40552 15787 -40488
rect 9488 -40568 15787 -40552
rect 9488 -40632 15703 -40568
rect 15767 -40632 15787 -40568
rect 9488 -40648 15787 -40632
rect 9488 -40712 15703 -40648
rect 15767 -40712 15787 -40648
rect 9488 -40728 15787 -40712
rect 9488 -40792 15703 -40728
rect 15767 -40792 15787 -40728
rect 9488 -40808 15787 -40792
rect 9488 -40872 15703 -40808
rect 15767 -40872 15787 -40808
rect 9488 -40900 15787 -40872
rect 15807 -34728 22106 -34700
rect 15807 -34792 22022 -34728
rect 22086 -34792 22106 -34728
rect 15807 -34808 22106 -34792
rect 15807 -34872 22022 -34808
rect 22086 -34872 22106 -34808
rect 15807 -34888 22106 -34872
rect 15807 -34952 22022 -34888
rect 22086 -34952 22106 -34888
rect 15807 -34968 22106 -34952
rect 15807 -35032 22022 -34968
rect 22086 -35032 22106 -34968
rect 15807 -35048 22106 -35032
rect 15807 -35112 22022 -35048
rect 22086 -35112 22106 -35048
rect 15807 -35128 22106 -35112
rect 15807 -35192 22022 -35128
rect 22086 -35192 22106 -35128
rect 15807 -35208 22106 -35192
rect 15807 -35272 22022 -35208
rect 22086 -35272 22106 -35208
rect 15807 -35288 22106 -35272
rect 15807 -35352 22022 -35288
rect 22086 -35352 22106 -35288
rect 15807 -35368 22106 -35352
rect 15807 -35432 22022 -35368
rect 22086 -35432 22106 -35368
rect 15807 -35448 22106 -35432
rect 15807 -35512 22022 -35448
rect 22086 -35512 22106 -35448
rect 15807 -35528 22106 -35512
rect 15807 -35592 22022 -35528
rect 22086 -35592 22106 -35528
rect 15807 -35608 22106 -35592
rect 15807 -35672 22022 -35608
rect 22086 -35672 22106 -35608
rect 15807 -35688 22106 -35672
rect 15807 -35752 22022 -35688
rect 22086 -35752 22106 -35688
rect 15807 -35768 22106 -35752
rect 15807 -35832 22022 -35768
rect 22086 -35832 22106 -35768
rect 15807 -35848 22106 -35832
rect 15807 -35912 22022 -35848
rect 22086 -35912 22106 -35848
rect 15807 -35928 22106 -35912
rect 15807 -35992 22022 -35928
rect 22086 -35992 22106 -35928
rect 15807 -36008 22106 -35992
rect 15807 -36072 22022 -36008
rect 22086 -36072 22106 -36008
rect 15807 -36088 22106 -36072
rect 15807 -36152 22022 -36088
rect 22086 -36152 22106 -36088
rect 15807 -36168 22106 -36152
rect 15807 -36232 22022 -36168
rect 22086 -36232 22106 -36168
rect 15807 -36248 22106 -36232
rect 15807 -36312 22022 -36248
rect 22086 -36312 22106 -36248
rect 15807 -36328 22106 -36312
rect 15807 -36392 22022 -36328
rect 22086 -36392 22106 -36328
rect 15807 -36408 22106 -36392
rect 15807 -36472 22022 -36408
rect 22086 -36472 22106 -36408
rect 15807 -36488 22106 -36472
rect 15807 -36552 22022 -36488
rect 22086 -36552 22106 -36488
rect 15807 -36568 22106 -36552
rect 15807 -36632 22022 -36568
rect 22086 -36632 22106 -36568
rect 15807 -36648 22106 -36632
rect 15807 -36712 22022 -36648
rect 22086 -36712 22106 -36648
rect 15807 -36728 22106 -36712
rect 15807 -36792 22022 -36728
rect 22086 -36792 22106 -36728
rect 15807 -36808 22106 -36792
rect 15807 -36872 22022 -36808
rect 22086 -36872 22106 -36808
rect 15807 -36888 22106 -36872
rect 15807 -36952 22022 -36888
rect 22086 -36952 22106 -36888
rect 15807 -36968 22106 -36952
rect 15807 -37032 22022 -36968
rect 22086 -37032 22106 -36968
rect 15807 -37048 22106 -37032
rect 15807 -37112 22022 -37048
rect 22086 -37112 22106 -37048
rect 15807 -37128 22106 -37112
rect 15807 -37192 22022 -37128
rect 22086 -37192 22106 -37128
rect 15807 -37208 22106 -37192
rect 15807 -37272 22022 -37208
rect 22086 -37272 22106 -37208
rect 15807 -37288 22106 -37272
rect 15807 -37352 22022 -37288
rect 22086 -37352 22106 -37288
rect 15807 -37368 22106 -37352
rect 15807 -37432 22022 -37368
rect 22086 -37432 22106 -37368
rect 15807 -37448 22106 -37432
rect 15807 -37512 22022 -37448
rect 22086 -37512 22106 -37448
rect 15807 -37528 22106 -37512
rect 15807 -37592 22022 -37528
rect 22086 -37592 22106 -37528
rect 15807 -37608 22106 -37592
rect 15807 -37672 22022 -37608
rect 22086 -37672 22106 -37608
rect 15807 -37688 22106 -37672
rect 15807 -37752 22022 -37688
rect 22086 -37752 22106 -37688
rect 15807 -37768 22106 -37752
rect 15807 -37832 22022 -37768
rect 22086 -37832 22106 -37768
rect 15807 -37848 22106 -37832
rect 15807 -37912 22022 -37848
rect 22086 -37912 22106 -37848
rect 15807 -37928 22106 -37912
rect 15807 -37992 22022 -37928
rect 22086 -37992 22106 -37928
rect 15807 -38008 22106 -37992
rect 15807 -38072 22022 -38008
rect 22086 -38072 22106 -38008
rect 15807 -38088 22106 -38072
rect 15807 -38152 22022 -38088
rect 22086 -38152 22106 -38088
rect 15807 -38168 22106 -38152
rect 15807 -38232 22022 -38168
rect 22086 -38232 22106 -38168
rect 15807 -38248 22106 -38232
rect 15807 -38312 22022 -38248
rect 22086 -38312 22106 -38248
rect 15807 -38328 22106 -38312
rect 15807 -38392 22022 -38328
rect 22086 -38392 22106 -38328
rect 15807 -38408 22106 -38392
rect 15807 -38472 22022 -38408
rect 22086 -38472 22106 -38408
rect 15807 -38488 22106 -38472
rect 15807 -38552 22022 -38488
rect 22086 -38552 22106 -38488
rect 15807 -38568 22106 -38552
rect 15807 -38632 22022 -38568
rect 22086 -38632 22106 -38568
rect 15807 -38648 22106 -38632
rect 15807 -38712 22022 -38648
rect 22086 -38712 22106 -38648
rect 15807 -38728 22106 -38712
rect 15807 -38792 22022 -38728
rect 22086 -38792 22106 -38728
rect 15807 -38808 22106 -38792
rect 15807 -38872 22022 -38808
rect 22086 -38872 22106 -38808
rect 15807 -38888 22106 -38872
rect 15807 -38952 22022 -38888
rect 22086 -38952 22106 -38888
rect 15807 -38968 22106 -38952
rect 15807 -39032 22022 -38968
rect 22086 -39032 22106 -38968
rect 15807 -39048 22106 -39032
rect 15807 -39112 22022 -39048
rect 22086 -39112 22106 -39048
rect 15807 -39128 22106 -39112
rect 15807 -39192 22022 -39128
rect 22086 -39192 22106 -39128
rect 15807 -39208 22106 -39192
rect 15807 -39272 22022 -39208
rect 22086 -39272 22106 -39208
rect 15807 -39288 22106 -39272
rect 15807 -39352 22022 -39288
rect 22086 -39352 22106 -39288
rect 15807 -39368 22106 -39352
rect 15807 -39432 22022 -39368
rect 22086 -39432 22106 -39368
rect 15807 -39448 22106 -39432
rect 15807 -39512 22022 -39448
rect 22086 -39512 22106 -39448
rect 15807 -39528 22106 -39512
rect 15807 -39592 22022 -39528
rect 22086 -39592 22106 -39528
rect 15807 -39608 22106 -39592
rect 15807 -39672 22022 -39608
rect 22086 -39672 22106 -39608
rect 15807 -39688 22106 -39672
rect 15807 -39752 22022 -39688
rect 22086 -39752 22106 -39688
rect 15807 -39768 22106 -39752
rect 15807 -39832 22022 -39768
rect 22086 -39832 22106 -39768
rect 15807 -39848 22106 -39832
rect 15807 -39912 22022 -39848
rect 22086 -39912 22106 -39848
rect 15807 -39928 22106 -39912
rect 15807 -39992 22022 -39928
rect 22086 -39992 22106 -39928
rect 15807 -40008 22106 -39992
rect 15807 -40072 22022 -40008
rect 22086 -40072 22106 -40008
rect 15807 -40088 22106 -40072
rect 15807 -40152 22022 -40088
rect 22086 -40152 22106 -40088
rect 15807 -40168 22106 -40152
rect 15807 -40232 22022 -40168
rect 22086 -40232 22106 -40168
rect 15807 -40248 22106 -40232
rect 15807 -40312 22022 -40248
rect 22086 -40312 22106 -40248
rect 15807 -40328 22106 -40312
rect 15807 -40392 22022 -40328
rect 22086 -40392 22106 -40328
rect 15807 -40408 22106 -40392
rect 15807 -40472 22022 -40408
rect 22086 -40472 22106 -40408
rect 15807 -40488 22106 -40472
rect 15807 -40552 22022 -40488
rect 22086 -40552 22106 -40488
rect 15807 -40568 22106 -40552
rect 15807 -40632 22022 -40568
rect 22086 -40632 22106 -40568
rect 15807 -40648 22106 -40632
rect 15807 -40712 22022 -40648
rect 22086 -40712 22106 -40648
rect 15807 -40728 22106 -40712
rect 15807 -40792 22022 -40728
rect 22086 -40792 22106 -40728
rect 15807 -40808 22106 -40792
rect 15807 -40872 22022 -40808
rect 22086 -40872 22106 -40808
rect 15807 -40900 22106 -40872
rect 22126 -34728 28425 -34700
rect 22126 -34792 28341 -34728
rect 28405 -34792 28425 -34728
rect 22126 -34808 28425 -34792
rect 22126 -34872 28341 -34808
rect 28405 -34872 28425 -34808
rect 22126 -34888 28425 -34872
rect 22126 -34952 28341 -34888
rect 28405 -34952 28425 -34888
rect 22126 -34968 28425 -34952
rect 22126 -35032 28341 -34968
rect 28405 -35032 28425 -34968
rect 22126 -35048 28425 -35032
rect 22126 -35112 28341 -35048
rect 28405 -35112 28425 -35048
rect 22126 -35128 28425 -35112
rect 22126 -35192 28341 -35128
rect 28405 -35192 28425 -35128
rect 22126 -35208 28425 -35192
rect 22126 -35272 28341 -35208
rect 28405 -35272 28425 -35208
rect 22126 -35288 28425 -35272
rect 22126 -35352 28341 -35288
rect 28405 -35352 28425 -35288
rect 22126 -35368 28425 -35352
rect 22126 -35432 28341 -35368
rect 28405 -35432 28425 -35368
rect 22126 -35448 28425 -35432
rect 22126 -35512 28341 -35448
rect 28405 -35512 28425 -35448
rect 22126 -35528 28425 -35512
rect 22126 -35592 28341 -35528
rect 28405 -35592 28425 -35528
rect 22126 -35608 28425 -35592
rect 22126 -35672 28341 -35608
rect 28405 -35672 28425 -35608
rect 22126 -35688 28425 -35672
rect 22126 -35752 28341 -35688
rect 28405 -35752 28425 -35688
rect 22126 -35768 28425 -35752
rect 22126 -35832 28341 -35768
rect 28405 -35832 28425 -35768
rect 22126 -35848 28425 -35832
rect 22126 -35912 28341 -35848
rect 28405 -35912 28425 -35848
rect 22126 -35928 28425 -35912
rect 22126 -35992 28341 -35928
rect 28405 -35992 28425 -35928
rect 22126 -36008 28425 -35992
rect 22126 -36072 28341 -36008
rect 28405 -36072 28425 -36008
rect 22126 -36088 28425 -36072
rect 22126 -36152 28341 -36088
rect 28405 -36152 28425 -36088
rect 22126 -36168 28425 -36152
rect 22126 -36232 28341 -36168
rect 28405 -36232 28425 -36168
rect 22126 -36248 28425 -36232
rect 22126 -36312 28341 -36248
rect 28405 -36312 28425 -36248
rect 22126 -36328 28425 -36312
rect 22126 -36392 28341 -36328
rect 28405 -36392 28425 -36328
rect 22126 -36408 28425 -36392
rect 22126 -36472 28341 -36408
rect 28405 -36472 28425 -36408
rect 22126 -36488 28425 -36472
rect 22126 -36552 28341 -36488
rect 28405 -36552 28425 -36488
rect 22126 -36568 28425 -36552
rect 22126 -36632 28341 -36568
rect 28405 -36632 28425 -36568
rect 22126 -36648 28425 -36632
rect 22126 -36712 28341 -36648
rect 28405 -36712 28425 -36648
rect 22126 -36728 28425 -36712
rect 22126 -36792 28341 -36728
rect 28405 -36792 28425 -36728
rect 22126 -36808 28425 -36792
rect 22126 -36872 28341 -36808
rect 28405 -36872 28425 -36808
rect 22126 -36888 28425 -36872
rect 22126 -36952 28341 -36888
rect 28405 -36952 28425 -36888
rect 22126 -36968 28425 -36952
rect 22126 -37032 28341 -36968
rect 28405 -37032 28425 -36968
rect 22126 -37048 28425 -37032
rect 22126 -37112 28341 -37048
rect 28405 -37112 28425 -37048
rect 22126 -37128 28425 -37112
rect 22126 -37192 28341 -37128
rect 28405 -37192 28425 -37128
rect 22126 -37208 28425 -37192
rect 22126 -37272 28341 -37208
rect 28405 -37272 28425 -37208
rect 22126 -37288 28425 -37272
rect 22126 -37352 28341 -37288
rect 28405 -37352 28425 -37288
rect 22126 -37368 28425 -37352
rect 22126 -37432 28341 -37368
rect 28405 -37432 28425 -37368
rect 22126 -37448 28425 -37432
rect 22126 -37512 28341 -37448
rect 28405 -37512 28425 -37448
rect 22126 -37528 28425 -37512
rect 22126 -37592 28341 -37528
rect 28405 -37592 28425 -37528
rect 22126 -37608 28425 -37592
rect 22126 -37672 28341 -37608
rect 28405 -37672 28425 -37608
rect 22126 -37688 28425 -37672
rect 22126 -37752 28341 -37688
rect 28405 -37752 28425 -37688
rect 22126 -37768 28425 -37752
rect 22126 -37832 28341 -37768
rect 28405 -37832 28425 -37768
rect 22126 -37848 28425 -37832
rect 22126 -37912 28341 -37848
rect 28405 -37912 28425 -37848
rect 22126 -37928 28425 -37912
rect 22126 -37992 28341 -37928
rect 28405 -37992 28425 -37928
rect 22126 -38008 28425 -37992
rect 22126 -38072 28341 -38008
rect 28405 -38072 28425 -38008
rect 22126 -38088 28425 -38072
rect 22126 -38152 28341 -38088
rect 28405 -38152 28425 -38088
rect 22126 -38168 28425 -38152
rect 22126 -38232 28341 -38168
rect 28405 -38232 28425 -38168
rect 22126 -38248 28425 -38232
rect 22126 -38312 28341 -38248
rect 28405 -38312 28425 -38248
rect 22126 -38328 28425 -38312
rect 22126 -38392 28341 -38328
rect 28405 -38392 28425 -38328
rect 22126 -38408 28425 -38392
rect 22126 -38472 28341 -38408
rect 28405 -38472 28425 -38408
rect 22126 -38488 28425 -38472
rect 22126 -38552 28341 -38488
rect 28405 -38552 28425 -38488
rect 22126 -38568 28425 -38552
rect 22126 -38632 28341 -38568
rect 28405 -38632 28425 -38568
rect 22126 -38648 28425 -38632
rect 22126 -38712 28341 -38648
rect 28405 -38712 28425 -38648
rect 22126 -38728 28425 -38712
rect 22126 -38792 28341 -38728
rect 28405 -38792 28425 -38728
rect 22126 -38808 28425 -38792
rect 22126 -38872 28341 -38808
rect 28405 -38872 28425 -38808
rect 22126 -38888 28425 -38872
rect 22126 -38952 28341 -38888
rect 28405 -38952 28425 -38888
rect 22126 -38968 28425 -38952
rect 22126 -39032 28341 -38968
rect 28405 -39032 28425 -38968
rect 22126 -39048 28425 -39032
rect 22126 -39112 28341 -39048
rect 28405 -39112 28425 -39048
rect 22126 -39128 28425 -39112
rect 22126 -39192 28341 -39128
rect 28405 -39192 28425 -39128
rect 22126 -39208 28425 -39192
rect 22126 -39272 28341 -39208
rect 28405 -39272 28425 -39208
rect 22126 -39288 28425 -39272
rect 22126 -39352 28341 -39288
rect 28405 -39352 28425 -39288
rect 22126 -39368 28425 -39352
rect 22126 -39432 28341 -39368
rect 28405 -39432 28425 -39368
rect 22126 -39448 28425 -39432
rect 22126 -39512 28341 -39448
rect 28405 -39512 28425 -39448
rect 22126 -39528 28425 -39512
rect 22126 -39592 28341 -39528
rect 28405 -39592 28425 -39528
rect 22126 -39608 28425 -39592
rect 22126 -39672 28341 -39608
rect 28405 -39672 28425 -39608
rect 22126 -39688 28425 -39672
rect 22126 -39752 28341 -39688
rect 28405 -39752 28425 -39688
rect 22126 -39768 28425 -39752
rect 22126 -39832 28341 -39768
rect 28405 -39832 28425 -39768
rect 22126 -39848 28425 -39832
rect 22126 -39912 28341 -39848
rect 28405 -39912 28425 -39848
rect 22126 -39928 28425 -39912
rect 22126 -39992 28341 -39928
rect 28405 -39992 28425 -39928
rect 22126 -40008 28425 -39992
rect 22126 -40072 28341 -40008
rect 28405 -40072 28425 -40008
rect 22126 -40088 28425 -40072
rect 22126 -40152 28341 -40088
rect 28405 -40152 28425 -40088
rect 22126 -40168 28425 -40152
rect 22126 -40232 28341 -40168
rect 28405 -40232 28425 -40168
rect 22126 -40248 28425 -40232
rect 22126 -40312 28341 -40248
rect 28405 -40312 28425 -40248
rect 22126 -40328 28425 -40312
rect 22126 -40392 28341 -40328
rect 28405 -40392 28425 -40328
rect 22126 -40408 28425 -40392
rect 22126 -40472 28341 -40408
rect 28405 -40472 28425 -40408
rect 22126 -40488 28425 -40472
rect 22126 -40552 28341 -40488
rect 28405 -40552 28425 -40488
rect 22126 -40568 28425 -40552
rect 22126 -40632 28341 -40568
rect 28405 -40632 28425 -40568
rect 22126 -40648 28425 -40632
rect 22126 -40712 28341 -40648
rect 28405 -40712 28425 -40648
rect 22126 -40728 28425 -40712
rect 22126 -40792 28341 -40728
rect 28405 -40792 28425 -40728
rect 22126 -40808 28425 -40792
rect 22126 -40872 28341 -40808
rect 28405 -40872 28425 -40808
rect 22126 -40900 28425 -40872
rect 28445 -34728 34744 -34700
rect 28445 -34792 34660 -34728
rect 34724 -34792 34744 -34728
rect 28445 -34808 34744 -34792
rect 28445 -34872 34660 -34808
rect 34724 -34872 34744 -34808
rect 28445 -34888 34744 -34872
rect 28445 -34952 34660 -34888
rect 34724 -34952 34744 -34888
rect 28445 -34968 34744 -34952
rect 28445 -35032 34660 -34968
rect 34724 -35032 34744 -34968
rect 28445 -35048 34744 -35032
rect 28445 -35112 34660 -35048
rect 34724 -35112 34744 -35048
rect 28445 -35128 34744 -35112
rect 28445 -35192 34660 -35128
rect 34724 -35192 34744 -35128
rect 28445 -35208 34744 -35192
rect 28445 -35272 34660 -35208
rect 34724 -35272 34744 -35208
rect 28445 -35288 34744 -35272
rect 28445 -35352 34660 -35288
rect 34724 -35352 34744 -35288
rect 28445 -35368 34744 -35352
rect 28445 -35432 34660 -35368
rect 34724 -35432 34744 -35368
rect 28445 -35448 34744 -35432
rect 28445 -35512 34660 -35448
rect 34724 -35512 34744 -35448
rect 28445 -35528 34744 -35512
rect 28445 -35592 34660 -35528
rect 34724 -35592 34744 -35528
rect 28445 -35608 34744 -35592
rect 28445 -35672 34660 -35608
rect 34724 -35672 34744 -35608
rect 28445 -35688 34744 -35672
rect 28445 -35752 34660 -35688
rect 34724 -35752 34744 -35688
rect 28445 -35768 34744 -35752
rect 28445 -35832 34660 -35768
rect 34724 -35832 34744 -35768
rect 28445 -35848 34744 -35832
rect 28445 -35912 34660 -35848
rect 34724 -35912 34744 -35848
rect 28445 -35928 34744 -35912
rect 28445 -35992 34660 -35928
rect 34724 -35992 34744 -35928
rect 28445 -36008 34744 -35992
rect 28445 -36072 34660 -36008
rect 34724 -36072 34744 -36008
rect 28445 -36088 34744 -36072
rect 28445 -36152 34660 -36088
rect 34724 -36152 34744 -36088
rect 28445 -36168 34744 -36152
rect 28445 -36232 34660 -36168
rect 34724 -36232 34744 -36168
rect 28445 -36248 34744 -36232
rect 28445 -36312 34660 -36248
rect 34724 -36312 34744 -36248
rect 28445 -36328 34744 -36312
rect 28445 -36392 34660 -36328
rect 34724 -36392 34744 -36328
rect 28445 -36408 34744 -36392
rect 28445 -36472 34660 -36408
rect 34724 -36472 34744 -36408
rect 28445 -36488 34744 -36472
rect 28445 -36552 34660 -36488
rect 34724 -36552 34744 -36488
rect 28445 -36568 34744 -36552
rect 28445 -36632 34660 -36568
rect 34724 -36632 34744 -36568
rect 28445 -36648 34744 -36632
rect 28445 -36712 34660 -36648
rect 34724 -36712 34744 -36648
rect 28445 -36728 34744 -36712
rect 28445 -36792 34660 -36728
rect 34724 -36792 34744 -36728
rect 28445 -36808 34744 -36792
rect 28445 -36872 34660 -36808
rect 34724 -36872 34744 -36808
rect 28445 -36888 34744 -36872
rect 28445 -36952 34660 -36888
rect 34724 -36952 34744 -36888
rect 28445 -36968 34744 -36952
rect 28445 -37032 34660 -36968
rect 34724 -37032 34744 -36968
rect 28445 -37048 34744 -37032
rect 28445 -37112 34660 -37048
rect 34724 -37112 34744 -37048
rect 28445 -37128 34744 -37112
rect 28445 -37192 34660 -37128
rect 34724 -37192 34744 -37128
rect 28445 -37208 34744 -37192
rect 28445 -37272 34660 -37208
rect 34724 -37272 34744 -37208
rect 28445 -37288 34744 -37272
rect 28445 -37352 34660 -37288
rect 34724 -37352 34744 -37288
rect 28445 -37368 34744 -37352
rect 28445 -37432 34660 -37368
rect 34724 -37432 34744 -37368
rect 28445 -37448 34744 -37432
rect 28445 -37512 34660 -37448
rect 34724 -37512 34744 -37448
rect 28445 -37528 34744 -37512
rect 28445 -37592 34660 -37528
rect 34724 -37592 34744 -37528
rect 28445 -37608 34744 -37592
rect 28445 -37672 34660 -37608
rect 34724 -37672 34744 -37608
rect 28445 -37688 34744 -37672
rect 28445 -37752 34660 -37688
rect 34724 -37752 34744 -37688
rect 28445 -37768 34744 -37752
rect 28445 -37832 34660 -37768
rect 34724 -37832 34744 -37768
rect 28445 -37848 34744 -37832
rect 28445 -37912 34660 -37848
rect 34724 -37912 34744 -37848
rect 28445 -37928 34744 -37912
rect 28445 -37992 34660 -37928
rect 34724 -37992 34744 -37928
rect 28445 -38008 34744 -37992
rect 28445 -38072 34660 -38008
rect 34724 -38072 34744 -38008
rect 28445 -38088 34744 -38072
rect 28445 -38152 34660 -38088
rect 34724 -38152 34744 -38088
rect 28445 -38168 34744 -38152
rect 28445 -38232 34660 -38168
rect 34724 -38232 34744 -38168
rect 28445 -38248 34744 -38232
rect 28445 -38312 34660 -38248
rect 34724 -38312 34744 -38248
rect 28445 -38328 34744 -38312
rect 28445 -38392 34660 -38328
rect 34724 -38392 34744 -38328
rect 28445 -38408 34744 -38392
rect 28445 -38472 34660 -38408
rect 34724 -38472 34744 -38408
rect 28445 -38488 34744 -38472
rect 28445 -38552 34660 -38488
rect 34724 -38552 34744 -38488
rect 28445 -38568 34744 -38552
rect 28445 -38632 34660 -38568
rect 34724 -38632 34744 -38568
rect 28445 -38648 34744 -38632
rect 28445 -38712 34660 -38648
rect 34724 -38712 34744 -38648
rect 28445 -38728 34744 -38712
rect 28445 -38792 34660 -38728
rect 34724 -38792 34744 -38728
rect 28445 -38808 34744 -38792
rect 28445 -38872 34660 -38808
rect 34724 -38872 34744 -38808
rect 28445 -38888 34744 -38872
rect 28445 -38952 34660 -38888
rect 34724 -38952 34744 -38888
rect 28445 -38968 34744 -38952
rect 28445 -39032 34660 -38968
rect 34724 -39032 34744 -38968
rect 28445 -39048 34744 -39032
rect 28445 -39112 34660 -39048
rect 34724 -39112 34744 -39048
rect 28445 -39128 34744 -39112
rect 28445 -39192 34660 -39128
rect 34724 -39192 34744 -39128
rect 28445 -39208 34744 -39192
rect 28445 -39272 34660 -39208
rect 34724 -39272 34744 -39208
rect 28445 -39288 34744 -39272
rect 28445 -39352 34660 -39288
rect 34724 -39352 34744 -39288
rect 28445 -39368 34744 -39352
rect 28445 -39432 34660 -39368
rect 34724 -39432 34744 -39368
rect 28445 -39448 34744 -39432
rect 28445 -39512 34660 -39448
rect 34724 -39512 34744 -39448
rect 28445 -39528 34744 -39512
rect 28445 -39592 34660 -39528
rect 34724 -39592 34744 -39528
rect 28445 -39608 34744 -39592
rect 28445 -39672 34660 -39608
rect 34724 -39672 34744 -39608
rect 28445 -39688 34744 -39672
rect 28445 -39752 34660 -39688
rect 34724 -39752 34744 -39688
rect 28445 -39768 34744 -39752
rect 28445 -39832 34660 -39768
rect 34724 -39832 34744 -39768
rect 28445 -39848 34744 -39832
rect 28445 -39912 34660 -39848
rect 34724 -39912 34744 -39848
rect 28445 -39928 34744 -39912
rect 28445 -39992 34660 -39928
rect 34724 -39992 34744 -39928
rect 28445 -40008 34744 -39992
rect 28445 -40072 34660 -40008
rect 34724 -40072 34744 -40008
rect 28445 -40088 34744 -40072
rect 28445 -40152 34660 -40088
rect 34724 -40152 34744 -40088
rect 28445 -40168 34744 -40152
rect 28445 -40232 34660 -40168
rect 34724 -40232 34744 -40168
rect 28445 -40248 34744 -40232
rect 28445 -40312 34660 -40248
rect 34724 -40312 34744 -40248
rect 28445 -40328 34744 -40312
rect 28445 -40392 34660 -40328
rect 34724 -40392 34744 -40328
rect 28445 -40408 34744 -40392
rect 28445 -40472 34660 -40408
rect 34724 -40472 34744 -40408
rect 28445 -40488 34744 -40472
rect 28445 -40552 34660 -40488
rect 34724 -40552 34744 -40488
rect 28445 -40568 34744 -40552
rect 28445 -40632 34660 -40568
rect 34724 -40632 34744 -40568
rect 28445 -40648 34744 -40632
rect 28445 -40712 34660 -40648
rect 34724 -40712 34744 -40648
rect 28445 -40728 34744 -40712
rect 28445 -40792 34660 -40728
rect 34724 -40792 34744 -40728
rect 28445 -40808 34744 -40792
rect 28445 -40872 34660 -40808
rect 34724 -40872 34744 -40808
rect 28445 -40900 34744 -40872
rect 34764 -34728 41063 -34700
rect 34764 -34792 40979 -34728
rect 41043 -34792 41063 -34728
rect 34764 -34808 41063 -34792
rect 34764 -34872 40979 -34808
rect 41043 -34872 41063 -34808
rect 34764 -34888 41063 -34872
rect 34764 -34952 40979 -34888
rect 41043 -34952 41063 -34888
rect 34764 -34968 41063 -34952
rect 34764 -35032 40979 -34968
rect 41043 -35032 41063 -34968
rect 34764 -35048 41063 -35032
rect 34764 -35112 40979 -35048
rect 41043 -35112 41063 -35048
rect 34764 -35128 41063 -35112
rect 34764 -35192 40979 -35128
rect 41043 -35192 41063 -35128
rect 34764 -35208 41063 -35192
rect 34764 -35272 40979 -35208
rect 41043 -35272 41063 -35208
rect 34764 -35288 41063 -35272
rect 34764 -35352 40979 -35288
rect 41043 -35352 41063 -35288
rect 34764 -35368 41063 -35352
rect 34764 -35432 40979 -35368
rect 41043 -35432 41063 -35368
rect 34764 -35448 41063 -35432
rect 34764 -35512 40979 -35448
rect 41043 -35512 41063 -35448
rect 34764 -35528 41063 -35512
rect 34764 -35592 40979 -35528
rect 41043 -35592 41063 -35528
rect 34764 -35608 41063 -35592
rect 34764 -35672 40979 -35608
rect 41043 -35672 41063 -35608
rect 34764 -35688 41063 -35672
rect 34764 -35752 40979 -35688
rect 41043 -35752 41063 -35688
rect 34764 -35768 41063 -35752
rect 34764 -35832 40979 -35768
rect 41043 -35832 41063 -35768
rect 34764 -35848 41063 -35832
rect 34764 -35912 40979 -35848
rect 41043 -35912 41063 -35848
rect 34764 -35928 41063 -35912
rect 34764 -35992 40979 -35928
rect 41043 -35992 41063 -35928
rect 34764 -36008 41063 -35992
rect 34764 -36072 40979 -36008
rect 41043 -36072 41063 -36008
rect 34764 -36088 41063 -36072
rect 34764 -36152 40979 -36088
rect 41043 -36152 41063 -36088
rect 34764 -36168 41063 -36152
rect 34764 -36232 40979 -36168
rect 41043 -36232 41063 -36168
rect 34764 -36248 41063 -36232
rect 34764 -36312 40979 -36248
rect 41043 -36312 41063 -36248
rect 34764 -36328 41063 -36312
rect 34764 -36392 40979 -36328
rect 41043 -36392 41063 -36328
rect 34764 -36408 41063 -36392
rect 34764 -36472 40979 -36408
rect 41043 -36472 41063 -36408
rect 34764 -36488 41063 -36472
rect 34764 -36552 40979 -36488
rect 41043 -36552 41063 -36488
rect 34764 -36568 41063 -36552
rect 34764 -36632 40979 -36568
rect 41043 -36632 41063 -36568
rect 34764 -36648 41063 -36632
rect 34764 -36712 40979 -36648
rect 41043 -36712 41063 -36648
rect 34764 -36728 41063 -36712
rect 34764 -36792 40979 -36728
rect 41043 -36792 41063 -36728
rect 34764 -36808 41063 -36792
rect 34764 -36872 40979 -36808
rect 41043 -36872 41063 -36808
rect 34764 -36888 41063 -36872
rect 34764 -36952 40979 -36888
rect 41043 -36952 41063 -36888
rect 34764 -36968 41063 -36952
rect 34764 -37032 40979 -36968
rect 41043 -37032 41063 -36968
rect 34764 -37048 41063 -37032
rect 34764 -37112 40979 -37048
rect 41043 -37112 41063 -37048
rect 34764 -37128 41063 -37112
rect 34764 -37192 40979 -37128
rect 41043 -37192 41063 -37128
rect 34764 -37208 41063 -37192
rect 34764 -37272 40979 -37208
rect 41043 -37272 41063 -37208
rect 34764 -37288 41063 -37272
rect 34764 -37352 40979 -37288
rect 41043 -37352 41063 -37288
rect 34764 -37368 41063 -37352
rect 34764 -37432 40979 -37368
rect 41043 -37432 41063 -37368
rect 34764 -37448 41063 -37432
rect 34764 -37512 40979 -37448
rect 41043 -37512 41063 -37448
rect 34764 -37528 41063 -37512
rect 34764 -37592 40979 -37528
rect 41043 -37592 41063 -37528
rect 34764 -37608 41063 -37592
rect 34764 -37672 40979 -37608
rect 41043 -37672 41063 -37608
rect 34764 -37688 41063 -37672
rect 34764 -37752 40979 -37688
rect 41043 -37752 41063 -37688
rect 34764 -37768 41063 -37752
rect 34764 -37832 40979 -37768
rect 41043 -37832 41063 -37768
rect 34764 -37848 41063 -37832
rect 34764 -37912 40979 -37848
rect 41043 -37912 41063 -37848
rect 34764 -37928 41063 -37912
rect 34764 -37992 40979 -37928
rect 41043 -37992 41063 -37928
rect 34764 -38008 41063 -37992
rect 34764 -38072 40979 -38008
rect 41043 -38072 41063 -38008
rect 34764 -38088 41063 -38072
rect 34764 -38152 40979 -38088
rect 41043 -38152 41063 -38088
rect 34764 -38168 41063 -38152
rect 34764 -38232 40979 -38168
rect 41043 -38232 41063 -38168
rect 34764 -38248 41063 -38232
rect 34764 -38312 40979 -38248
rect 41043 -38312 41063 -38248
rect 34764 -38328 41063 -38312
rect 34764 -38392 40979 -38328
rect 41043 -38392 41063 -38328
rect 34764 -38408 41063 -38392
rect 34764 -38472 40979 -38408
rect 41043 -38472 41063 -38408
rect 34764 -38488 41063 -38472
rect 34764 -38552 40979 -38488
rect 41043 -38552 41063 -38488
rect 34764 -38568 41063 -38552
rect 34764 -38632 40979 -38568
rect 41043 -38632 41063 -38568
rect 34764 -38648 41063 -38632
rect 34764 -38712 40979 -38648
rect 41043 -38712 41063 -38648
rect 34764 -38728 41063 -38712
rect 34764 -38792 40979 -38728
rect 41043 -38792 41063 -38728
rect 34764 -38808 41063 -38792
rect 34764 -38872 40979 -38808
rect 41043 -38872 41063 -38808
rect 34764 -38888 41063 -38872
rect 34764 -38952 40979 -38888
rect 41043 -38952 41063 -38888
rect 34764 -38968 41063 -38952
rect 34764 -39032 40979 -38968
rect 41043 -39032 41063 -38968
rect 34764 -39048 41063 -39032
rect 34764 -39112 40979 -39048
rect 41043 -39112 41063 -39048
rect 34764 -39128 41063 -39112
rect 34764 -39192 40979 -39128
rect 41043 -39192 41063 -39128
rect 34764 -39208 41063 -39192
rect 34764 -39272 40979 -39208
rect 41043 -39272 41063 -39208
rect 34764 -39288 41063 -39272
rect 34764 -39352 40979 -39288
rect 41043 -39352 41063 -39288
rect 34764 -39368 41063 -39352
rect 34764 -39432 40979 -39368
rect 41043 -39432 41063 -39368
rect 34764 -39448 41063 -39432
rect 34764 -39512 40979 -39448
rect 41043 -39512 41063 -39448
rect 34764 -39528 41063 -39512
rect 34764 -39592 40979 -39528
rect 41043 -39592 41063 -39528
rect 34764 -39608 41063 -39592
rect 34764 -39672 40979 -39608
rect 41043 -39672 41063 -39608
rect 34764 -39688 41063 -39672
rect 34764 -39752 40979 -39688
rect 41043 -39752 41063 -39688
rect 34764 -39768 41063 -39752
rect 34764 -39832 40979 -39768
rect 41043 -39832 41063 -39768
rect 34764 -39848 41063 -39832
rect 34764 -39912 40979 -39848
rect 41043 -39912 41063 -39848
rect 34764 -39928 41063 -39912
rect 34764 -39992 40979 -39928
rect 41043 -39992 41063 -39928
rect 34764 -40008 41063 -39992
rect 34764 -40072 40979 -40008
rect 41043 -40072 41063 -40008
rect 34764 -40088 41063 -40072
rect 34764 -40152 40979 -40088
rect 41043 -40152 41063 -40088
rect 34764 -40168 41063 -40152
rect 34764 -40232 40979 -40168
rect 41043 -40232 41063 -40168
rect 34764 -40248 41063 -40232
rect 34764 -40312 40979 -40248
rect 41043 -40312 41063 -40248
rect 34764 -40328 41063 -40312
rect 34764 -40392 40979 -40328
rect 41043 -40392 41063 -40328
rect 34764 -40408 41063 -40392
rect 34764 -40472 40979 -40408
rect 41043 -40472 41063 -40408
rect 34764 -40488 41063 -40472
rect 34764 -40552 40979 -40488
rect 41043 -40552 41063 -40488
rect 34764 -40568 41063 -40552
rect 34764 -40632 40979 -40568
rect 41043 -40632 41063 -40568
rect 34764 -40648 41063 -40632
rect 34764 -40712 40979 -40648
rect 41043 -40712 41063 -40648
rect 34764 -40728 41063 -40712
rect 34764 -40792 40979 -40728
rect 41043 -40792 41063 -40728
rect 34764 -40808 41063 -40792
rect 34764 -40872 40979 -40808
rect 41043 -40872 41063 -40808
rect 34764 -40900 41063 -40872
rect 41083 -34728 47382 -34700
rect 41083 -34792 47298 -34728
rect 47362 -34792 47382 -34728
rect 41083 -34808 47382 -34792
rect 41083 -34872 47298 -34808
rect 47362 -34872 47382 -34808
rect 41083 -34888 47382 -34872
rect 41083 -34952 47298 -34888
rect 47362 -34952 47382 -34888
rect 41083 -34968 47382 -34952
rect 41083 -35032 47298 -34968
rect 47362 -35032 47382 -34968
rect 41083 -35048 47382 -35032
rect 41083 -35112 47298 -35048
rect 47362 -35112 47382 -35048
rect 41083 -35128 47382 -35112
rect 41083 -35192 47298 -35128
rect 47362 -35192 47382 -35128
rect 41083 -35208 47382 -35192
rect 41083 -35272 47298 -35208
rect 47362 -35272 47382 -35208
rect 41083 -35288 47382 -35272
rect 41083 -35352 47298 -35288
rect 47362 -35352 47382 -35288
rect 41083 -35368 47382 -35352
rect 41083 -35432 47298 -35368
rect 47362 -35432 47382 -35368
rect 41083 -35448 47382 -35432
rect 41083 -35512 47298 -35448
rect 47362 -35512 47382 -35448
rect 41083 -35528 47382 -35512
rect 41083 -35592 47298 -35528
rect 47362 -35592 47382 -35528
rect 41083 -35608 47382 -35592
rect 41083 -35672 47298 -35608
rect 47362 -35672 47382 -35608
rect 41083 -35688 47382 -35672
rect 41083 -35752 47298 -35688
rect 47362 -35752 47382 -35688
rect 41083 -35768 47382 -35752
rect 41083 -35832 47298 -35768
rect 47362 -35832 47382 -35768
rect 41083 -35848 47382 -35832
rect 41083 -35912 47298 -35848
rect 47362 -35912 47382 -35848
rect 41083 -35928 47382 -35912
rect 41083 -35992 47298 -35928
rect 47362 -35992 47382 -35928
rect 41083 -36008 47382 -35992
rect 41083 -36072 47298 -36008
rect 47362 -36072 47382 -36008
rect 41083 -36088 47382 -36072
rect 41083 -36152 47298 -36088
rect 47362 -36152 47382 -36088
rect 41083 -36168 47382 -36152
rect 41083 -36232 47298 -36168
rect 47362 -36232 47382 -36168
rect 41083 -36248 47382 -36232
rect 41083 -36312 47298 -36248
rect 47362 -36312 47382 -36248
rect 41083 -36328 47382 -36312
rect 41083 -36392 47298 -36328
rect 47362 -36392 47382 -36328
rect 41083 -36408 47382 -36392
rect 41083 -36472 47298 -36408
rect 47362 -36472 47382 -36408
rect 41083 -36488 47382 -36472
rect 41083 -36552 47298 -36488
rect 47362 -36552 47382 -36488
rect 41083 -36568 47382 -36552
rect 41083 -36632 47298 -36568
rect 47362 -36632 47382 -36568
rect 41083 -36648 47382 -36632
rect 41083 -36712 47298 -36648
rect 47362 -36712 47382 -36648
rect 41083 -36728 47382 -36712
rect 41083 -36792 47298 -36728
rect 47362 -36792 47382 -36728
rect 41083 -36808 47382 -36792
rect 41083 -36872 47298 -36808
rect 47362 -36872 47382 -36808
rect 41083 -36888 47382 -36872
rect 41083 -36952 47298 -36888
rect 47362 -36952 47382 -36888
rect 41083 -36968 47382 -36952
rect 41083 -37032 47298 -36968
rect 47362 -37032 47382 -36968
rect 41083 -37048 47382 -37032
rect 41083 -37112 47298 -37048
rect 47362 -37112 47382 -37048
rect 41083 -37128 47382 -37112
rect 41083 -37192 47298 -37128
rect 47362 -37192 47382 -37128
rect 41083 -37208 47382 -37192
rect 41083 -37272 47298 -37208
rect 47362 -37272 47382 -37208
rect 41083 -37288 47382 -37272
rect 41083 -37352 47298 -37288
rect 47362 -37352 47382 -37288
rect 41083 -37368 47382 -37352
rect 41083 -37432 47298 -37368
rect 47362 -37432 47382 -37368
rect 41083 -37448 47382 -37432
rect 41083 -37512 47298 -37448
rect 47362 -37512 47382 -37448
rect 41083 -37528 47382 -37512
rect 41083 -37592 47298 -37528
rect 47362 -37592 47382 -37528
rect 41083 -37608 47382 -37592
rect 41083 -37672 47298 -37608
rect 47362 -37672 47382 -37608
rect 41083 -37688 47382 -37672
rect 41083 -37752 47298 -37688
rect 47362 -37752 47382 -37688
rect 41083 -37768 47382 -37752
rect 41083 -37832 47298 -37768
rect 47362 -37832 47382 -37768
rect 41083 -37848 47382 -37832
rect 41083 -37912 47298 -37848
rect 47362 -37912 47382 -37848
rect 41083 -37928 47382 -37912
rect 41083 -37992 47298 -37928
rect 47362 -37992 47382 -37928
rect 41083 -38008 47382 -37992
rect 41083 -38072 47298 -38008
rect 47362 -38072 47382 -38008
rect 41083 -38088 47382 -38072
rect 41083 -38152 47298 -38088
rect 47362 -38152 47382 -38088
rect 41083 -38168 47382 -38152
rect 41083 -38232 47298 -38168
rect 47362 -38232 47382 -38168
rect 41083 -38248 47382 -38232
rect 41083 -38312 47298 -38248
rect 47362 -38312 47382 -38248
rect 41083 -38328 47382 -38312
rect 41083 -38392 47298 -38328
rect 47362 -38392 47382 -38328
rect 41083 -38408 47382 -38392
rect 41083 -38472 47298 -38408
rect 47362 -38472 47382 -38408
rect 41083 -38488 47382 -38472
rect 41083 -38552 47298 -38488
rect 47362 -38552 47382 -38488
rect 41083 -38568 47382 -38552
rect 41083 -38632 47298 -38568
rect 47362 -38632 47382 -38568
rect 41083 -38648 47382 -38632
rect 41083 -38712 47298 -38648
rect 47362 -38712 47382 -38648
rect 41083 -38728 47382 -38712
rect 41083 -38792 47298 -38728
rect 47362 -38792 47382 -38728
rect 41083 -38808 47382 -38792
rect 41083 -38872 47298 -38808
rect 47362 -38872 47382 -38808
rect 41083 -38888 47382 -38872
rect 41083 -38952 47298 -38888
rect 47362 -38952 47382 -38888
rect 41083 -38968 47382 -38952
rect 41083 -39032 47298 -38968
rect 47362 -39032 47382 -38968
rect 41083 -39048 47382 -39032
rect 41083 -39112 47298 -39048
rect 47362 -39112 47382 -39048
rect 41083 -39128 47382 -39112
rect 41083 -39192 47298 -39128
rect 47362 -39192 47382 -39128
rect 41083 -39208 47382 -39192
rect 41083 -39272 47298 -39208
rect 47362 -39272 47382 -39208
rect 41083 -39288 47382 -39272
rect 41083 -39352 47298 -39288
rect 47362 -39352 47382 -39288
rect 41083 -39368 47382 -39352
rect 41083 -39432 47298 -39368
rect 47362 -39432 47382 -39368
rect 41083 -39448 47382 -39432
rect 41083 -39512 47298 -39448
rect 47362 -39512 47382 -39448
rect 41083 -39528 47382 -39512
rect 41083 -39592 47298 -39528
rect 47362 -39592 47382 -39528
rect 41083 -39608 47382 -39592
rect 41083 -39672 47298 -39608
rect 47362 -39672 47382 -39608
rect 41083 -39688 47382 -39672
rect 41083 -39752 47298 -39688
rect 47362 -39752 47382 -39688
rect 41083 -39768 47382 -39752
rect 41083 -39832 47298 -39768
rect 47362 -39832 47382 -39768
rect 41083 -39848 47382 -39832
rect 41083 -39912 47298 -39848
rect 47362 -39912 47382 -39848
rect 41083 -39928 47382 -39912
rect 41083 -39992 47298 -39928
rect 47362 -39992 47382 -39928
rect 41083 -40008 47382 -39992
rect 41083 -40072 47298 -40008
rect 47362 -40072 47382 -40008
rect 41083 -40088 47382 -40072
rect 41083 -40152 47298 -40088
rect 47362 -40152 47382 -40088
rect 41083 -40168 47382 -40152
rect 41083 -40232 47298 -40168
rect 47362 -40232 47382 -40168
rect 41083 -40248 47382 -40232
rect 41083 -40312 47298 -40248
rect 47362 -40312 47382 -40248
rect 41083 -40328 47382 -40312
rect 41083 -40392 47298 -40328
rect 47362 -40392 47382 -40328
rect 41083 -40408 47382 -40392
rect 41083 -40472 47298 -40408
rect 47362 -40472 47382 -40408
rect 41083 -40488 47382 -40472
rect 41083 -40552 47298 -40488
rect 47362 -40552 47382 -40488
rect 41083 -40568 47382 -40552
rect 41083 -40632 47298 -40568
rect 47362 -40632 47382 -40568
rect 41083 -40648 47382 -40632
rect 41083 -40712 47298 -40648
rect 47362 -40712 47382 -40648
rect 41083 -40728 47382 -40712
rect 41083 -40792 47298 -40728
rect 47362 -40792 47382 -40728
rect 41083 -40808 47382 -40792
rect 41083 -40872 47298 -40808
rect 47362 -40872 47382 -40808
rect 41083 -40900 47382 -40872
rect -47383 -41028 -41084 -41000
rect -47383 -41092 -41168 -41028
rect -41104 -41092 -41084 -41028
rect -47383 -41108 -41084 -41092
rect -47383 -41172 -41168 -41108
rect -41104 -41172 -41084 -41108
rect -47383 -41188 -41084 -41172
rect -47383 -41252 -41168 -41188
rect -41104 -41252 -41084 -41188
rect -47383 -41268 -41084 -41252
rect -47383 -41332 -41168 -41268
rect -41104 -41332 -41084 -41268
rect -47383 -41348 -41084 -41332
rect -47383 -41412 -41168 -41348
rect -41104 -41412 -41084 -41348
rect -47383 -41428 -41084 -41412
rect -47383 -41492 -41168 -41428
rect -41104 -41492 -41084 -41428
rect -47383 -41508 -41084 -41492
rect -47383 -41572 -41168 -41508
rect -41104 -41572 -41084 -41508
rect -47383 -41588 -41084 -41572
rect -47383 -41652 -41168 -41588
rect -41104 -41652 -41084 -41588
rect -47383 -41668 -41084 -41652
rect -47383 -41732 -41168 -41668
rect -41104 -41732 -41084 -41668
rect -47383 -41748 -41084 -41732
rect -47383 -41812 -41168 -41748
rect -41104 -41812 -41084 -41748
rect -47383 -41828 -41084 -41812
rect -47383 -41892 -41168 -41828
rect -41104 -41892 -41084 -41828
rect -47383 -41908 -41084 -41892
rect -47383 -41972 -41168 -41908
rect -41104 -41972 -41084 -41908
rect -47383 -41988 -41084 -41972
rect -47383 -42052 -41168 -41988
rect -41104 -42052 -41084 -41988
rect -47383 -42068 -41084 -42052
rect -47383 -42132 -41168 -42068
rect -41104 -42132 -41084 -42068
rect -47383 -42148 -41084 -42132
rect -47383 -42212 -41168 -42148
rect -41104 -42212 -41084 -42148
rect -47383 -42228 -41084 -42212
rect -47383 -42292 -41168 -42228
rect -41104 -42292 -41084 -42228
rect -47383 -42308 -41084 -42292
rect -47383 -42372 -41168 -42308
rect -41104 -42372 -41084 -42308
rect -47383 -42388 -41084 -42372
rect -47383 -42452 -41168 -42388
rect -41104 -42452 -41084 -42388
rect -47383 -42468 -41084 -42452
rect -47383 -42532 -41168 -42468
rect -41104 -42532 -41084 -42468
rect -47383 -42548 -41084 -42532
rect -47383 -42612 -41168 -42548
rect -41104 -42612 -41084 -42548
rect -47383 -42628 -41084 -42612
rect -47383 -42692 -41168 -42628
rect -41104 -42692 -41084 -42628
rect -47383 -42708 -41084 -42692
rect -47383 -42772 -41168 -42708
rect -41104 -42772 -41084 -42708
rect -47383 -42788 -41084 -42772
rect -47383 -42852 -41168 -42788
rect -41104 -42852 -41084 -42788
rect -47383 -42868 -41084 -42852
rect -47383 -42932 -41168 -42868
rect -41104 -42932 -41084 -42868
rect -47383 -42948 -41084 -42932
rect -47383 -43012 -41168 -42948
rect -41104 -43012 -41084 -42948
rect -47383 -43028 -41084 -43012
rect -47383 -43092 -41168 -43028
rect -41104 -43092 -41084 -43028
rect -47383 -43108 -41084 -43092
rect -47383 -43172 -41168 -43108
rect -41104 -43172 -41084 -43108
rect -47383 -43188 -41084 -43172
rect -47383 -43252 -41168 -43188
rect -41104 -43252 -41084 -43188
rect -47383 -43268 -41084 -43252
rect -47383 -43332 -41168 -43268
rect -41104 -43332 -41084 -43268
rect -47383 -43348 -41084 -43332
rect -47383 -43412 -41168 -43348
rect -41104 -43412 -41084 -43348
rect -47383 -43428 -41084 -43412
rect -47383 -43492 -41168 -43428
rect -41104 -43492 -41084 -43428
rect -47383 -43508 -41084 -43492
rect -47383 -43572 -41168 -43508
rect -41104 -43572 -41084 -43508
rect -47383 -43588 -41084 -43572
rect -47383 -43652 -41168 -43588
rect -41104 -43652 -41084 -43588
rect -47383 -43668 -41084 -43652
rect -47383 -43732 -41168 -43668
rect -41104 -43732 -41084 -43668
rect -47383 -43748 -41084 -43732
rect -47383 -43812 -41168 -43748
rect -41104 -43812 -41084 -43748
rect -47383 -43828 -41084 -43812
rect -47383 -43892 -41168 -43828
rect -41104 -43892 -41084 -43828
rect -47383 -43908 -41084 -43892
rect -47383 -43972 -41168 -43908
rect -41104 -43972 -41084 -43908
rect -47383 -43988 -41084 -43972
rect -47383 -44052 -41168 -43988
rect -41104 -44052 -41084 -43988
rect -47383 -44068 -41084 -44052
rect -47383 -44132 -41168 -44068
rect -41104 -44132 -41084 -44068
rect -47383 -44148 -41084 -44132
rect -47383 -44212 -41168 -44148
rect -41104 -44212 -41084 -44148
rect -47383 -44228 -41084 -44212
rect -47383 -44292 -41168 -44228
rect -41104 -44292 -41084 -44228
rect -47383 -44308 -41084 -44292
rect -47383 -44372 -41168 -44308
rect -41104 -44372 -41084 -44308
rect -47383 -44388 -41084 -44372
rect -47383 -44452 -41168 -44388
rect -41104 -44452 -41084 -44388
rect -47383 -44468 -41084 -44452
rect -47383 -44532 -41168 -44468
rect -41104 -44532 -41084 -44468
rect -47383 -44548 -41084 -44532
rect -47383 -44612 -41168 -44548
rect -41104 -44612 -41084 -44548
rect -47383 -44628 -41084 -44612
rect -47383 -44692 -41168 -44628
rect -41104 -44692 -41084 -44628
rect -47383 -44708 -41084 -44692
rect -47383 -44772 -41168 -44708
rect -41104 -44772 -41084 -44708
rect -47383 -44788 -41084 -44772
rect -47383 -44852 -41168 -44788
rect -41104 -44852 -41084 -44788
rect -47383 -44868 -41084 -44852
rect -47383 -44932 -41168 -44868
rect -41104 -44932 -41084 -44868
rect -47383 -44948 -41084 -44932
rect -47383 -45012 -41168 -44948
rect -41104 -45012 -41084 -44948
rect -47383 -45028 -41084 -45012
rect -47383 -45092 -41168 -45028
rect -41104 -45092 -41084 -45028
rect -47383 -45108 -41084 -45092
rect -47383 -45172 -41168 -45108
rect -41104 -45172 -41084 -45108
rect -47383 -45188 -41084 -45172
rect -47383 -45252 -41168 -45188
rect -41104 -45252 -41084 -45188
rect -47383 -45268 -41084 -45252
rect -47383 -45332 -41168 -45268
rect -41104 -45332 -41084 -45268
rect -47383 -45348 -41084 -45332
rect -47383 -45412 -41168 -45348
rect -41104 -45412 -41084 -45348
rect -47383 -45428 -41084 -45412
rect -47383 -45492 -41168 -45428
rect -41104 -45492 -41084 -45428
rect -47383 -45508 -41084 -45492
rect -47383 -45572 -41168 -45508
rect -41104 -45572 -41084 -45508
rect -47383 -45588 -41084 -45572
rect -47383 -45652 -41168 -45588
rect -41104 -45652 -41084 -45588
rect -47383 -45668 -41084 -45652
rect -47383 -45732 -41168 -45668
rect -41104 -45732 -41084 -45668
rect -47383 -45748 -41084 -45732
rect -47383 -45812 -41168 -45748
rect -41104 -45812 -41084 -45748
rect -47383 -45828 -41084 -45812
rect -47383 -45892 -41168 -45828
rect -41104 -45892 -41084 -45828
rect -47383 -45908 -41084 -45892
rect -47383 -45972 -41168 -45908
rect -41104 -45972 -41084 -45908
rect -47383 -45988 -41084 -45972
rect -47383 -46052 -41168 -45988
rect -41104 -46052 -41084 -45988
rect -47383 -46068 -41084 -46052
rect -47383 -46132 -41168 -46068
rect -41104 -46132 -41084 -46068
rect -47383 -46148 -41084 -46132
rect -47383 -46212 -41168 -46148
rect -41104 -46212 -41084 -46148
rect -47383 -46228 -41084 -46212
rect -47383 -46292 -41168 -46228
rect -41104 -46292 -41084 -46228
rect -47383 -46308 -41084 -46292
rect -47383 -46372 -41168 -46308
rect -41104 -46372 -41084 -46308
rect -47383 -46388 -41084 -46372
rect -47383 -46452 -41168 -46388
rect -41104 -46452 -41084 -46388
rect -47383 -46468 -41084 -46452
rect -47383 -46532 -41168 -46468
rect -41104 -46532 -41084 -46468
rect -47383 -46548 -41084 -46532
rect -47383 -46612 -41168 -46548
rect -41104 -46612 -41084 -46548
rect -47383 -46628 -41084 -46612
rect -47383 -46692 -41168 -46628
rect -41104 -46692 -41084 -46628
rect -47383 -46708 -41084 -46692
rect -47383 -46772 -41168 -46708
rect -41104 -46772 -41084 -46708
rect -47383 -46788 -41084 -46772
rect -47383 -46852 -41168 -46788
rect -41104 -46852 -41084 -46788
rect -47383 -46868 -41084 -46852
rect -47383 -46932 -41168 -46868
rect -41104 -46932 -41084 -46868
rect -47383 -46948 -41084 -46932
rect -47383 -47012 -41168 -46948
rect -41104 -47012 -41084 -46948
rect -47383 -47028 -41084 -47012
rect -47383 -47092 -41168 -47028
rect -41104 -47092 -41084 -47028
rect -47383 -47108 -41084 -47092
rect -47383 -47172 -41168 -47108
rect -41104 -47172 -41084 -47108
rect -47383 -47200 -41084 -47172
rect -41064 -41028 -34765 -41000
rect -41064 -41092 -34849 -41028
rect -34785 -41092 -34765 -41028
rect -41064 -41108 -34765 -41092
rect -41064 -41172 -34849 -41108
rect -34785 -41172 -34765 -41108
rect -41064 -41188 -34765 -41172
rect -41064 -41252 -34849 -41188
rect -34785 -41252 -34765 -41188
rect -41064 -41268 -34765 -41252
rect -41064 -41332 -34849 -41268
rect -34785 -41332 -34765 -41268
rect -41064 -41348 -34765 -41332
rect -41064 -41412 -34849 -41348
rect -34785 -41412 -34765 -41348
rect -41064 -41428 -34765 -41412
rect -41064 -41492 -34849 -41428
rect -34785 -41492 -34765 -41428
rect -41064 -41508 -34765 -41492
rect -41064 -41572 -34849 -41508
rect -34785 -41572 -34765 -41508
rect -41064 -41588 -34765 -41572
rect -41064 -41652 -34849 -41588
rect -34785 -41652 -34765 -41588
rect -41064 -41668 -34765 -41652
rect -41064 -41732 -34849 -41668
rect -34785 -41732 -34765 -41668
rect -41064 -41748 -34765 -41732
rect -41064 -41812 -34849 -41748
rect -34785 -41812 -34765 -41748
rect -41064 -41828 -34765 -41812
rect -41064 -41892 -34849 -41828
rect -34785 -41892 -34765 -41828
rect -41064 -41908 -34765 -41892
rect -41064 -41972 -34849 -41908
rect -34785 -41972 -34765 -41908
rect -41064 -41988 -34765 -41972
rect -41064 -42052 -34849 -41988
rect -34785 -42052 -34765 -41988
rect -41064 -42068 -34765 -42052
rect -41064 -42132 -34849 -42068
rect -34785 -42132 -34765 -42068
rect -41064 -42148 -34765 -42132
rect -41064 -42212 -34849 -42148
rect -34785 -42212 -34765 -42148
rect -41064 -42228 -34765 -42212
rect -41064 -42292 -34849 -42228
rect -34785 -42292 -34765 -42228
rect -41064 -42308 -34765 -42292
rect -41064 -42372 -34849 -42308
rect -34785 -42372 -34765 -42308
rect -41064 -42388 -34765 -42372
rect -41064 -42452 -34849 -42388
rect -34785 -42452 -34765 -42388
rect -41064 -42468 -34765 -42452
rect -41064 -42532 -34849 -42468
rect -34785 -42532 -34765 -42468
rect -41064 -42548 -34765 -42532
rect -41064 -42612 -34849 -42548
rect -34785 -42612 -34765 -42548
rect -41064 -42628 -34765 -42612
rect -41064 -42692 -34849 -42628
rect -34785 -42692 -34765 -42628
rect -41064 -42708 -34765 -42692
rect -41064 -42772 -34849 -42708
rect -34785 -42772 -34765 -42708
rect -41064 -42788 -34765 -42772
rect -41064 -42852 -34849 -42788
rect -34785 -42852 -34765 -42788
rect -41064 -42868 -34765 -42852
rect -41064 -42932 -34849 -42868
rect -34785 -42932 -34765 -42868
rect -41064 -42948 -34765 -42932
rect -41064 -43012 -34849 -42948
rect -34785 -43012 -34765 -42948
rect -41064 -43028 -34765 -43012
rect -41064 -43092 -34849 -43028
rect -34785 -43092 -34765 -43028
rect -41064 -43108 -34765 -43092
rect -41064 -43172 -34849 -43108
rect -34785 -43172 -34765 -43108
rect -41064 -43188 -34765 -43172
rect -41064 -43252 -34849 -43188
rect -34785 -43252 -34765 -43188
rect -41064 -43268 -34765 -43252
rect -41064 -43332 -34849 -43268
rect -34785 -43332 -34765 -43268
rect -41064 -43348 -34765 -43332
rect -41064 -43412 -34849 -43348
rect -34785 -43412 -34765 -43348
rect -41064 -43428 -34765 -43412
rect -41064 -43492 -34849 -43428
rect -34785 -43492 -34765 -43428
rect -41064 -43508 -34765 -43492
rect -41064 -43572 -34849 -43508
rect -34785 -43572 -34765 -43508
rect -41064 -43588 -34765 -43572
rect -41064 -43652 -34849 -43588
rect -34785 -43652 -34765 -43588
rect -41064 -43668 -34765 -43652
rect -41064 -43732 -34849 -43668
rect -34785 -43732 -34765 -43668
rect -41064 -43748 -34765 -43732
rect -41064 -43812 -34849 -43748
rect -34785 -43812 -34765 -43748
rect -41064 -43828 -34765 -43812
rect -41064 -43892 -34849 -43828
rect -34785 -43892 -34765 -43828
rect -41064 -43908 -34765 -43892
rect -41064 -43972 -34849 -43908
rect -34785 -43972 -34765 -43908
rect -41064 -43988 -34765 -43972
rect -41064 -44052 -34849 -43988
rect -34785 -44052 -34765 -43988
rect -41064 -44068 -34765 -44052
rect -41064 -44132 -34849 -44068
rect -34785 -44132 -34765 -44068
rect -41064 -44148 -34765 -44132
rect -41064 -44212 -34849 -44148
rect -34785 -44212 -34765 -44148
rect -41064 -44228 -34765 -44212
rect -41064 -44292 -34849 -44228
rect -34785 -44292 -34765 -44228
rect -41064 -44308 -34765 -44292
rect -41064 -44372 -34849 -44308
rect -34785 -44372 -34765 -44308
rect -41064 -44388 -34765 -44372
rect -41064 -44452 -34849 -44388
rect -34785 -44452 -34765 -44388
rect -41064 -44468 -34765 -44452
rect -41064 -44532 -34849 -44468
rect -34785 -44532 -34765 -44468
rect -41064 -44548 -34765 -44532
rect -41064 -44612 -34849 -44548
rect -34785 -44612 -34765 -44548
rect -41064 -44628 -34765 -44612
rect -41064 -44692 -34849 -44628
rect -34785 -44692 -34765 -44628
rect -41064 -44708 -34765 -44692
rect -41064 -44772 -34849 -44708
rect -34785 -44772 -34765 -44708
rect -41064 -44788 -34765 -44772
rect -41064 -44852 -34849 -44788
rect -34785 -44852 -34765 -44788
rect -41064 -44868 -34765 -44852
rect -41064 -44932 -34849 -44868
rect -34785 -44932 -34765 -44868
rect -41064 -44948 -34765 -44932
rect -41064 -45012 -34849 -44948
rect -34785 -45012 -34765 -44948
rect -41064 -45028 -34765 -45012
rect -41064 -45092 -34849 -45028
rect -34785 -45092 -34765 -45028
rect -41064 -45108 -34765 -45092
rect -41064 -45172 -34849 -45108
rect -34785 -45172 -34765 -45108
rect -41064 -45188 -34765 -45172
rect -41064 -45252 -34849 -45188
rect -34785 -45252 -34765 -45188
rect -41064 -45268 -34765 -45252
rect -41064 -45332 -34849 -45268
rect -34785 -45332 -34765 -45268
rect -41064 -45348 -34765 -45332
rect -41064 -45412 -34849 -45348
rect -34785 -45412 -34765 -45348
rect -41064 -45428 -34765 -45412
rect -41064 -45492 -34849 -45428
rect -34785 -45492 -34765 -45428
rect -41064 -45508 -34765 -45492
rect -41064 -45572 -34849 -45508
rect -34785 -45572 -34765 -45508
rect -41064 -45588 -34765 -45572
rect -41064 -45652 -34849 -45588
rect -34785 -45652 -34765 -45588
rect -41064 -45668 -34765 -45652
rect -41064 -45732 -34849 -45668
rect -34785 -45732 -34765 -45668
rect -41064 -45748 -34765 -45732
rect -41064 -45812 -34849 -45748
rect -34785 -45812 -34765 -45748
rect -41064 -45828 -34765 -45812
rect -41064 -45892 -34849 -45828
rect -34785 -45892 -34765 -45828
rect -41064 -45908 -34765 -45892
rect -41064 -45972 -34849 -45908
rect -34785 -45972 -34765 -45908
rect -41064 -45988 -34765 -45972
rect -41064 -46052 -34849 -45988
rect -34785 -46052 -34765 -45988
rect -41064 -46068 -34765 -46052
rect -41064 -46132 -34849 -46068
rect -34785 -46132 -34765 -46068
rect -41064 -46148 -34765 -46132
rect -41064 -46212 -34849 -46148
rect -34785 -46212 -34765 -46148
rect -41064 -46228 -34765 -46212
rect -41064 -46292 -34849 -46228
rect -34785 -46292 -34765 -46228
rect -41064 -46308 -34765 -46292
rect -41064 -46372 -34849 -46308
rect -34785 -46372 -34765 -46308
rect -41064 -46388 -34765 -46372
rect -41064 -46452 -34849 -46388
rect -34785 -46452 -34765 -46388
rect -41064 -46468 -34765 -46452
rect -41064 -46532 -34849 -46468
rect -34785 -46532 -34765 -46468
rect -41064 -46548 -34765 -46532
rect -41064 -46612 -34849 -46548
rect -34785 -46612 -34765 -46548
rect -41064 -46628 -34765 -46612
rect -41064 -46692 -34849 -46628
rect -34785 -46692 -34765 -46628
rect -41064 -46708 -34765 -46692
rect -41064 -46772 -34849 -46708
rect -34785 -46772 -34765 -46708
rect -41064 -46788 -34765 -46772
rect -41064 -46852 -34849 -46788
rect -34785 -46852 -34765 -46788
rect -41064 -46868 -34765 -46852
rect -41064 -46932 -34849 -46868
rect -34785 -46932 -34765 -46868
rect -41064 -46948 -34765 -46932
rect -41064 -47012 -34849 -46948
rect -34785 -47012 -34765 -46948
rect -41064 -47028 -34765 -47012
rect -41064 -47092 -34849 -47028
rect -34785 -47092 -34765 -47028
rect -41064 -47108 -34765 -47092
rect -41064 -47172 -34849 -47108
rect -34785 -47172 -34765 -47108
rect -41064 -47200 -34765 -47172
rect -34745 -41028 -28446 -41000
rect -34745 -41092 -28530 -41028
rect -28466 -41092 -28446 -41028
rect -34745 -41108 -28446 -41092
rect -34745 -41172 -28530 -41108
rect -28466 -41172 -28446 -41108
rect -34745 -41188 -28446 -41172
rect -34745 -41252 -28530 -41188
rect -28466 -41252 -28446 -41188
rect -34745 -41268 -28446 -41252
rect -34745 -41332 -28530 -41268
rect -28466 -41332 -28446 -41268
rect -34745 -41348 -28446 -41332
rect -34745 -41412 -28530 -41348
rect -28466 -41412 -28446 -41348
rect -34745 -41428 -28446 -41412
rect -34745 -41492 -28530 -41428
rect -28466 -41492 -28446 -41428
rect -34745 -41508 -28446 -41492
rect -34745 -41572 -28530 -41508
rect -28466 -41572 -28446 -41508
rect -34745 -41588 -28446 -41572
rect -34745 -41652 -28530 -41588
rect -28466 -41652 -28446 -41588
rect -34745 -41668 -28446 -41652
rect -34745 -41732 -28530 -41668
rect -28466 -41732 -28446 -41668
rect -34745 -41748 -28446 -41732
rect -34745 -41812 -28530 -41748
rect -28466 -41812 -28446 -41748
rect -34745 -41828 -28446 -41812
rect -34745 -41892 -28530 -41828
rect -28466 -41892 -28446 -41828
rect -34745 -41908 -28446 -41892
rect -34745 -41972 -28530 -41908
rect -28466 -41972 -28446 -41908
rect -34745 -41988 -28446 -41972
rect -34745 -42052 -28530 -41988
rect -28466 -42052 -28446 -41988
rect -34745 -42068 -28446 -42052
rect -34745 -42132 -28530 -42068
rect -28466 -42132 -28446 -42068
rect -34745 -42148 -28446 -42132
rect -34745 -42212 -28530 -42148
rect -28466 -42212 -28446 -42148
rect -34745 -42228 -28446 -42212
rect -34745 -42292 -28530 -42228
rect -28466 -42292 -28446 -42228
rect -34745 -42308 -28446 -42292
rect -34745 -42372 -28530 -42308
rect -28466 -42372 -28446 -42308
rect -34745 -42388 -28446 -42372
rect -34745 -42452 -28530 -42388
rect -28466 -42452 -28446 -42388
rect -34745 -42468 -28446 -42452
rect -34745 -42532 -28530 -42468
rect -28466 -42532 -28446 -42468
rect -34745 -42548 -28446 -42532
rect -34745 -42612 -28530 -42548
rect -28466 -42612 -28446 -42548
rect -34745 -42628 -28446 -42612
rect -34745 -42692 -28530 -42628
rect -28466 -42692 -28446 -42628
rect -34745 -42708 -28446 -42692
rect -34745 -42772 -28530 -42708
rect -28466 -42772 -28446 -42708
rect -34745 -42788 -28446 -42772
rect -34745 -42852 -28530 -42788
rect -28466 -42852 -28446 -42788
rect -34745 -42868 -28446 -42852
rect -34745 -42932 -28530 -42868
rect -28466 -42932 -28446 -42868
rect -34745 -42948 -28446 -42932
rect -34745 -43012 -28530 -42948
rect -28466 -43012 -28446 -42948
rect -34745 -43028 -28446 -43012
rect -34745 -43092 -28530 -43028
rect -28466 -43092 -28446 -43028
rect -34745 -43108 -28446 -43092
rect -34745 -43172 -28530 -43108
rect -28466 -43172 -28446 -43108
rect -34745 -43188 -28446 -43172
rect -34745 -43252 -28530 -43188
rect -28466 -43252 -28446 -43188
rect -34745 -43268 -28446 -43252
rect -34745 -43332 -28530 -43268
rect -28466 -43332 -28446 -43268
rect -34745 -43348 -28446 -43332
rect -34745 -43412 -28530 -43348
rect -28466 -43412 -28446 -43348
rect -34745 -43428 -28446 -43412
rect -34745 -43492 -28530 -43428
rect -28466 -43492 -28446 -43428
rect -34745 -43508 -28446 -43492
rect -34745 -43572 -28530 -43508
rect -28466 -43572 -28446 -43508
rect -34745 -43588 -28446 -43572
rect -34745 -43652 -28530 -43588
rect -28466 -43652 -28446 -43588
rect -34745 -43668 -28446 -43652
rect -34745 -43732 -28530 -43668
rect -28466 -43732 -28446 -43668
rect -34745 -43748 -28446 -43732
rect -34745 -43812 -28530 -43748
rect -28466 -43812 -28446 -43748
rect -34745 -43828 -28446 -43812
rect -34745 -43892 -28530 -43828
rect -28466 -43892 -28446 -43828
rect -34745 -43908 -28446 -43892
rect -34745 -43972 -28530 -43908
rect -28466 -43972 -28446 -43908
rect -34745 -43988 -28446 -43972
rect -34745 -44052 -28530 -43988
rect -28466 -44052 -28446 -43988
rect -34745 -44068 -28446 -44052
rect -34745 -44132 -28530 -44068
rect -28466 -44132 -28446 -44068
rect -34745 -44148 -28446 -44132
rect -34745 -44212 -28530 -44148
rect -28466 -44212 -28446 -44148
rect -34745 -44228 -28446 -44212
rect -34745 -44292 -28530 -44228
rect -28466 -44292 -28446 -44228
rect -34745 -44308 -28446 -44292
rect -34745 -44372 -28530 -44308
rect -28466 -44372 -28446 -44308
rect -34745 -44388 -28446 -44372
rect -34745 -44452 -28530 -44388
rect -28466 -44452 -28446 -44388
rect -34745 -44468 -28446 -44452
rect -34745 -44532 -28530 -44468
rect -28466 -44532 -28446 -44468
rect -34745 -44548 -28446 -44532
rect -34745 -44612 -28530 -44548
rect -28466 -44612 -28446 -44548
rect -34745 -44628 -28446 -44612
rect -34745 -44692 -28530 -44628
rect -28466 -44692 -28446 -44628
rect -34745 -44708 -28446 -44692
rect -34745 -44772 -28530 -44708
rect -28466 -44772 -28446 -44708
rect -34745 -44788 -28446 -44772
rect -34745 -44852 -28530 -44788
rect -28466 -44852 -28446 -44788
rect -34745 -44868 -28446 -44852
rect -34745 -44932 -28530 -44868
rect -28466 -44932 -28446 -44868
rect -34745 -44948 -28446 -44932
rect -34745 -45012 -28530 -44948
rect -28466 -45012 -28446 -44948
rect -34745 -45028 -28446 -45012
rect -34745 -45092 -28530 -45028
rect -28466 -45092 -28446 -45028
rect -34745 -45108 -28446 -45092
rect -34745 -45172 -28530 -45108
rect -28466 -45172 -28446 -45108
rect -34745 -45188 -28446 -45172
rect -34745 -45252 -28530 -45188
rect -28466 -45252 -28446 -45188
rect -34745 -45268 -28446 -45252
rect -34745 -45332 -28530 -45268
rect -28466 -45332 -28446 -45268
rect -34745 -45348 -28446 -45332
rect -34745 -45412 -28530 -45348
rect -28466 -45412 -28446 -45348
rect -34745 -45428 -28446 -45412
rect -34745 -45492 -28530 -45428
rect -28466 -45492 -28446 -45428
rect -34745 -45508 -28446 -45492
rect -34745 -45572 -28530 -45508
rect -28466 -45572 -28446 -45508
rect -34745 -45588 -28446 -45572
rect -34745 -45652 -28530 -45588
rect -28466 -45652 -28446 -45588
rect -34745 -45668 -28446 -45652
rect -34745 -45732 -28530 -45668
rect -28466 -45732 -28446 -45668
rect -34745 -45748 -28446 -45732
rect -34745 -45812 -28530 -45748
rect -28466 -45812 -28446 -45748
rect -34745 -45828 -28446 -45812
rect -34745 -45892 -28530 -45828
rect -28466 -45892 -28446 -45828
rect -34745 -45908 -28446 -45892
rect -34745 -45972 -28530 -45908
rect -28466 -45972 -28446 -45908
rect -34745 -45988 -28446 -45972
rect -34745 -46052 -28530 -45988
rect -28466 -46052 -28446 -45988
rect -34745 -46068 -28446 -46052
rect -34745 -46132 -28530 -46068
rect -28466 -46132 -28446 -46068
rect -34745 -46148 -28446 -46132
rect -34745 -46212 -28530 -46148
rect -28466 -46212 -28446 -46148
rect -34745 -46228 -28446 -46212
rect -34745 -46292 -28530 -46228
rect -28466 -46292 -28446 -46228
rect -34745 -46308 -28446 -46292
rect -34745 -46372 -28530 -46308
rect -28466 -46372 -28446 -46308
rect -34745 -46388 -28446 -46372
rect -34745 -46452 -28530 -46388
rect -28466 -46452 -28446 -46388
rect -34745 -46468 -28446 -46452
rect -34745 -46532 -28530 -46468
rect -28466 -46532 -28446 -46468
rect -34745 -46548 -28446 -46532
rect -34745 -46612 -28530 -46548
rect -28466 -46612 -28446 -46548
rect -34745 -46628 -28446 -46612
rect -34745 -46692 -28530 -46628
rect -28466 -46692 -28446 -46628
rect -34745 -46708 -28446 -46692
rect -34745 -46772 -28530 -46708
rect -28466 -46772 -28446 -46708
rect -34745 -46788 -28446 -46772
rect -34745 -46852 -28530 -46788
rect -28466 -46852 -28446 -46788
rect -34745 -46868 -28446 -46852
rect -34745 -46932 -28530 -46868
rect -28466 -46932 -28446 -46868
rect -34745 -46948 -28446 -46932
rect -34745 -47012 -28530 -46948
rect -28466 -47012 -28446 -46948
rect -34745 -47028 -28446 -47012
rect -34745 -47092 -28530 -47028
rect -28466 -47092 -28446 -47028
rect -34745 -47108 -28446 -47092
rect -34745 -47172 -28530 -47108
rect -28466 -47172 -28446 -47108
rect -34745 -47200 -28446 -47172
rect -28426 -41028 -22127 -41000
rect -28426 -41092 -22211 -41028
rect -22147 -41092 -22127 -41028
rect -28426 -41108 -22127 -41092
rect -28426 -41172 -22211 -41108
rect -22147 -41172 -22127 -41108
rect -28426 -41188 -22127 -41172
rect -28426 -41252 -22211 -41188
rect -22147 -41252 -22127 -41188
rect -28426 -41268 -22127 -41252
rect -28426 -41332 -22211 -41268
rect -22147 -41332 -22127 -41268
rect -28426 -41348 -22127 -41332
rect -28426 -41412 -22211 -41348
rect -22147 -41412 -22127 -41348
rect -28426 -41428 -22127 -41412
rect -28426 -41492 -22211 -41428
rect -22147 -41492 -22127 -41428
rect -28426 -41508 -22127 -41492
rect -28426 -41572 -22211 -41508
rect -22147 -41572 -22127 -41508
rect -28426 -41588 -22127 -41572
rect -28426 -41652 -22211 -41588
rect -22147 -41652 -22127 -41588
rect -28426 -41668 -22127 -41652
rect -28426 -41732 -22211 -41668
rect -22147 -41732 -22127 -41668
rect -28426 -41748 -22127 -41732
rect -28426 -41812 -22211 -41748
rect -22147 -41812 -22127 -41748
rect -28426 -41828 -22127 -41812
rect -28426 -41892 -22211 -41828
rect -22147 -41892 -22127 -41828
rect -28426 -41908 -22127 -41892
rect -28426 -41972 -22211 -41908
rect -22147 -41972 -22127 -41908
rect -28426 -41988 -22127 -41972
rect -28426 -42052 -22211 -41988
rect -22147 -42052 -22127 -41988
rect -28426 -42068 -22127 -42052
rect -28426 -42132 -22211 -42068
rect -22147 -42132 -22127 -42068
rect -28426 -42148 -22127 -42132
rect -28426 -42212 -22211 -42148
rect -22147 -42212 -22127 -42148
rect -28426 -42228 -22127 -42212
rect -28426 -42292 -22211 -42228
rect -22147 -42292 -22127 -42228
rect -28426 -42308 -22127 -42292
rect -28426 -42372 -22211 -42308
rect -22147 -42372 -22127 -42308
rect -28426 -42388 -22127 -42372
rect -28426 -42452 -22211 -42388
rect -22147 -42452 -22127 -42388
rect -28426 -42468 -22127 -42452
rect -28426 -42532 -22211 -42468
rect -22147 -42532 -22127 -42468
rect -28426 -42548 -22127 -42532
rect -28426 -42612 -22211 -42548
rect -22147 -42612 -22127 -42548
rect -28426 -42628 -22127 -42612
rect -28426 -42692 -22211 -42628
rect -22147 -42692 -22127 -42628
rect -28426 -42708 -22127 -42692
rect -28426 -42772 -22211 -42708
rect -22147 -42772 -22127 -42708
rect -28426 -42788 -22127 -42772
rect -28426 -42852 -22211 -42788
rect -22147 -42852 -22127 -42788
rect -28426 -42868 -22127 -42852
rect -28426 -42932 -22211 -42868
rect -22147 -42932 -22127 -42868
rect -28426 -42948 -22127 -42932
rect -28426 -43012 -22211 -42948
rect -22147 -43012 -22127 -42948
rect -28426 -43028 -22127 -43012
rect -28426 -43092 -22211 -43028
rect -22147 -43092 -22127 -43028
rect -28426 -43108 -22127 -43092
rect -28426 -43172 -22211 -43108
rect -22147 -43172 -22127 -43108
rect -28426 -43188 -22127 -43172
rect -28426 -43252 -22211 -43188
rect -22147 -43252 -22127 -43188
rect -28426 -43268 -22127 -43252
rect -28426 -43332 -22211 -43268
rect -22147 -43332 -22127 -43268
rect -28426 -43348 -22127 -43332
rect -28426 -43412 -22211 -43348
rect -22147 -43412 -22127 -43348
rect -28426 -43428 -22127 -43412
rect -28426 -43492 -22211 -43428
rect -22147 -43492 -22127 -43428
rect -28426 -43508 -22127 -43492
rect -28426 -43572 -22211 -43508
rect -22147 -43572 -22127 -43508
rect -28426 -43588 -22127 -43572
rect -28426 -43652 -22211 -43588
rect -22147 -43652 -22127 -43588
rect -28426 -43668 -22127 -43652
rect -28426 -43732 -22211 -43668
rect -22147 -43732 -22127 -43668
rect -28426 -43748 -22127 -43732
rect -28426 -43812 -22211 -43748
rect -22147 -43812 -22127 -43748
rect -28426 -43828 -22127 -43812
rect -28426 -43892 -22211 -43828
rect -22147 -43892 -22127 -43828
rect -28426 -43908 -22127 -43892
rect -28426 -43972 -22211 -43908
rect -22147 -43972 -22127 -43908
rect -28426 -43988 -22127 -43972
rect -28426 -44052 -22211 -43988
rect -22147 -44052 -22127 -43988
rect -28426 -44068 -22127 -44052
rect -28426 -44132 -22211 -44068
rect -22147 -44132 -22127 -44068
rect -28426 -44148 -22127 -44132
rect -28426 -44212 -22211 -44148
rect -22147 -44212 -22127 -44148
rect -28426 -44228 -22127 -44212
rect -28426 -44292 -22211 -44228
rect -22147 -44292 -22127 -44228
rect -28426 -44308 -22127 -44292
rect -28426 -44372 -22211 -44308
rect -22147 -44372 -22127 -44308
rect -28426 -44388 -22127 -44372
rect -28426 -44452 -22211 -44388
rect -22147 -44452 -22127 -44388
rect -28426 -44468 -22127 -44452
rect -28426 -44532 -22211 -44468
rect -22147 -44532 -22127 -44468
rect -28426 -44548 -22127 -44532
rect -28426 -44612 -22211 -44548
rect -22147 -44612 -22127 -44548
rect -28426 -44628 -22127 -44612
rect -28426 -44692 -22211 -44628
rect -22147 -44692 -22127 -44628
rect -28426 -44708 -22127 -44692
rect -28426 -44772 -22211 -44708
rect -22147 -44772 -22127 -44708
rect -28426 -44788 -22127 -44772
rect -28426 -44852 -22211 -44788
rect -22147 -44852 -22127 -44788
rect -28426 -44868 -22127 -44852
rect -28426 -44932 -22211 -44868
rect -22147 -44932 -22127 -44868
rect -28426 -44948 -22127 -44932
rect -28426 -45012 -22211 -44948
rect -22147 -45012 -22127 -44948
rect -28426 -45028 -22127 -45012
rect -28426 -45092 -22211 -45028
rect -22147 -45092 -22127 -45028
rect -28426 -45108 -22127 -45092
rect -28426 -45172 -22211 -45108
rect -22147 -45172 -22127 -45108
rect -28426 -45188 -22127 -45172
rect -28426 -45252 -22211 -45188
rect -22147 -45252 -22127 -45188
rect -28426 -45268 -22127 -45252
rect -28426 -45332 -22211 -45268
rect -22147 -45332 -22127 -45268
rect -28426 -45348 -22127 -45332
rect -28426 -45412 -22211 -45348
rect -22147 -45412 -22127 -45348
rect -28426 -45428 -22127 -45412
rect -28426 -45492 -22211 -45428
rect -22147 -45492 -22127 -45428
rect -28426 -45508 -22127 -45492
rect -28426 -45572 -22211 -45508
rect -22147 -45572 -22127 -45508
rect -28426 -45588 -22127 -45572
rect -28426 -45652 -22211 -45588
rect -22147 -45652 -22127 -45588
rect -28426 -45668 -22127 -45652
rect -28426 -45732 -22211 -45668
rect -22147 -45732 -22127 -45668
rect -28426 -45748 -22127 -45732
rect -28426 -45812 -22211 -45748
rect -22147 -45812 -22127 -45748
rect -28426 -45828 -22127 -45812
rect -28426 -45892 -22211 -45828
rect -22147 -45892 -22127 -45828
rect -28426 -45908 -22127 -45892
rect -28426 -45972 -22211 -45908
rect -22147 -45972 -22127 -45908
rect -28426 -45988 -22127 -45972
rect -28426 -46052 -22211 -45988
rect -22147 -46052 -22127 -45988
rect -28426 -46068 -22127 -46052
rect -28426 -46132 -22211 -46068
rect -22147 -46132 -22127 -46068
rect -28426 -46148 -22127 -46132
rect -28426 -46212 -22211 -46148
rect -22147 -46212 -22127 -46148
rect -28426 -46228 -22127 -46212
rect -28426 -46292 -22211 -46228
rect -22147 -46292 -22127 -46228
rect -28426 -46308 -22127 -46292
rect -28426 -46372 -22211 -46308
rect -22147 -46372 -22127 -46308
rect -28426 -46388 -22127 -46372
rect -28426 -46452 -22211 -46388
rect -22147 -46452 -22127 -46388
rect -28426 -46468 -22127 -46452
rect -28426 -46532 -22211 -46468
rect -22147 -46532 -22127 -46468
rect -28426 -46548 -22127 -46532
rect -28426 -46612 -22211 -46548
rect -22147 -46612 -22127 -46548
rect -28426 -46628 -22127 -46612
rect -28426 -46692 -22211 -46628
rect -22147 -46692 -22127 -46628
rect -28426 -46708 -22127 -46692
rect -28426 -46772 -22211 -46708
rect -22147 -46772 -22127 -46708
rect -28426 -46788 -22127 -46772
rect -28426 -46852 -22211 -46788
rect -22147 -46852 -22127 -46788
rect -28426 -46868 -22127 -46852
rect -28426 -46932 -22211 -46868
rect -22147 -46932 -22127 -46868
rect -28426 -46948 -22127 -46932
rect -28426 -47012 -22211 -46948
rect -22147 -47012 -22127 -46948
rect -28426 -47028 -22127 -47012
rect -28426 -47092 -22211 -47028
rect -22147 -47092 -22127 -47028
rect -28426 -47108 -22127 -47092
rect -28426 -47172 -22211 -47108
rect -22147 -47172 -22127 -47108
rect -28426 -47200 -22127 -47172
rect -22107 -41028 -15808 -41000
rect -22107 -41092 -15892 -41028
rect -15828 -41092 -15808 -41028
rect -22107 -41108 -15808 -41092
rect -22107 -41172 -15892 -41108
rect -15828 -41172 -15808 -41108
rect -22107 -41188 -15808 -41172
rect -22107 -41252 -15892 -41188
rect -15828 -41252 -15808 -41188
rect -22107 -41268 -15808 -41252
rect -22107 -41332 -15892 -41268
rect -15828 -41332 -15808 -41268
rect -22107 -41348 -15808 -41332
rect -22107 -41412 -15892 -41348
rect -15828 -41412 -15808 -41348
rect -22107 -41428 -15808 -41412
rect -22107 -41492 -15892 -41428
rect -15828 -41492 -15808 -41428
rect -22107 -41508 -15808 -41492
rect -22107 -41572 -15892 -41508
rect -15828 -41572 -15808 -41508
rect -22107 -41588 -15808 -41572
rect -22107 -41652 -15892 -41588
rect -15828 -41652 -15808 -41588
rect -22107 -41668 -15808 -41652
rect -22107 -41732 -15892 -41668
rect -15828 -41732 -15808 -41668
rect -22107 -41748 -15808 -41732
rect -22107 -41812 -15892 -41748
rect -15828 -41812 -15808 -41748
rect -22107 -41828 -15808 -41812
rect -22107 -41892 -15892 -41828
rect -15828 -41892 -15808 -41828
rect -22107 -41908 -15808 -41892
rect -22107 -41972 -15892 -41908
rect -15828 -41972 -15808 -41908
rect -22107 -41988 -15808 -41972
rect -22107 -42052 -15892 -41988
rect -15828 -42052 -15808 -41988
rect -22107 -42068 -15808 -42052
rect -22107 -42132 -15892 -42068
rect -15828 -42132 -15808 -42068
rect -22107 -42148 -15808 -42132
rect -22107 -42212 -15892 -42148
rect -15828 -42212 -15808 -42148
rect -22107 -42228 -15808 -42212
rect -22107 -42292 -15892 -42228
rect -15828 -42292 -15808 -42228
rect -22107 -42308 -15808 -42292
rect -22107 -42372 -15892 -42308
rect -15828 -42372 -15808 -42308
rect -22107 -42388 -15808 -42372
rect -22107 -42452 -15892 -42388
rect -15828 -42452 -15808 -42388
rect -22107 -42468 -15808 -42452
rect -22107 -42532 -15892 -42468
rect -15828 -42532 -15808 -42468
rect -22107 -42548 -15808 -42532
rect -22107 -42612 -15892 -42548
rect -15828 -42612 -15808 -42548
rect -22107 -42628 -15808 -42612
rect -22107 -42692 -15892 -42628
rect -15828 -42692 -15808 -42628
rect -22107 -42708 -15808 -42692
rect -22107 -42772 -15892 -42708
rect -15828 -42772 -15808 -42708
rect -22107 -42788 -15808 -42772
rect -22107 -42852 -15892 -42788
rect -15828 -42852 -15808 -42788
rect -22107 -42868 -15808 -42852
rect -22107 -42932 -15892 -42868
rect -15828 -42932 -15808 -42868
rect -22107 -42948 -15808 -42932
rect -22107 -43012 -15892 -42948
rect -15828 -43012 -15808 -42948
rect -22107 -43028 -15808 -43012
rect -22107 -43092 -15892 -43028
rect -15828 -43092 -15808 -43028
rect -22107 -43108 -15808 -43092
rect -22107 -43172 -15892 -43108
rect -15828 -43172 -15808 -43108
rect -22107 -43188 -15808 -43172
rect -22107 -43252 -15892 -43188
rect -15828 -43252 -15808 -43188
rect -22107 -43268 -15808 -43252
rect -22107 -43332 -15892 -43268
rect -15828 -43332 -15808 -43268
rect -22107 -43348 -15808 -43332
rect -22107 -43412 -15892 -43348
rect -15828 -43412 -15808 -43348
rect -22107 -43428 -15808 -43412
rect -22107 -43492 -15892 -43428
rect -15828 -43492 -15808 -43428
rect -22107 -43508 -15808 -43492
rect -22107 -43572 -15892 -43508
rect -15828 -43572 -15808 -43508
rect -22107 -43588 -15808 -43572
rect -22107 -43652 -15892 -43588
rect -15828 -43652 -15808 -43588
rect -22107 -43668 -15808 -43652
rect -22107 -43732 -15892 -43668
rect -15828 -43732 -15808 -43668
rect -22107 -43748 -15808 -43732
rect -22107 -43812 -15892 -43748
rect -15828 -43812 -15808 -43748
rect -22107 -43828 -15808 -43812
rect -22107 -43892 -15892 -43828
rect -15828 -43892 -15808 -43828
rect -22107 -43908 -15808 -43892
rect -22107 -43972 -15892 -43908
rect -15828 -43972 -15808 -43908
rect -22107 -43988 -15808 -43972
rect -22107 -44052 -15892 -43988
rect -15828 -44052 -15808 -43988
rect -22107 -44068 -15808 -44052
rect -22107 -44132 -15892 -44068
rect -15828 -44132 -15808 -44068
rect -22107 -44148 -15808 -44132
rect -22107 -44212 -15892 -44148
rect -15828 -44212 -15808 -44148
rect -22107 -44228 -15808 -44212
rect -22107 -44292 -15892 -44228
rect -15828 -44292 -15808 -44228
rect -22107 -44308 -15808 -44292
rect -22107 -44372 -15892 -44308
rect -15828 -44372 -15808 -44308
rect -22107 -44388 -15808 -44372
rect -22107 -44452 -15892 -44388
rect -15828 -44452 -15808 -44388
rect -22107 -44468 -15808 -44452
rect -22107 -44532 -15892 -44468
rect -15828 -44532 -15808 -44468
rect -22107 -44548 -15808 -44532
rect -22107 -44612 -15892 -44548
rect -15828 -44612 -15808 -44548
rect -22107 -44628 -15808 -44612
rect -22107 -44692 -15892 -44628
rect -15828 -44692 -15808 -44628
rect -22107 -44708 -15808 -44692
rect -22107 -44772 -15892 -44708
rect -15828 -44772 -15808 -44708
rect -22107 -44788 -15808 -44772
rect -22107 -44852 -15892 -44788
rect -15828 -44852 -15808 -44788
rect -22107 -44868 -15808 -44852
rect -22107 -44932 -15892 -44868
rect -15828 -44932 -15808 -44868
rect -22107 -44948 -15808 -44932
rect -22107 -45012 -15892 -44948
rect -15828 -45012 -15808 -44948
rect -22107 -45028 -15808 -45012
rect -22107 -45092 -15892 -45028
rect -15828 -45092 -15808 -45028
rect -22107 -45108 -15808 -45092
rect -22107 -45172 -15892 -45108
rect -15828 -45172 -15808 -45108
rect -22107 -45188 -15808 -45172
rect -22107 -45252 -15892 -45188
rect -15828 -45252 -15808 -45188
rect -22107 -45268 -15808 -45252
rect -22107 -45332 -15892 -45268
rect -15828 -45332 -15808 -45268
rect -22107 -45348 -15808 -45332
rect -22107 -45412 -15892 -45348
rect -15828 -45412 -15808 -45348
rect -22107 -45428 -15808 -45412
rect -22107 -45492 -15892 -45428
rect -15828 -45492 -15808 -45428
rect -22107 -45508 -15808 -45492
rect -22107 -45572 -15892 -45508
rect -15828 -45572 -15808 -45508
rect -22107 -45588 -15808 -45572
rect -22107 -45652 -15892 -45588
rect -15828 -45652 -15808 -45588
rect -22107 -45668 -15808 -45652
rect -22107 -45732 -15892 -45668
rect -15828 -45732 -15808 -45668
rect -22107 -45748 -15808 -45732
rect -22107 -45812 -15892 -45748
rect -15828 -45812 -15808 -45748
rect -22107 -45828 -15808 -45812
rect -22107 -45892 -15892 -45828
rect -15828 -45892 -15808 -45828
rect -22107 -45908 -15808 -45892
rect -22107 -45972 -15892 -45908
rect -15828 -45972 -15808 -45908
rect -22107 -45988 -15808 -45972
rect -22107 -46052 -15892 -45988
rect -15828 -46052 -15808 -45988
rect -22107 -46068 -15808 -46052
rect -22107 -46132 -15892 -46068
rect -15828 -46132 -15808 -46068
rect -22107 -46148 -15808 -46132
rect -22107 -46212 -15892 -46148
rect -15828 -46212 -15808 -46148
rect -22107 -46228 -15808 -46212
rect -22107 -46292 -15892 -46228
rect -15828 -46292 -15808 -46228
rect -22107 -46308 -15808 -46292
rect -22107 -46372 -15892 -46308
rect -15828 -46372 -15808 -46308
rect -22107 -46388 -15808 -46372
rect -22107 -46452 -15892 -46388
rect -15828 -46452 -15808 -46388
rect -22107 -46468 -15808 -46452
rect -22107 -46532 -15892 -46468
rect -15828 -46532 -15808 -46468
rect -22107 -46548 -15808 -46532
rect -22107 -46612 -15892 -46548
rect -15828 -46612 -15808 -46548
rect -22107 -46628 -15808 -46612
rect -22107 -46692 -15892 -46628
rect -15828 -46692 -15808 -46628
rect -22107 -46708 -15808 -46692
rect -22107 -46772 -15892 -46708
rect -15828 -46772 -15808 -46708
rect -22107 -46788 -15808 -46772
rect -22107 -46852 -15892 -46788
rect -15828 -46852 -15808 -46788
rect -22107 -46868 -15808 -46852
rect -22107 -46932 -15892 -46868
rect -15828 -46932 -15808 -46868
rect -22107 -46948 -15808 -46932
rect -22107 -47012 -15892 -46948
rect -15828 -47012 -15808 -46948
rect -22107 -47028 -15808 -47012
rect -22107 -47092 -15892 -47028
rect -15828 -47092 -15808 -47028
rect -22107 -47108 -15808 -47092
rect -22107 -47172 -15892 -47108
rect -15828 -47172 -15808 -47108
rect -22107 -47200 -15808 -47172
rect -15788 -41028 -9489 -41000
rect -15788 -41092 -9573 -41028
rect -9509 -41092 -9489 -41028
rect -15788 -41108 -9489 -41092
rect -15788 -41172 -9573 -41108
rect -9509 -41172 -9489 -41108
rect -15788 -41188 -9489 -41172
rect -15788 -41252 -9573 -41188
rect -9509 -41252 -9489 -41188
rect -15788 -41268 -9489 -41252
rect -15788 -41332 -9573 -41268
rect -9509 -41332 -9489 -41268
rect -15788 -41348 -9489 -41332
rect -15788 -41412 -9573 -41348
rect -9509 -41412 -9489 -41348
rect -15788 -41428 -9489 -41412
rect -15788 -41492 -9573 -41428
rect -9509 -41492 -9489 -41428
rect -15788 -41508 -9489 -41492
rect -15788 -41572 -9573 -41508
rect -9509 -41572 -9489 -41508
rect -15788 -41588 -9489 -41572
rect -15788 -41652 -9573 -41588
rect -9509 -41652 -9489 -41588
rect -15788 -41668 -9489 -41652
rect -15788 -41732 -9573 -41668
rect -9509 -41732 -9489 -41668
rect -15788 -41748 -9489 -41732
rect -15788 -41812 -9573 -41748
rect -9509 -41812 -9489 -41748
rect -15788 -41828 -9489 -41812
rect -15788 -41892 -9573 -41828
rect -9509 -41892 -9489 -41828
rect -15788 -41908 -9489 -41892
rect -15788 -41972 -9573 -41908
rect -9509 -41972 -9489 -41908
rect -15788 -41988 -9489 -41972
rect -15788 -42052 -9573 -41988
rect -9509 -42052 -9489 -41988
rect -15788 -42068 -9489 -42052
rect -15788 -42132 -9573 -42068
rect -9509 -42132 -9489 -42068
rect -15788 -42148 -9489 -42132
rect -15788 -42212 -9573 -42148
rect -9509 -42212 -9489 -42148
rect -15788 -42228 -9489 -42212
rect -15788 -42292 -9573 -42228
rect -9509 -42292 -9489 -42228
rect -15788 -42308 -9489 -42292
rect -15788 -42372 -9573 -42308
rect -9509 -42372 -9489 -42308
rect -15788 -42388 -9489 -42372
rect -15788 -42452 -9573 -42388
rect -9509 -42452 -9489 -42388
rect -15788 -42468 -9489 -42452
rect -15788 -42532 -9573 -42468
rect -9509 -42532 -9489 -42468
rect -15788 -42548 -9489 -42532
rect -15788 -42612 -9573 -42548
rect -9509 -42612 -9489 -42548
rect -15788 -42628 -9489 -42612
rect -15788 -42692 -9573 -42628
rect -9509 -42692 -9489 -42628
rect -15788 -42708 -9489 -42692
rect -15788 -42772 -9573 -42708
rect -9509 -42772 -9489 -42708
rect -15788 -42788 -9489 -42772
rect -15788 -42852 -9573 -42788
rect -9509 -42852 -9489 -42788
rect -15788 -42868 -9489 -42852
rect -15788 -42932 -9573 -42868
rect -9509 -42932 -9489 -42868
rect -15788 -42948 -9489 -42932
rect -15788 -43012 -9573 -42948
rect -9509 -43012 -9489 -42948
rect -15788 -43028 -9489 -43012
rect -15788 -43092 -9573 -43028
rect -9509 -43092 -9489 -43028
rect -15788 -43108 -9489 -43092
rect -15788 -43172 -9573 -43108
rect -9509 -43172 -9489 -43108
rect -15788 -43188 -9489 -43172
rect -15788 -43252 -9573 -43188
rect -9509 -43252 -9489 -43188
rect -15788 -43268 -9489 -43252
rect -15788 -43332 -9573 -43268
rect -9509 -43332 -9489 -43268
rect -15788 -43348 -9489 -43332
rect -15788 -43412 -9573 -43348
rect -9509 -43412 -9489 -43348
rect -15788 -43428 -9489 -43412
rect -15788 -43492 -9573 -43428
rect -9509 -43492 -9489 -43428
rect -15788 -43508 -9489 -43492
rect -15788 -43572 -9573 -43508
rect -9509 -43572 -9489 -43508
rect -15788 -43588 -9489 -43572
rect -15788 -43652 -9573 -43588
rect -9509 -43652 -9489 -43588
rect -15788 -43668 -9489 -43652
rect -15788 -43732 -9573 -43668
rect -9509 -43732 -9489 -43668
rect -15788 -43748 -9489 -43732
rect -15788 -43812 -9573 -43748
rect -9509 -43812 -9489 -43748
rect -15788 -43828 -9489 -43812
rect -15788 -43892 -9573 -43828
rect -9509 -43892 -9489 -43828
rect -15788 -43908 -9489 -43892
rect -15788 -43972 -9573 -43908
rect -9509 -43972 -9489 -43908
rect -15788 -43988 -9489 -43972
rect -15788 -44052 -9573 -43988
rect -9509 -44052 -9489 -43988
rect -15788 -44068 -9489 -44052
rect -15788 -44132 -9573 -44068
rect -9509 -44132 -9489 -44068
rect -15788 -44148 -9489 -44132
rect -15788 -44212 -9573 -44148
rect -9509 -44212 -9489 -44148
rect -15788 -44228 -9489 -44212
rect -15788 -44292 -9573 -44228
rect -9509 -44292 -9489 -44228
rect -15788 -44308 -9489 -44292
rect -15788 -44372 -9573 -44308
rect -9509 -44372 -9489 -44308
rect -15788 -44388 -9489 -44372
rect -15788 -44452 -9573 -44388
rect -9509 -44452 -9489 -44388
rect -15788 -44468 -9489 -44452
rect -15788 -44532 -9573 -44468
rect -9509 -44532 -9489 -44468
rect -15788 -44548 -9489 -44532
rect -15788 -44612 -9573 -44548
rect -9509 -44612 -9489 -44548
rect -15788 -44628 -9489 -44612
rect -15788 -44692 -9573 -44628
rect -9509 -44692 -9489 -44628
rect -15788 -44708 -9489 -44692
rect -15788 -44772 -9573 -44708
rect -9509 -44772 -9489 -44708
rect -15788 -44788 -9489 -44772
rect -15788 -44852 -9573 -44788
rect -9509 -44852 -9489 -44788
rect -15788 -44868 -9489 -44852
rect -15788 -44932 -9573 -44868
rect -9509 -44932 -9489 -44868
rect -15788 -44948 -9489 -44932
rect -15788 -45012 -9573 -44948
rect -9509 -45012 -9489 -44948
rect -15788 -45028 -9489 -45012
rect -15788 -45092 -9573 -45028
rect -9509 -45092 -9489 -45028
rect -15788 -45108 -9489 -45092
rect -15788 -45172 -9573 -45108
rect -9509 -45172 -9489 -45108
rect -15788 -45188 -9489 -45172
rect -15788 -45252 -9573 -45188
rect -9509 -45252 -9489 -45188
rect -15788 -45268 -9489 -45252
rect -15788 -45332 -9573 -45268
rect -9509 -45332 -9489 -45268
rect -15788 -45348 -9489 -45332
rect -15788 -45412 -9573 -45348
rect -9509 -45412 -9489 -45348
rect -15788 -45428 -9489 -45412
rect -15788 -45492 -9573 -45428
rect -9509 -45492 -9489 -45428
rect -15788 -45508 -9489 -45492
rect -15788 -45572 -9573 -45508
rect -9509 -45572 -9489 -45508
rect -15788 -45588 -9489 -45572
rect -15788 -45652 -9573 -45588
rect -9509 -45652 -9489 -45588
rect -15788 -45668 -9489 -45652
rect -15788 -45732 -9573 -45668
rect -9509 -45732 -9489 -45668
rect -15788 -45748 -9489 -45732
rect -15788 -45812 -9573 -45748
rect -9509 -45812 -9489 -45748
rect -15788 -45828 -9489 -45812
rect -15788 -45892 -9573 -45828
rect -9509 -45892 -9489 -45828
rect -15788 -45908 -9489 -45892
rect -15788 -45972 -9573 -45908
rect -9509 -45972 -9489 -45908
rect -15788 -45988 -9489 -45972
rect -15788 -46052 -9573 -45988
rect -9509 -46052 -9489 -45988
rect -15788 -46068 -9489 -46052
rect -15788 -46132 -9573 -46068
rect -9509 -46132 -9489 -46068
rect -15788 -46148 -9489 -46132
rect -15788 -46212 -9573 -46148
rect -9509 -46212 -9489 -46148
rect -15788 -46228 -9489 -46212
rect -15788 -46292 -9573 -46228
rect -9509 -46292 -9489 -46228
rect -15788 -46308 -9489 -46292
rect -15788 -46372 -9573 -46308
rect -9509 -46372 -9489 -46308
rect -15788 -46388 -9489 -46372
rect -15788 -46452 -9573 -46388
rect -9509 -46452 -9489 -46388
rect -15788 -46468 -9489 -46452
rect -15788 -46532 -9573 -46468
rect -9509 -46532 -9489 -46468
rect -15788 -46548 -9489 -46532
rect -15788 -46612 -9573 -46548
rect -9509 -46612 -9489 -46548
rect -15788 -46628 -9489 -46612
rect -15788 -46692 -9573 -46628
rect -9509 -46692 -9489 -46628
rect -15788 -46708 -9489 -46692
rect -15788 -46772 -9573 -46708
rect -9509 -46772 -9489 -46708
rect -15788 -46788 -9489 -46772
rect -15788 -46852 -9573 -46788
rect -9509 -46852 -9489 -46788
rect -15788 -46868 -9489 -46852
rect -15788 -46932 -9573 -46868
rect -9509 -46932 -9489 -46868
rect -15788 -46948 -9489 -46932
rect -15788 -47012 -9573 -46948
rect -9509 -47012 -9489 -46948
rect -15788 -47028 -9489 -47012
rect -15788 -47092 -9573 -47028
rect -9509 -47092 -9489 -47028
rect -15788 -47108 -9489 -47092
rect -15788 -47172 -9573 -47108
rect -9509 -47172 -9489 -47108
rect -15788 -47200 -9489 -47172
rect -9469 -41028 -3170 -41000
rect -9469 -41092 -3254 -41028
rect -3190 -41092 -3170 -41028
rect -9469 -41108 -3170 -41092
rect -9469 -41172 -3254 -41108
rect -3190 -41172 -3170 -41108
rect -9469 -41188 -3170 -41172
rect -9469 -41252 -3254 -41188
rect -3190 -41252 -3170 -41188
rect -9469 -41268 -3170 -41252
rect -9469 -41332 -3254 -41268
rect -3190 -41332 -3170 -41268
rect -9469 -41348 -3170 -41332
rect -9469 -41412 -3254 -41348
rect -3190 -41412 -3170 -41348
rect -9469 -41428 -3170 -41412
rect -9469 -41492 -3254 -41428
rect -3190 -41492 -3170 -41428
rect -9469 -41508 -3170 -41492
rect -9469 -41572 -3254 -41508
rect -3190 -41572 -3170 -41508
rect -9469 -41588 -3170 -41572
rect -9469 -41652 -3254 -41588
rect -3190 -41652 -3170 -41588
rect -9469 -41668 -3170 -41652
rect -9469 -41732 -3254 -41668
rect -3190 -41732 -3170 -41668
rect -9469 -41748 -3170 -41732
rect -9469 -41812 -3254 -41748
rect -3190 -41812 -3170 -41748
rect -9469 -41828 -3170 -41812
rect -9469 -41892 -3254 -41828
rect -3190 -41892 -3170 -41828
rect -9469 -41908 -3170 -41892
rect -9469 -41972 -3254 -41908
rect -3190 -41972 -3170 -41908
rect -9469 -41988 -3170 -41972
rect -9469 -42052 -3254 -41988
rect -3190 -42052 -3170 -41988
rect -9469 -42068 -3170 -42052
rect -9469 -42132 -3254 -42068
rect -3190 -42132 -3170 -42068
rect -9469 -42148 -3170 -42132
rect -9469 -42212 -3254 -42148
rect -3190 -42212 -3170 -42148
rect -9469 -42228 -3170 -42212
rect -9469 -42292 -3254 -42228
rect -3190 -42292 -3170 -42228
rect -9469 -42308 -3170 -42292
rect -9469 -42372 -3254 -42308
rect -3190 -42372 -3170 -42308
rect -9469 -42388 -3170 -42372
rect -9469 -42452 -3254 -42388
rect -3190 -42452 -3170 -42388
rect -9469 -42468 -3170 -42452
rect -9469 -42532 -3254 -42468
rect -3190 -42532 -3170 -42468
rect -9469 -42548 -3170 -42532
rect -9469 -42612 -3254 -42548
rect -3190 -42612 -3170 -42548
rect -9469 -42628 -3170 -42612
rect -9469 -42692 -3254 -42628
rect -3190 -42692 -3170 -42628
rect -9469 -42708 -3170 -42692
rect -9469 -42772 -3254 -42708
rect -3190 -42772 -3170 -42708
rect -9469 -42788 -3170 -42772
rect -9469 -42852 -3254 -42788
rect -3190 -42852 -3170 -42788
rect -9469 -42868 -3170 -42852
rect -9469 -42932 -3254 -42868
rect -3190 -42932 -3170 -42868
rect -9469 -42948 -3170 -42932
rect -9469 -43012 -3254 -42948
rect -3190 -43012 -3170 -42948
rect -9469 -43028 -3170 -43012
rect -9469 -43092 -3254 -43028
rect -3190 -43092 -3170 -43028
rect -9469 -43108 -3170 -43092
rect -9469 -43172 -3254 -43108
rect -3190 -43172 -3170 -43108
rect -9469 -43188 -3170 -43172
rect -9469 -43252 -3254 -43188
rect -3190 -43252 -3170 -43188
rect -9469 -43268 -3170 -43252
rect -9469 -43332 -3254 -43268
rect -3190 -43332 -3170 -43268
rect -9469 -43348 -3170 -43332
rect -9469 -43412 -3254 -43348
rect -3190 -43412 -3170 -43348
rect -9469 -43428 -3170 -43412
rect -9469 -43492 -3254 -43428
rect -3190 -43492 -3170 -43428
rect -9469 -43508 -3170 -43492
rect -9469 -43572 -3254 -43508
rect -3190 -43572 -3170 -43508
rect -9469 -43588 -3170 -43572
rect -9469 -43652 -3254 -43588
rect -3190 -43652 -3170 -43588
rect -9469 -43668 -3170 -43652
rect -9469 -43732 -3254 -43668
rect -3190 -43732 -3170 -43668
rect -9469 -43748 -3170 -43732
rect -9469 -43812 -3254 -43748
rect -3190 -43812 -3170 -43748
rect -9469 -43828 -3170 -43812
rect -9469 -43892 -3254 -43828
rect -3190 -43892 -3170 -43828
rect -9469 -43908 -3170 -43892
rect -9469 -43972 -3254 -43908
rect -3190 -43972 -3170 -43908
rect -9469 -43988 -3170 -43972
rect -9469 -44052 -3254 -43988
rect -3190 -44052 -3170 -43988
rect -9469 -44068 -3170 -44052
rect -9469 -44132 -3254 -44068
rect -3190 -44132 -3170 -44068
rect -9469 -44148 -3170 -44132
rect -9469 -44212 -3254 -44148
rect -3190 -44212 -3170 -44148
rect -9469 -44228 -3170 -44212
rect -9469 -44292 -3254 -44228
rect -3190 -44292 -3170 -44228
rect -9469 -44308 -3170 -44292
rect -9469 -44372 -3254 -44308
rect -3190 -44372 -3170 -44308
rect -9469 -44388 -3170 -44372
rect -9469 -44452 -3254 -44388
rect -3190 -44452 -3170 -44388
rect -9469 -44468 -3170 -44452
rect -9469 -44532 -3254 -44468
rect -3190 -44532 -3170 -44468
rect -9469 -44548 -3170 -44532
rect -9469 -44612 -3254 -44548
rect -3190 -44612 -3170 -44548
rect -9469 -44628 -3170 -44612
rect -9469 -44692 -3254 -44628
rect -3190 -44692 -3170 -44628
rect -9469 -44708 -3170 -44692
rect -9469 -44772 -3254 -44708
rect -3190 -44772 -3170 -44708
rect -9469 -44788 -3170 -44772
rect -9469 -44852 -3254 -44788
rect -3190 -44852 -3170 -44788
rect -9469 -44868 -3170 -44852
rect -9469 -44932 -3254 -44868
rect -3190 -44932 -3170 -44868
rect -9469 -44948 -3170 -44932
rect -9469 -45012 -3254 -44948
rect -3190 -45012 -3170 -44948
rect -9469 -45028 -3170 -45012
rect -9469 -45092 -3254 -45028
rect -3190 -45092 -3170 -45028
rect -9469 -45108 -3170 -45092
rect -9469 -45172 -3254 -45108
rect -3190 -45172 -3170 -45108
rect -9469 -45188 -3170 -45172
rect -9469 -45252 -3254 -45188
rect -3190 -45252 -3170 -45188
rect -9469 -45268 -3170 -45252
rect -9469 -45332 -3254 -45268
rect -3190 -45332 -3170 -45268
rect -9469 -45348 -3170 -45332
rect -9469 -45412 -3254 -45348
rect -3190 -45412 -3170 -45348
rect -9469 -45428 -3170 -45412
rect -9469 -45492 -3254 -45428
rect -3190 -45492 -3170 -45428
rect -9469 -45508 -3170 -45492
rect -9469 -45572 -3254 -45508
rect -3190 -45572 -3170 -45508
rect -9469 -45588 -3170 -45572
rect -9469 -45652 -3254 -45588
rect -3190 -45652 -3170 -45588
rect -9469 -45668 -3170 -45652
rect -9469 -45732 -3254 -45668
rect -3190 -45732 -3170 -45668
rect -9469 -45748 -3170 -45732
rect -9469 -45812 -3254 -45748
rect -3190 -45812 -3170 -45748
rect -9469 -45828 -3170 -45812
rect -9469 -45892 -3254 -45828
rect -3190 -45892 -3170 -45828
rect -9469 -45908 -3170 -45892
rect -9469 -45972 -3254 -45908
rect -3190 -45972 -3170 -45908
rect -9469 -45988 -3170 -45972
rect -9469 -46052 -3254 -45988
rect -3190 -46052 -3170 -45988
rect -9469 -46068 -3170 -46052
rect -9469 -46132 -3254 -46068
rect -3190 -46132 -3170 -46068
rect -9469 -46148 -3170 -46132
rect -9469 -46212 -3254 -46148
rect -3190 -46212 -3170 -46148
rect -9469 -46228 -3170 -46212
rect -9469 -46292 -3254 -46228
rect -3190 -46292 -3170 -46228
rect -9469 -46308 -3170 -46292
rect -9469 -46372 -3254 -46308
rect -3190 -46372 -3170 -46308
rect -9469 -46388 -3170 -46372
rect -9469 -46452 -3254 -46388
rect -3190 -46452 -3170 -46388
rect -9469 -46468 -3170 -46452
rect -9469 -46532 -3254 -46468
rect -3190 -46532 -3170 -46468
rect -9469 -46548 -3170 -46532
rect -9469 -46612 -3254 -46548
rect -3190 -46612 -3170 -46548
rect -9469 -46628 -3170 -46612
rect -9469 -46692 -3254 -46628
rect -3190 -46692 -3170 -46628
rect -9469 -46708 -3170 -46692
rect -9469 -46772 -3254 -46708
rect -3190 -46772 -3170 -46708
rect -9469 -46788 -3170 -46772
rect -9469 -46852 -3254 -46788
rect -3190 -46852 -3170 -46788
rect -9469 -46868 -3170 -46852
rect -9469 -46932 -3254 -46868
rect -3190 -46932 -3170 -46868
rect -9469 -46948 -3170 -46932
rect -9469 -47012 -3254 -46948
rect -3190 -47012 -3170 -46948
rect -9469 -47028 -3170 -47012
rect -9469 -47092 -3254 -47028
rect -3190 -47092 -3170 -47028
rect -9469 -47108 -3170 -47092
rect -9469 -47172 -3254 -47108
rect -3190 -47172 -3170 -47108
rect -9469 -47200 -3170 -47172
rect -3150 -41028 3149 -41000
rect -3150 -41092 3065 -41028
rect 3129 -41092 3149 -41028
rect -3150 -41108 3149 -41092
rect -3150 -41172 3065 -41108
rect 3129 -41172 3149 -41108
rect -3150 -41188 3149 -41172
rect -3150 -41252 3065 -41188
rect 3129 -41252 3149 -41188
rect -3150 -41268 3149 -41252
rect -3150 -41332 3065 -41268
rect 3129 -41332 3149 -41268
rect -3150 -41348 3149 -41332
rect -3150 -41412 3065 -41348
rect 3129 -41412 3149 -41348
rect -3150 -41428 3149 -41412
rect -3150 -41492 3065 -41428
rect 3129 -41492 3149 -41428
rect -3150 -41508 3149 -41492
rect -3150 -41572 3065 -41508
rect 3129 -41572 3149 -41508
rect -3150 -41588 3149 -41572
rect -3150 -41652 3065 -41588
rect 3129 -41652 3149 -41588
rect -3150 -41668 3149 -41652
rect -3150 -41732 3065 -41668
rect 3129 -41732 3149 -41668
rect -3150 -41748 3149 -41732
rect -3150 -41812 3065 -41748
rect 3129 -41812 3149 -41748
rect -3150 -41828 3149 -41812
rect -3150 -41892 3065 -41828
rect 3129 -41892 3149 -41828
rect -3150 -41908 3149 -41892
rect -3150 -41972 3065 -41908
rect 3129 -41972 3149 -41908
rect -3150 -41988 3149 -41972
rect -3150 -42052 3065 -41988
rect 3129 -42052 3149 -41988
rect -3150 -42068 3149 -42052
rect -3150 -42132 3065 -42068
rect 3129 -42132 3149 -42068
rect -3150 -42148 3149 -42132
rect -3150 -42212 3065 -42148
rect 3129 -42212 3149 -42148
rect -3150 -42228 3149 -42212
rect -3150 -42292 3065 -42228
rect 3129 -42292 3149 -42228
rect -3150 -42308 3149 -42292
rect -3150 -42372 3065 -42308
rect 3129 -42372 3149 -42308
rect -3150 -42388 3149 -42372
rect -3150 -42452 3065 -42388
rect 3129 -42452 3149 -42388
rect -3150 -42468 3149 -42452
rect -3150 -42532 3065 -42468
rect 3129 -42532 3149 -42468
rect -3150 -42548 3149 -42532
rect -3150 -42612 3065 -42548
rect 3129 -42612 3149 -42548
rect -3150 -42628 3149 -42612
rect -3150 -42692 3065 -42628
rect 3129 -42692 3149 -42628
rect -3150 -42708 3149 -42692
rect -3150 -42772 3065 -42708
rect 3129 -42772 3149 -42708
rect -3150 -42788 3149 -42772
rect -3150 -42852 3065 -42788
rect 3129 -42852 3149 -42788
rect -3150 -42868 3149 -42852
rect -3150 -42932 3065 -42868
rect 3129 -42932 3149 -42868
rect -3150 -42948 3149 -42932
rect -3150 -43012 3065 -42948
rect 3129 -43012 3149 -42948
rect -3150 -43028 3149 -43012
rect -3150 -43092 3065 -43028
rect 3129 -43092 3149 -43028
rect -3150 -43108 3149 -43092
rect -3150 -43172 3065 -43108
rect 3129 -43172 3149 -43108
rect -3150 -43188 3149 -43172
rect -3150 -43252 3065 -43188
rect 3129 -43252 3149 -43188
rect -3150 -43268 3149 -43252
rect -3150 -43332 3065 -43268
rect 3129 -43332 3149 -43268
rect -3150 -43348 3149 -43332
rect -3150 -43412 3065 -43348
rect 3129 -43412 3149 -43348
rect -3150 -43428 3149 -43412
rect -3150 -43492 3065 -43428
rect 3129 -43492 3149 -43428
rect -3150 -43508 3149 -43492
rect -3150 -43572 3065 -43508
rect 3129 -43572 3149 -43508
rect -3150 -43588 3149 -43572
rect -3150 -43652 3065 -43588
rect 3129 -43652 3149 -43588
rect -3150 -43668 3149 -43652
rect -3150 -43732 3065 -43668
rect 3129 -43732 3149 -43668
rect -3150 -43748 3149 -43732
rect -3150 -43812 3065 -43748
rect 3129 -43812 3149 -43748
rect -3150 -43828 3149 -43812
rect -3150 -43892 3065 -43828
rect 3129 -43892 3149 -43828
rect -3150 -43908 3149 -43892
rect -3150 -43972 3065 -43908
rect 3129 -43972 3149 -43908
rect -3150 -43988 3149 -43972
rect -3150 -44052 3065 -43988
rect 3129 -44052 3149 -43988
rect -3150 -44068 3149 -44052
rect -3150 -44132 3065 -44068
rect 3129 -44132 3149 -44068
rect -3150 -44148 3149 -44132
rect -3150 -44212 3065 -44148
rect 3129 -44212 3149 -44148
rect -3150 -44228 3149 -44212
rect -3150 -44292 3065 -44228
rect 3129 -44292 3149 -44228
rect -3150 -44308 3149 -44292
rect -3150 -44372 3065 -44308
rect 3129 -44372 3149 -44308
rect -3150 -44388 3149 -44372
rect -3150 -44452 3065 -44388
rect 3129 -44452 3149 -44388
rect -3150 -44468 3149 -44452
rect -3150 -44532 3065 -44468
rect 3129 -44532 3149 -44468
rect -3150 -44548 3149 -44532
rect -3150 -44612 3065 -44548
rect 3129 -44612 3149 -44548
rect -3150 -44628 3149 -44612
rect -3150 -44692 3065 -44628
rect 3129 -44692 3149 -44628
rect -3150 -44708 3149 -44692
rect -3150 -44772 3065 -44708
rect 3129 -44772 3149 -44708
rect -3150 -44788 3149 -44772
rect -3150 -44852 3065 -44788
rect 3129 -44852 3149 -44788
rect -3150 -44868 3149 -44852
rect -3150 -44932 3065 -44868
rect 3129 -44932 3149 -44868
rect -3150 -44948 3149 -44932
rect -3150 -45012 3065 -44948
rect 3129 -45012 3149 -44948
rect -3150 -45028 3149 -45012
rect -3150 -45092 3065 -45028
rect 3129 -45092 3149 -45028
rect -3150 -45108 3149 -45092
rect -3150 -45172 3065 -45108
rect 3129 -45172 3149 -45108
rect -3150 -45188 3149 -45172
rect -3150 -45252 3065 -45188
rect 3129 -45252 3149 -45188
rect -3150 -45268 3149 -45252
rect -3150 -45332 3065 -45268
rect 3129 -45332 3149 -45268
rect -3150 -45348 3149 -45332
rect -3150 -45412 3065 -45348
rect 3129 -45412 3149 -45348
rect -3150 -45428 3149 -45412
rect -3150 -45492 3065 -45428
rect 3129 -45492 3149 -45428
rect -3150 -45508 3149 -45492
rect -3150 -45572 3065 -45508
rect 3129 -45572 3149 -45508
rect -3150 -45588 3149 -45572
rect -3150 -45652 3065 -45588
rect 3129 -45652 3149 -45588
rect -3150 -45668 3149 -45652
rect -3150 -45732 3065 -45668
rect 3129 -45732 3149 -45668
rect -3150 -45748 3149 -45732
rect -3150 -45812 3065 -45748
rect 3129 -45812 3149 -45748
rect -3150 -45828 3149 -45812
rect -3150 -45892 3065 -45828
rect 3129 -45892 3149 -45828
rect -3150 -45908 3149 -45892
rect -3150 -45972 3065 -45908
rect 3129 -45972 3149 -45908
rect -3150 -45988 3149 -45972
rect -3150 -46052 3065 -45988
rect 3129 -46052 3149 -45988
rect -3150 -46068 3149 -46052
rect -3150 -46132 3065 -46068
rect 3129 -46132 3149 -46068
rect -3150 -46148 3149 -46132
rect -3150 -46212 3065 -46148
rect 3129 -46212 3149 -46148
rect -3150 -46228 3149 -46212
rect -3150 -46292 3065 -46228
rect 3129 -46292 3149 -46228
rect -3150 -46308 3149 -46292
rect -3150 -46372 3065 -46308
rect 3129 -46372 3149 -46308
rect -3150 -46388 3149 -46372
rect -3150 -46452 3065 -46388
rect 3129 -46452 3149 -46388
rect -3150 -46468 3149 -46452
rect -3150 -46532 3065 -46468
rect 3129 -46532 3149 -46468
rect -3150 -46548 3149 -46532
rect -3150 -46612 3065 -46548
rect 3129 -46612 3149 -46548
rect -3150 -46628 3149 -46612
rect -3150 -46692 3065 -46628
rect 3129 -46692 3149 -46628
rect -3150 -46708 3149 -46692
rect -3150 -46772 3065 -46708
rect 3129 -46772 3149 -46708
rect -3150 -46788 3149 -46772
rect -3150 -46852 3065 -46788
rect 3129 -46852 3149 -46788
rect -3150 -46868 3149 -46852
rect -3150 -46932 3065 -46868
rect 3129 -46932 3149 -46868
rect -3150 -46948 3149 -46932
rect -3150 -47012 3065 -46948
rect 3129 -47012 3149 -46948
rect -3150 -47028 3149 -47012
rect -3150 -47092 3065 -47028
rect 3129 -47092 3149 -47028
rect -3150 -47108 3149 -47092
rect -3150 -47172 3065 -47108
rect 3129 -47172 3149 -47108
rect -3150 -47200 3149 -47172
rect 3169 -41028 9468 -41000
rect 3169 -41092 9384 -41028
rect 9448 -41092 9468 -41028
rect 3169 -41108 9468 -41092
rect 3169 -41172 9384 -41108
rect 9448 -41172 9468 -41108
rect 3169 -41188 9468 -41172
rect 3169 -41252 9384 -41188
rect 9448 -41252 9468 -41188
rect 3169 -41268 9468 -41252
rect 3169 -41332 9384 -41268
rect 9448 -41332 9468 -41268
rect 3169 -41348 9468 -41332
rect 3169 -41412 9384 -41348
rect 9448 -41412 9468 -41348
rect 3169 -41428 9468 -41412
rect 3169 -41492 9384 -41428
rect 9448 -41492 9468 -41428
rect 3169 -41508 9468 -41492
rect 3169 -41572 9384 -41508
rect 9448 -41572 9468 -41508
rect 3169 -41588 9468 -41572
rect 3169 -41652 9384 -41588
rect 9448 -41652 9468 -41588
rect 3169 -41668 9468 -41652
rect 3169 -41732 9384 -41668
rect 9448 -41732 9468 -41668
rect 3169 -41748 9468 -41732
rect 3169 -41812 9384 -41748
rect 9448 -41812 9468 -41748
rect 3169 -41828 9468 -41812
rect 3169 -41892 9384 -41828
rect 9448 -41892 9468 -41828
rect 3169 -41908 9468 -41892
rect 3169 -41972 9384 -41908
rect 9448 -41972 9468 -41908
rect 3169 -41988 9468 -41972
rect 3169 -42052 9384 -41988
rect 9448 -42052 9468 -41988
rect 3169 -42068 9468 -42052
rect 3169 -42132 9384 -42068
rect 9448 -42132 9468 -42068
rect 3169 -42148 9468 -42132
rect 3169 -42212 9384 -42148
rect 9448 -42212 9468 -42148
rect 3169 -42228 9468 -42212
rect 3169 -42292 9384 -42228
rect 9448 -42292 9468 -42228
rect 3169 -42308 9468 -42292
rect 3169 -42372 9384 -42308
rect 9448 -42372 9468 -42308
rect 3169 -42388 9468 -42372
rect 3169 -42452 9384 -42388
rect 9448 -42452 9468 -42388
rect 3169 -42468 9468 -42452
rect 3169 -42532 9384 -42468
rect 9448 -42532 9468 -42468
rect 3169 -42548 9468 -42532
rect 3169 -42612 9384 -42548
rect 9448 -42612 9468 -42548
rect 3169 -42628 9468 -42612
rect 3169 -42692 9384 -42628
rect 9448 -42692 9468 -42628
rect 3169 -42708 9468 -42692
rect 3169 -42772 9384 -42708
rect 9448 -42772 9468 -42708
rect 3169 -42788 9468 -42772
rect 3169 -42852 9384 -42788
rect 9448 -42852 9468 -42788
rect 3169 -42868 9468 -42852
rect 3169 -42932 9384 -42868
rect 9448 -42932 9468 -42868
rect 3169 -42948 9468 -42932
rect 3169 -43012 9384 -42948
rect 9448 -43012 9468 -42948
rect 3169 -43028 9468 -43012
rect 3169 -43092 9384 -43028
rect 9448 -43092 9468 -43028
rect 3169 -43108 9468 -43092
rect 3169 -43172 9384 -43108
rect 9448 -43172 9468 -43108
rect 3169 -43188 9468 -43172
rect 3169 -43252 9384 -43188
rect 9448 -43252 9468 -43188
rect 3169 -43268 9468 -43252
rect 3169 -43332 9384 -43268
rect 9448 -43332 9468 -43268
rect 3169 -43348 9468 -43332
rect 3169 -43412 9384 -43348
rect 9448 -43412 9468 -43348
rect 3169 -43428 9468 -43412
rect 3169 -43492 9384 -43428
rect 9448 -43492 9468 -43428
rect 3169 -43508 9468 -43492
rect 3169 -43572 9384 -43508
rect 9448 -43572 9468 -43508
rect 3169 -43588 9468 -43572
rect 3169 -43652 9384 -43588
rect 9448 -43652 9468 -43588
rect 3169 -43668 9468 -43652
rect 3169 -43732 9384 -43668
rect 9448 -43732 9468 -43668
rect 3169 -43748 9468 -43732
rect 3169 -43812 9384 -43748
rect 9448 -43812 9468 -43748
rect 3169 -43828 9468 -43812
rect 3169 -43892 9384 -43828
rect 9448 -43892 9468 -43828
rect 3169 -43908 9468 -43892
rect 3169 -43972 9384 -43908
rect 9448 -43972 9468 -43908
rect 3169 -43988 9468 -43972
rect 3169 -44052 9384 -43988
rect 9448 -44052 9468 -43988
rect 3169 -44068 9468 -44052
rect 3169 -44132 9384 -44068
rect 9448 -44132 9468 -44068
rect 3169 -44148 9468 -44132
rect 3169 -44212 9384 -44148
rect 9448 -44212 9468 -44148
rect 3169 -44228 9468 -44212
rect 3169 -44292 9384 -44228
rect 9448 -44292 9468 -44228
rect 3169 -44308 9468 -44292
rect 3169 -44372 9384 -44308
rect 9448 -44372 9468 -44308
rect 3169 -44388 9468 -44372
rect 3169 -44452 9384 -44388
rect 9448 -44452 9468 -44388
rect 3169 -44468 9468 -44452
rect 3169 -44532 9384 -44468
rect 9448 -44532 9468 -44468
rect 3169 -44548 9468 -44532
rect 3169 -44612 9384 -44548
rect 9448 -44612 9468 -44548
rect 3169 -44628 9468 -44612
rect 3169 -44692 9384 -44628
rect 9448 -44692 9468 -44628
rect 3169 -44708 9468 -44692
rect 3169 -44772 9384 -44708
rect 9448 -44772 9468 -44708
rect 3169 -44788 9468 -44772
rect 3169 -44852 9384 -44788
rect 9448 -44852 9468 -44788
rect 3169 -44868 9468 -44852
rect 3169 -44932 9384 -44868
rect 9448 -44932 9468 -44868
rect 3169 -44948 9468 -44932
rect 3169 -45012 9384 -44948
rect 9448 -45012 9468 -44948
rect 3169 -45028 9468 -45012
rect 3169 -45092 9384 -45028
rect 9448 -45092 9468 -45028
rect 3169 -45108 9468 -45092
rect 3169 -45172 9384 -45108
rect 9448 -45172 9468 -45108
rect 3169 -45188 9468 -45172
rect 3169 -45252 9384 -45188
rect 9448 -45252 9468 -45188
rect 3169 -45268 9468 -45252
rect 3169 -45332 9384 -45268
rect 9448 -45332 9468 -45268
rect 3169 -45348 9468 -45332
rect 3169 -45412 9384 -45348
rect 9448 -45412 9468 -45348
rect 3169 -45428 9468 -45412
rect 3169 -45492 9384 -45428
rect 9448 -45492 9468 -45428
rect 3169 -45508 9468 -45492
rect 3169 -45572 9384 -45508
rect 9448 -45572 9468 -45508
rect 3169 -45588 9468 -45572
rect 3169 -45652 9384 -45588
rect 9448 -45652 9468 -45588
rect 3169 -45668 9468 -45652
rect 3169 -45732 9384 -45668
rect 9448 -45732 9468 -45668
rect 3169 -45748 9468 -45732
rect 3169 -45812 9384 -45748
rect 9448 -45812 9468 -45748
rect 3169 -45828 9468 -45812
rect 3169 -45892 9384 -45828
rect 9448 -45892 9468 -45828
rect 3169 -45908 9468 -45892
rect 3169 -45972 9384 -45908
rect 9448 -45972 9468 -45908
rect 3169 -45988 9468 -45972
rect 3169 -46052 9384 -45988
rect 9448 -46052 9468 -45988
rect 3169 -46068 9468 -46052
rect 3169 -46132 9384 -46068
rect 9448 -46132 9468 -46068
rect 3169 -46148 9468 -46132
rect 3169 -46212 9384 -46148
rect 9448 -46212 9468 -46148
rect 3169 -46228 9468 -46212
rect 3169 -46292 9384 -46228
rect 9448 -46292 9468 -46228
rect 3169 -46308 9468 -46292
rect 3169 -46372 9384 -46308
rect 9448 -46372 9468 -46308
rect 3169 -46388 9468 -46372
rect 3169 -46452 9384 -46388
rect 9448 -46452 9468 -46388
rect 3169 -46468 9468 -46452
rect 3169 -46532 9384 -46468
rect 9448 -46532 9468 -46468
rect 3169 -46548 9468 -46532
rect 3169 -46612 9384 -46548
rect 9448 -46612 9468 -46548
rect 3169 -46628 9468 -46612
rect 3169 -46692 9384 -46628
rect 9448 -46692 9468 -46628
rect 3169 -46708 9468 -46692
rect 3169 -46772 9384 -46708
rect 9448 -46772 9468 -46708
rect 3169 -46788 9468 -46772
rect 3169 -46852 9384 -46788
rect 9448 -46852 9468 -46788
rect 3169 -46868 9468 -46852
rect 3169 -46932 9384 -46868
rect 9448 -46932 9468 -46868
rect 3169 -46948 9468 -46932
rect 3169 -47012 9384 -46948
rect 9448 -47012 9468 -46948
rect 3169 -47028 9468 -47012
rect 3169 -47092 9384 -47028
rect 9448 -47092 9468 -47028
rect 3169 -47108 9468 -47092
rect 3169 -47172 9384 -47108
rect 9448 -47172 9468 -47108
rect 3169 -47200 9468 -47172
rect 9488 -41028 15787 -41000
rect 9488 -41092 15703 -41028
rect 15767 -41092 15787 -41028
rect 9488 -41108 15787 -41092
rect 9488 -41172 15703 -41108
rect 15767 -41172 15787 -41108
rect 9488 -41188 15787 -41172
rect 9488 -41252 15703 -41188
rect 15767 -41252 15787 -41188
rect 9488 -41268 15787 -41252
rect 9488 -41332 15703 -41268
rect 15767 -41332 15787 -41268
rect 9488 -41348 15787 -41332
rect 9488 -41412 15703 -41348
rect 15767 -41412 15787 -41348
rect 9488 -41428 15787 -41412
rect 9488 -41492 15703 -41428
rect 15767 -41492 15787 -41428
rect 9488 -41508 15787 -41492
rect 9488 -41572 15703 -41508
rect 15767 -41572 15787 -41508
rect 9488 -41588 15787 -41572
rect 9488 -41652 15703 -41588
rect 15767 -41652 15787 -41588
rect 9488 -41668 15787 -41652
rect 9488 -41732 15703 -41668
rect 15767 -41732 15787 -41668
rect 9488 -41748 15787 -41732
rect 9488 -41812 15703 -41748
rect 15767 -41812 15787 -41748
rect 9488 -41828 15787 -41812
rect 9488 -41892 15703 -41828
rect 15767 -41892 15787 -41828
rect 9488 -41908 15787 -41892
rect 9488 -41972 15703 -41908
rect 15767 -41972 15787 -41908
rect 9488 -41988 15787 -41972
rect 9488 -42052 15703 -41988
rect 15767 -42052 15787 -41988
rect 9488 -42068 15787 -42052
rect 9488 -42132 15703 -42068
rect 15767 -42132 15787 -42068
rect 9488 -42148 15787 -42132
rect 9488 -42212 15703 -42148
rect 15767 -42212 15787 -42148
rect 9488 -42228 15787 -42212
rect 9488 -42292 15703 -42228
rect 15767 -42292 15787 -42228
rect 9488 -42308 15787 -42292
rect 9488 -42372 15703 -42308
rect 15767 -42372 15787 -42308
rect 9488 -42388 15787 -42372
rect 9488 -42452 15703 -42388
rect 15767 -42452 15787 -42388
rect 9488 -42468 15787 -42452
rect 9488 -42532 15703 -42468
rect 15767 -42532 15787 -42468
rect 9488 -42548 15787 -42532
rect 9488 -42612 15703 -42548
rect 15767 -42612 15787 -42548
rect 9488 -42628 15787 -42612
rect 9488 -42692 15703 -42628
rect 15767 -42692 15787 -42628
rect 9488 -42708 15787 -42692
rect 9488 -42772 15703 -42708
rect 15767 -42772 15787 -42708
rect 9488 -42788 15787 -42772
rect 9488 -42852 15703 -42788
rect 15767 -42852 15787 -42788
rect 9488 -42868 15787 -42852
rect 9488 -42932 15703 -42868
rect 15767 -42932 15787 -42868
rect 9488 -42948 15787 -42932
rect 9488 -43012 15703 -42948
rect 15767 -43012 15787 -42948
rect 9488 -43028 15787 -43012
rect 9488 -43092 15703 -43028
rect 15767 -43092 15787 -43028
rect 9488 -43108 15787 -43092
rect 9488 -43172 15703 -43108
rect 15767 -43172 15787 -43108
rect 9488 -43188 15787 -43172
rect 9488 -43252 15703 -43188
rect 15767 -43252 15787 -43188
rect 9488 -43268 15787 -43252
rect 9488 -43332 15703 -43268
rect 15767 -43332 15787 -43268
rect 9488 -43348 15787 -43332
rect 9488 -43412 15703 -43348
rect 15767 -43412 15787 -43348
rect 9488 -43428 15787 -43412
rect 9488 -43492 15703 -43428
rect 15767 -43492 15787 -43428
rect 9488 -43508 15787 -43492
rect 9488 -43572 15703 -43508
rect 15767 -43572 15787 -43508
rect 9488 -43588 15787 -43572
rect 9488 -43652 15703 -43588
rect 15767 -43652 15787 -43588
rect 9488 -43668 15787 -43652
rect 9488 -43732 15703 -43668
rect 15767 -43732 15787 -43668
rect 9488 -43748 15787 -43732
rect 9488 -43812 15703 -43748
rect 15767 -43812 15787 -43748
rect 9488 -43828 15787 -43812
rect 9488 -43892 15703 -43828
rect 15767 -43892 15787 -43828
rect 9488 -43908 15787 -43892
rect 9488 -43972 15703 -43908
rect 15767 -43972 15787 -43908
rect 9488 -43988 15787 -43972
rect 9488 -44052 15703 -43988
rect 15767 -44052 15787 -43988
rect 9488 -44068 15787 -44052
rect 9488 -44132 15703 -44068
rect 15767 -44132 15787 -44068
rect 9488 -44148 15787 -44132
rect 9488 -44212 15703 -44148
rect 15767 -44212 15787 -44148
rect 9488 -44228 15787 -44212
rect 9488 -44292 15703 -44228
rect 15767 -44292 15787 -44228
rect 9488 -44308 15787 -44292
rect 9488 -44372 15703 -44308
rect 15767 -44372 15787 -44308
rect 9488 -44388 15787 -44372
rect 9488 -44452 15703 -44388
rect 15767 -44452 15787 -44388
rect 9488 -44468 15787 -44452
rect 9488 -44532 15703 -44468
rect 15767 -44532 15787 -44468
rect 9488 -44548 15787 -44532
rect 9488 -44612 15703 -44548
rect 15767 -44612 15787 -44548
rect 9488 -44628 15787 -44612
rect 9488 -44692 15703 -44628
rect 15767 -44692 15787 -44628
rect 9488 -44708 15787 -44692
rect 9488 -44772 15703 -44708
rect 15767 -44772 15787 -44708
rect 9488 -44788 15787 -44772
rect 9488 -44852 15703 -44788
rect 15767 -44852 15787 -44788
rect 9488 -44868 15787 -44852
rect 9488 -44932 15703 -44868
rect 15767 -44932 15787 -44868
rect 9488 -44948 15787 -44932
rect 9488 -45012 15703 -44948
rect 15767 -45012 15787 -44948
rect 9488 -45028 15787 -45012
rect 9488 -45092 15703 -45028
rect 15767 -45092 15787 -45028
rect 9488 -45108 15787 -45092
rect 9488 -45172 15703 -45108
rect 15767 -45172 15787 -45108
rect 9488 -45188 15787 -45172
rect 9488 -45252 15703 -45188
rect 15767 -45252 15787 -45188
rect 9488 -45268 15787 -45252
rect 9488 -45332 15703 -45268
rect 15767 -45332 15787 -45268
rect 9488 -45348 15787 -45332
rect 9488 -45412 15703 -45348
rect 15767 -45412 15787 -45348
rect 9488 -45428 15787 -45412
rect 9488 -45492 15703 -45428
rect 15767 -45492 15787 -45428
rect 9488 -45508 15787 -45492
rect 9488 -45572 15703 -45508
rect 15767 -45572 15787 -45508
rect 9488 -45588 15787 -45572
rect 9488 -45652 15703 -45588
rect 15767 -45652 15787 -45588
rect 9488 -45668 15787 -45652
rect 9488 -45732 15703 -45668
rect 15767 -45732 15787 -45668
rect 9488 -45748 15787 -45732
rect 9488 -45812 15703 -45748
rect 15767 -45812 15787 -45748
rect 9488 -45828 15787 -45812
rect 9488 -45892 15703 -45828
rect 15767 -45892 15787 -45828
rect 9488 -45908 15787 -45892
rect 9488 -45972 15703 -45908
rect 15767 -45972 15787 -45908
rect 9488 -45988 15787 -45972
rect 9488 -46052 15703 -45988
rect 15767 -46052 15787 -45988
rect 9488 -46068 15787 -46052
rect 9488 -46132 15703 -46068
rect 15767 -46132 15787 -46068
rect 9488 -46148 15787 -46132
rect 9488 -46212 15703 -46148
rect 15767 -46212 15787 -46148
rect 9488 -46228 15787 -46212
rect 9488 -46292 15703 -46228
rect 15767 -46292 15787 -46228
rect 9488 -46308 15787 -46292
rect 9488 -46372 15703 -46308
rect 15767 -46372 15787 -46308
rect 9488 -46388 15787 -46372
rect 9488 -46452 15703 -46388
rect 15767 -46452 15787 -46388
rect 9488 -46468 15787 -46452
rect 9488 -46532 15703 -46468
rect 15767 -46532 15787 -46468
rect 9488 -46548 15787 -46532
rect 9488 -46612 15703 -46548
rect 15767 -46612 15787 -46548
rect 9488 -46628 15787 -46612
rect 9488 -46692 15703 -46628
rect 15767 -46692 15787 -46628
rect 9488 -46708 15787 -46692
rect 9488 -46772 15703 -46708
rect 15767 -46772 15787 -46708
rect 9488 -46788 15787 -46772
rect 9488 -46852 15703 -46788
rect 15767 -46852 15787 -46788
rect 9488 -46868 15787 -46852
rect 9488 -46932 15703 -46868
rect 15767 -46932 15787 -46868
rect 9488 -46948 15787 -46932
rect 9488 -47012 15703 -46948
rect 15767 -47012 15787 -46948
rect 9488 -47028 15787 -47012
rect 9488 -47092 15703 -47028
rect 15767 -47092 15787 -47028
rect 9488 -47108 15787 -47092
rect 9488 -47172 15703 -47108
rect 15767 -47172 15787 -47108
rect 9488 -47200 15787 -47172
rect 15807 -41028 22106 -41000
rect 15807 -41092 22022 -41028
rect 22086 -41092 22106 -41028
rect 15807 -41108 22106 -41092
rect 15807 -41172 22022 -41108
rect 22086 -41172 22106 -41108
rect 15807 -41188 22106 -41172
rect 15807 -41252 22022 -41188
rect 22086 -41252 22106 -41188
rect 15807 -41268 22106 -41252
rect 15807 -41332 22022 -41268
rect 22086 -41332 22106 -41268
rect 15807 -41348 22106 -41332
rect 15807 -41412 22022 -41348
rect 22086 -41412 22106 -41348
rect 15807 -41428 22106 -41412
rect 15807 -41492 22022 -41428
rect 22086 -41492 22106 -41428
rect 15807 -41508 22106 -41492
rect 15807 -41572 22022 -41508
rect 22086 -41572 22106 -41508
rect 15807 -41588 22106 -41572
rect 15807 -41652 22022 -41588
rect 22086 -41652 22106 -41588
rect 15807 -41668 22106 -41652
rect 15807 -41732 22022 -41668
rect 22086 -41732 22106 -41668
rect 15807 -41748 22106 -41732
rect 15807 -41812 22022 -41748
rect 22086 -41812 22106 -41748
rect 15807 -41828 22106 -41812
rect 15807 -41892 22022 -41828
rect 22086 -41892 22106 -41828
rect 15807 -41908 22106 -41892
rect 15807 -41972 22022 -41908
rect 22086 -41972 22106 -41908
rect 15807 -41988 22106 -41972
rect 15807 -42052 22022 -41988
rect 22086 -42052 22106 -41988
rect 15807 -42068 22106 -42052
rect 15807 -42132 22022 -42068
rect 22086 -42132 22106 -42068
rect 15807 -42148 22106 -42132
rect 15807 -42212 22022 -42148
rect 22086 -42212 22106 -42148
rect 15807 -42228 22106 -42212
rect 15807 -42292 22022 -42228
rect 22086 -42292 22106 -42228
rect 15807 -42308 22106 -42292
rect 15807 -42372 22022 -42308
rect 22086 -42372 22106 -42308
rect 15807 -42388 22106 -42372
rect 15807 -42452 22022 -42388
rect 22086 -42452 22106 -42388
rect 15807 -42468 22106 -42452
rect 15807 -42532 22022 -42468
rect 22086 -42532 22106 -42468
rect 15807 -42548 22106 -42532
rect 15807 -42612 22022 -42548
rect 22086 -42612 22106 -42548
rect 15807 -42628 22106 -42612
rect 15807 -42692 22022 -42628
rect 22086 -42692 22106 -42628
rect 15807 -42708 22106 -42692
rect 15807 -42772 22022 -42708
rect 22086 -42772 22106 -42708
rect 15807 -42788 22106 -42772
rect 15807 -42852 22022 -42788
rect 22086 -42852 22106 -42788
rect 15807 -42868 22106 -42852
rect 15807 -42932 22022 -42868
rect 22086 -42932 22106 -42868
rect 15807 -42948 22106 -42932
rect 15807 -43012 22022 -42948
rect 22086 -43012 22106 -42948
rect 15807 -43028 22106 -43012
rect 15807 -43092 22022 -43028
rect 22086 -43092 22106 -43028
rect 15807 -43108 22106 -43092
rect 15807 -43172 22022 -43108
rect 22086 -43172 22106 -43108
rect 15807 -43188 22106 -43172
rect 15807 -43252 22022 -43188
rect 22086 -43252 22106 -43188
rect 15807 -43268 22106 -43252
rect 15807 -43332 22022 -43268
rect 22086 -43332 22106 -43268
rect 15807 -43348 22106 -43332
rect 15807 -43412 22022 -43348
rect 22086 -43412 22106 -43348
rect 15807 -43428 22106 -43412
rect 15807 -43492 22022 -43428
rect 22086 -43492 22106 -43428
rect 15807 -43508 22106 -43492
rect 15807 -43572 22022 -43508
rect 22086 -43572 22106 -43508
rect 15807 -43588 22106 -43572
rect 15807 -43652 22022 -43588
rect 22086 -43652 22106 -43588
rect 15807 -43668 22106 -43652
rect 15807 -43732 22022 -43668
rect 22086 -43732 22106 -43668
rect 15807 -43748 22106 -43732
rect 15807 -43812 22022 -43748
rect 22086 -43812 22106 -43748
rect 15807 -43828 22106 -43812
rect 15807 -43892 22022 -43828
rect 22086 -43892 22106 -43828
rect 15807 -43908 22106 -43892
rect 15807 -43972 22022 -43908
rect 22086 -43972 22106 -43908
rect 15807 -43988 22106 -43972
rect 15807 -44052 22022 -43988
rect 22086 -44052 22106 -43988
rect 15807 -44068 22106 -44052
rect 15807 -44132 22022 -44068
rect 22086 -44132 22106 -44068
rect 15807 -44148 22106 -44132
rect 15807 -44212 22022 -44148
rect 22086 -44212 22106 -44148
rect 15807 -44228 22106 -44212
rect 15807 -44292 22022 -44228
rect 22086 -44292 22106 -44228
rect 15807 -44308 22106 -44292
rect 15807 -44372 22022 -44308
rect 22086 -44372 22106 -44308
rect 15807 -44388 22106 -44372
rect 15807 -44452 22022 -44388
rect 22086 -44452 22106 -44388
rect 15807 -44468 22106 -44452
rect 15807 -44532 22022 -44468
rect 22086 -44532 22106 -44468
rect 15807 -44548 22106 -44532
rect 15807 -44612 22022 -44548
rect 22086 -44612 22106 -44548
rect 15807 -44628 22106 -44612
rect 15807 -44692 22022 -44628
rect 22086 -44692 22106 -44628
rect 15807 -44708 22106 -44692
rect 15807 -44772 22022 -44708
rect 22086 -44772 22106 -44708
rect 15807 -44788 22106 -44772
rect 15807 -44852 22022 -44788
rect 22086 -44852 22106 -44788
rect 15807 -44868 22106 -44852
rect 15807 -44932 22022 -44868
rect 22086 -44932 22106 -44868
rect 15807 -44948 22106 -44932
rect 15807 -45012 22022 -44948
rect 22086 -45012 22106 -44948
rect 15807 -45028 22106 -45012
rect 15807 -45092 22022 -45028
rect 22086 -45092 22106 -45028
rect 15807 -45108 22106 -45092
rect 15807 -45172 22022 -45108
rect 22086 -45172 22106 -45108
rect 15807 -45188 22106 -45172
rect 15807 -45252 22022 -45188
rect 22086 -45252 22106 -45188
rect 15807 -45268 22106 -45252
rect 15807 -45332 22022 -45268
rect 22086 -45332 22106 -45268
rect 15807 -45348 22106 -45332
rect 15807 -45412 22022 -45348
rect 22086 -45412 22106 -45348
rect 15807 -45428 22106 -45412
rect 15807 -45492 22022 -45428
rect 22086 -45492 22106 -45428
rect 15807 -45508 22106 -45492
rect 15807 -45572 22022 -45508
rect 22086 -45572 22106 -45508
rect 15807 -45588 22106 -45572
rect 15807 -45652 22022 -45588
rect 22086 -45652 22106 -45588
rect 15807 -45668 22106 -45652
rect 15807 -45732 22022 -45668
rect 22086 -45732 22106 -45668
rect 15807 -45748 22106 -45732
rect 15807 -45812 22022 -45748
rect 22086 -45812 22106 -45748
rect 15807 -45828 22106 -45812
rect 15807 -45892 22022 -45828
rect 22086 -45892 22106 -45828
rect 15807 -45908 22106 -45892
rect 15807 -45972 22022 -45908
rect 22086 -45972 22106 -45908
rect 15807 -45988 22106 -45972
rect 15807 -46052 22022 -45988
rect 22086 -46052 22106 -45988
rect 15807 -46068 22106 -46052
rect 15807 -46132 22022 -46068
rect 22086 -46132 22106 -46068
rect 15807 -46148 22106 -46132
rect 15807 -46212 22022 -46148
rect 22086 -46212 22106 -46148
rect 15807 -46228 22106 -46212
rect 15807 -46292 22022 -46228
rect 22086 -46292 22106 -46228
rect 15807 -46308 22106 -46292
rect 15807 -46372 22022 -46308
rect 22086 -46372 22106 -46308
rect 15807 -46388 22106 -46372
rect 15807 -46452 22022 -46388
rect 22086 -46452 22106 -46388
rect 15807 -46468 22106 -46452
rect 15807 -46532 22022 -46468
rect 22086 -46532 22106 -46468
rect 15807 -46548 22106 -46532
rect 15807 -46612 22022 -46548
rect 22086 -46612 22106 -46548
rect 15807 -46628 22106 -46612
rect 15807 -46692 22022 -46628
rect 22086 -46692 22106 -46628
rect 15807 -46708 22106 -46692
rect 15807 -46772 22022 -46708
rect 22086 -46772 22106 -46708
rect 15807 -46788 22106 -46772
rect 15807 -46852 22022 -46788
rect 22086 -46852 22106 -46788
rect 15807 -46868 22106 -46852
rect 15807 -46932 22022 -46868
rect 22086 -46932 22106 -46868
rect 15807 -46948 22106 -46932
rect 15807 -47012 22022 -46948
rect 22086 -47012 22106 -46948
rect 15807 -47028 22106 -47012
rect 15807 -47092 22022 -47028
rect 22086 -47092 22106 -47028
rect 15807 -47108 22106 -47092
rect 15807 -47172 22022 -47108
rect 22086 -47172 22106 -47108
rect 15807 -47200 22106 -47172
rect 22126 -41028 28425 -41000
rect 22126 -41092 28341 -41028
rect 28405 -41092 28425 -41028
rect 22126 -41108 28425 -41092
rect 22126 -41172 28341 -41108
rect 28405 -41172 28425 -41108
rect 22126 -41188 28425 -41172
rect 22126 -41252 28341 -41188
rect 28405 -41252 28425 -41188
rect 22126 -41268 28425 -41252
rect 22126 -41332 28341 -41268
rect 28405 -41332 28425 -41268
rect 22126 -41348 28425 -41332
rect 22126 -41412 28341 -41348
rect 28405 -41412 28425 -41348
rect 22126 -41428 28425 -41412
rect 22126 -41492 28341 -41428
rect 28405 -41492 28425 -41428
rect 22126 -41508 28425 -41492
rect 22126 -41572 28341 -41508
rect 28405 -41572 28425 -41508
rect 22126 -41588 28425 -41572
rect 22126 -41652 28341 -41588
rect 28405 -41652 28425 -41588
rect 22126 -41668 28425 -41652
rect 22126 -41732 28341 -41668
rect 28405 -41732 28425 -41668
rect 22126 -41748 28425 -41732
rect 22126 -41812 28341 -41748
rect 28405 -41812 28425 -41748
rect 22126 -41828 28425 -41812
rect 22126 -41892 28341 -41828
rect 28405 -41892 28425 -41828
rect 22126 -41908 28425 -41892
rect 22126 -41972 28341 -41908
rect 28405 -41972 28425 -41908
rect 22126 -41988 28425 -41972
rect 22126 -42052 28341 -41988
rect 28405 -42052 28425 -41988
rect 22126 -42068 28425 -42052
rect 22126 -42132 28341 -42068
rect 28405 -42132 28425 -42068
rect 22126 -42148 28425 -42132
rect 22126 -42212 28341 -42148
rect 28405 -42212 28425 -42148
rect 22126 -42228 28425 -42212
rect 22126 -42292 28341 -42228
rect 28405 -42292 28425 -42228
rect 22126 -42308 28425 -42292
rect 22126 -42372 28341 -42308
rect 28405 -42372 28425 -42308
rect 22126 -42388 28425 -42372
rect 22126 -42452 28341 -42388
rect 28405 -42452 28425 -42388
rect 22126 -42468 28425 -42452
rect 22126 -42532 28341 -42468
rect 28405 -42532 28425 -42468
rect 22126 -42548 28425 -42532
rect 22126 -42612 28341 -42548
rect 28405 -42612 28425 -42548
rect 22126 -42628 28425 -42612
rect 22126 -42692 28341 -42628
rect 28405 -42692 28425 -42628
rect 22126 -42708 28425 -42692
rect 22126 -42772 28341 -42708
rect 28405 -42772 28425 -42708
rect 22126 -42788 28425 -42772
rect 22126 -42852 28341 -42788
rect 28405 -42852 28425 -42788
rect 22126 -42868 28425 -42852
rect 22126 -42932 28341 -42868
rect 28405 -42932 28425 -42868
rect 22126 -42948 28425 -42932
rect 22126 -43012 28341 -42948
rect 28405 -43012 28425 -42948
rect 22126 -43028 28425 -43012
rect 22126 -43092 28341 -43028
rect 28405 -43092 28425 -43028
rect 22126 -43108 28425 -43092
rect 22126 -43172 28341 -43108
rect 28405 -43172 28425 -43108
rect 22126 -43188 28425 -43172
rect 22126 -43252 28341 -43188
rect 28405 -43252 28425 -43188
rect 22126 -43268 28425 -43252
rect 22126 -43332 28341 -43268
rect 28405 -43332 28425 -43268
rect 22126 -43348 28425 -43332
rect 22126 -43412 28341 -43348
rect 28405 -43412 28425 -43348
rect 22126 -43428 28425 -43412
rect 22126 -43492 28341 -43428
rect 28405 -43492 28425 -43428
rect 22126 -43508 28425 -43492
rect 22126 -43572 28341 -43508
rect 28405 -43572 28425 -43508
rect 22126 -43588 28425 -43572
rect 22126 -43652 28341 -43588
rect 28405 -43652 28425 -43588
rect 22126 -43668 28425 -43652
rect 22126 -43732 28341 -43668
rect 28405 -43732 28425 -43668
rect 22126 -43748 28425 -43732
rect 22126 -43812 28341 -43748
rect 28405 -43812 28425 -43748
rect 22126 -43828 28425 -43812
rect 22126 -43892 28341 -43828
rect 28405 -43892 28425 -43828
rect 22126 -43908 28425 -43892
rect 22126 -43972 28341 -43908
rect 28405 -43972 28425 -43908
rect 22126 -43988 28425 -43972
rect 22126 -44052 28341 -43988
rect 28405 -44052 28425 -43988
rect 22126 -44068 28425 -44052
rect 22126 -44132 28341 -44068
rect 28405 -44132 28425 -44068
rect 22126 -44148 28425 -44132
rect 22126 -44212 28341 -44148
rect 28405 -44212 28425 -44148
rect 22126 -44228 28425 -44212
rect 22126 -44292 28341 -44228
rect 28405 -44292 28425 -44228
rect 22126 -44308 28425 -44292
rect 22126 -44372 28341 -44308
rect 28405 -44372 28425 -44308
rect 22126 -44388 28425 -44372
rect 22126 -44452 28341 -44388
rect 28405 -44452 28425 -44388
rect 22126 -44468 28425 -44452
rect 22126 -44532 28341 -44468
rect 28405 -44532 28425 -44468
rect 22126 -44548 28425 -44532
rect 22126 -44612 28341 -44548
rect 28405 -44612 28425 -44548
rect 22126 -44628 28425 -44612
rect 22126 -44692 28341 -44628
rect 28405 -44692 28425 -44628
rect 22126 -44708 28425 -44692
rect 22126 -44772 28341 -44708
rect 28405 -44772 28425 -44708
rect 22126 -44788 28425 -44772
rect 22126 -44852 28341 -44788
rect 28405 -44852 28425 -44788
rect 22126 -44868 28425 -44852
rect 22126 -44932 28341 -44868
rect 28405 -44932 28425 -44868
rect 22126 -44948 28425 -44932
rect 22126 -45012 28341 -44948
rect 28405 -45012 28425 -44948
rect 22126 -45028 28425 -45012
rect 22126 -45092 28341 -45028
rect 28405 -45092 28425 -45028
rect 22126 -45108 28425 -45092
rect 22126 -45172 28341 -45108
rect 28405 -45172 28425 -45108
rect 22126 -45188 28425 -45172
rect 22126 -45252 28341 -45188
rect 28405 -45252 28425 -45188
rect 22126 -45268 28425 -45252
rect 22126 -45332 28341 -45268
rect 28405 -45332 28425 -45268
rect 22126 -45348 28425 -45332
rect 22126 -45412 28341 -45348
rect 28405 -45412 28425 -45348
rect 22126 -45428 28425 -45412
rect 22126 -45492 28341 -45428
rect 28405 -45492 28425 -45428
rect 22126 -45508 28425 -45492
rect 22126 -45572 28341 -45508
rect 28405 -45572 28425 -45508
rect 22126 -45588 28425 -45572
rect 22126 -45652 28341 -45588
rect 28405 -45652 28425 -45588
rect 22126 -45668 28425 -45652
rect 22126 -45732 28341 -45668
rect 28405 -45732 28425 -45668
rect 22126 -45748 28425 -45732
rect 22126 -45812 28341 -45748
rect 28405 -45812 28425 -45748
rect 22126 -45828 28425 -45812
rect 22126 -45892 28341 -45828
rect 28405 -45892 28425 -45828
rect 22126 -45908 28425 -45892
rect 22126 -45972 28341 -45908
rect 28405 -45972 28425 -45908
rect 22126 -45988 28425 -45972
rect 22126 -46052 28341 -45988
rect 28405 -46052 28425 -45988
rect 22126 -46068 28425 -46052
rect 22126 -46132 28341 -46068
rect 28405 -46132 28425 -46068
rect 22126 -46148 28425 -46132
rect 22126 -46212 28341 -46148
rect 28405 -46212 28425 -46148
rect 22126 -46228 28425 -46212
rect 22126 -46292 28341 -46228
rect 28405 -46292 28425 -46228
rect 22126 -46308 28425 -46292
rect 22126 -46372 28341 -46308
rect 28405 -46372 28425 -46308
rect 22126 -46388 28425 -46372
rect 22126 -46452 28341 -46388
rect 28405 -46452 28425 -46388
rect 22126 -46468 28425 -46452
rect 22126 -46532 28341 -46468
rect 28405 -46532 28425 -46468
rect 22126 -46548 28425 -46532
rect 22126 -46612 28341 -46548
rect 28405 -46612 28425 -46548
rect 22126 -46628 28425 -46612
rect 22126 -46692 28341 -46628
rect 28405 -46692 28425 -46628
rect 22126 -46708 28425 -46692
rect 22126 -46772 28341 -46708
rect 28405 -46772 28425 -46708
rect 22126 -46788 28425 -46772
rect 22126 -46852 28341 -46788
rect 28405 -46852 28425 -46788
rect 22126 -46868 28425 -46852
rect 22126 -46932 28341 -46868
rect 28405 -46932 28425 -46868
rect 22126 -46948 28425 -46932
rect 22126 -47012 28341 -46948
rect 28405 -47012 28425 -46948
rect 22126 -47028 28425 -47012
rect 22126 -47092 28341 -47028
rect 28405 -47092 28425 -47028
rect 22126 -47108 28425 -47092
rect 22126 -47172 28341 -47108
rect 28405 -47172 28425 -47108
rect 22126 -47200 28425 -47172
rect 28445 -41028 34744 -41000
rect 28445 -41092 34660 -41028
rect 34724 -41092 34744 -41028
rect 28445 -41108 34744 -41092
rect 28445 -41172 34660 -41108
rect 34724 -41172 34744 -41108
rect 28445 -41188 34744 -41172
rect 28445 -41252 34660 -41188
rect 34724 -41252 34744 -41188
rect 28445 -41268 34744 -41252
rect 28445 -41332 34660 -41268
rect 34724 -41332 34744 -41268
rect 28445 -41348 34744 -41332
rect 28445 -41412 34660 -41348
rect 34724 -41412 34744 -41348
rect 28445 -41428 34744 -41412
rect 28445 -41492 34660 -41428
rect 34724 -41492 34744 -41428
rect 28445 -41508 34744 -41492
rect 28445 -41572 34660 -41508
rect 34724 -41572 34744 -41508
rect 28445 -41588 34744 -41572
rect 28445 -41652 34660 -41588
rect 34724 -41652 34744 -41588
rect 28445 -41668 34744 -41652
rect 28445 -41732 34660 -41668
rect 34724 -41732 34744 -41668
rect 28445 -41748 34744 -41732
rect 28445 -41812 34660 -41748
rect 34724 -41812 34744 -41748
rect 28445 -41828 34744 -41812
rect 28445 -41892 34660 -41828
rect 34724 -41892 34744 -41828
rect 28445 -41908 34744 -41892
rect 28445 -41972 34660 -41908
rect 34724 -41972 34744 -41908
rect 28445 -41988 34744 -41972
rect 28445 -42052 34660 -41988
rect 34724 -42052 34744 -41988
rect 28445 -42068 34744 -42052
rect 28445 -42132 34660 -42068
rect 34724 -42132 34744 -42068
rect 28445 -42148 34744 -42132
rect 28445 -42212 34660 -42148
rect 34724 -42212 34744 -42148
rect 28445 -42228 34744 -42212
rect 28445 -42292 34660 -42228
rect 34724 -42292 34744 -42228
rect 28445 -42308 34744 -42292
rect 28445 -42372 34660 -42308
rect 34724 -42372 34744 -42308
rect 28445 -42388 34744 -42372
rect 28445 -42452 34660 -42388
rect 34724 -42452 34744 -42388
rect 28445 -42468 34744 -42452
rect 28445 -42532 34660 -42468
rect 34724 -42532 34744 -42468
rect 28445 -42548 34744 -42532
rect 28445 -42612 34660 -42548
rect 34724 -42612 34744 -42548
rect 28445 -42628 34744 -42612
rect 28445 -42692 34660 -42628
rect 34724 -42692 34744 -42628
rect 28445 -42708 34744 -42692
rect 28445 -42772 34660 -42708
rect 34724 -42772 34744 -42708
rect 28445 -42788 34744 -42772
rect 28445 -42852 34660 -42788
rect 34724 -42852 34744 -42788
rect 28445 -42868 34744 -42852
rect 28445 -42932 34660 -42868
rect 34724 -42932 34744 -42868
rect 28445 -42948 34744 -42932
rect 28445 -43012 34660 -42948
rect 34724 -43012 34744 -42948
rect 28445 -43028 34744 -43012
rect 28445 -43092 34660 -43028
rect 34724 -43092 34744 -43028
rect 28445 -43108 34744 -43092
rect 28445 -43172 34660 -43108
rect 34724 -43172 34744 -43108
rect 28445 -43188 34744 -43172
rect 28445 -43252 34660 -43188
rect 34724 -43252 34744 -43188
rect 28445 -43268 34744 -43252
rect 28445 -43332 34660 -43268
rect 34724 -43332 34744 -43268
rect 28445 -43348 34744 -43332
rect 28445 -43412 34660 -43348
rect 34724 -43412 34744 -43348
rect 28445 -43428 34744 -43412
rect 28445 -43492 34660 -43428
rect 34724 -43492 34744 -43428
rect 28445 -43508 34744 -43492
rect 28445 -43572 34660 -43508
rect 34724 -43572 34744 -43508
rect 28445 -43588 34744 -43572
rect 28445 -43652 34660 -43588
rect 34724 -43652 34744 -43588
rect 28445 -43668 34744 -43652
rect 28445 -43732 34660 -43668
rect 34724 -43732 34744 -43668
rect 28445 -43748 34744 -43732
rect 28445 -43812 34660 -43748
rect 34724 -43812 34744 -43748
rect 28445 -43828 34744 -43812
rect 28445 -43892 34660 -43828
rect 34724 -43892 34744 -43828
rect 28445 -43908 34744 -43892
rect 28445 -43972 34660 -43908
rect 34724 -43972 34744 -43908
rect 28445 -43988 34744 -43972
rect 28445 -44052 34660 -43988
rect 34724 -44052 34744 -43988
rect 28445 -44068 34744 -44052
rect 28445 -44132 34660 -44068
rect 34724 -44132 34744 -44068
rect 28445 -44148 34744 -44132
rect 28445 -44212 34660 -44148
rect 34724 -44212 34744 -44148
rect 28445 -44228 34744 -44212
rect 28445 -44292 34660 -44228
rect 34724 -44292 34744 -44228
rect 28445 -44308 34744 -44292
rect 28445 -44372 34660 -44308
rect 34724 -44372 34744 -44308
rect 28445 -44388 34744 -44372
rect 28445 -44452 34660 -44388
rect 34724 -44452 34744 -44388
rect 28445 -44468 34744 -44452
rect 28445 -44532 34660 -44468
rect 34724 -44532 34744 -44468
rect 28445 -44548 34744 -44532
rect 28445 -44612 34660 -44548
rect 34724 -44612 34744 -44548
rect 28445 -44628 34744 -44612
rect 28445 -44692 34660 -44628
rect 34724 -44692 34744 -44628
rect 28445 -44708 34744 -44692
rect 28445 -44772 34660 -44708
rect 34724 -44772 34744 -44708
rect 28445 -44788 34744 -44772
rect 28445 -44852 34660 -44788
rect 34724 -44852 34744 -44788
rect 28445 -44868 34744 -44852
rect 28445 -44932 34660 -44868
rect 34724 -44932 34744 -44868
rect 28445 -44948 34744 -44932
rect 28445 -45012 34660 -44948
rect 34724 -45012 34744 -44948
rect 28445 -45028 34744 -45012
rect 28445 -45092 34660 -45028
rect 34724 -45092 34744 -45028
rect 28445 -45108 34744 -45092
rect 28445 -45172 34660 -45108
rect 34724 -45172 34744 -45108
rect 28445 -45188 34744 -45172
rect 28445 -45252 34660 -45188
rect 34724 -45252 34744 -45188
rect 28445 -45268 34744 -45252
rect 28445 -45332 34660 -45268
rect 34724 -45332 34744 -45268
rect 28445 -45348 34744 -45332
rect 28445 -45412 34660 -45348
rect 34724 -45412 34744 -45348
rect 28445 -45428 34744 -45412
rect 28445 -45492 34660 -45428
rect 34724 -45492 34744 -45428
rect 28445 -45508 34744 -45492
rect 28445 -45572 34660 -45508
rect 34724 -45572 34744 -45508
rect 28445 -45588 34744 -45572
rect 28445 -45652 34660 -45588
rect 34724 -45652 34744 -45588
rect 28445 -45668 34744 -45652
rect 28445 -45732 34660 -45668
rect 34724 -45732 34744 -45668
rect 28445 -45748 34744 -45732
rect 28445 -45812 34660 -45748
rect 34724 -45812 34744 -45748
rect 28445 -45828 34744 -45812
rect 28445 -45892 34660 -45828
rect 34724 -45892 34744 -45828
rect 28445 -45908 34744 -45892
rect 28445 -45972 34660 -45908
rect 34724 -45972 34744 -45908
rect 28445 -45988 34744 -45972
rect 28445 -46052 34660 -45988
rect 34724 -46052 34744 -45988
rect 28445 -46068 34744 -46052
rect 28445 -46132 34660 -46068
rect 34724 -46132 34744 -46068
rect 28445 -46148 34744 -46132
rect 28445 -46212 34660 -46148
rect 34724 -46212 34744 -46148
rect 28445 -46228 34744 -46212
rect 28445 -46292 34660 -46228
rect 34724 -46292 34744 -46228
rect 28445 -46308 34744 -46292
rect 28445 -46372 34660 -46308
rect 34724 -46372 34744 -46308
rect 28445 -46388 34744 -46372
rect 28445 -46452 34660 -46388
rect 34724 -46452 34744 -46388
rect 28445 -46468 34744 -46452
rect 28445 -46532 34660 -46468
rect 34724 -46532 34744 -46468
rect 28445 -46548 34744 -46532
rect 28445 -46612 34660 -46548
rect 34724 -46612 34744 -46548
rect 28445 -46628 34744 -46612
rect 28445 -46692 34660 -46628
rect 34724 -46692 34744 -46628
rect 28445 -46708 34744 -46692
rect 28445 -46772 34660 -46708
rect 34724 -46772 34744 -46708
rect 28445 -46788 34744 -46772
rect 28445 -46852 34660 -46788
rect 34724 -46852 34744 -46788
rect 28445 -46868 34744 -46852
rect 28445 -46932 34660 -46868
rect 34724 -46932 34744 -46868
rect 28445 -46948 34744 -46932
rect 28445 -47012 34660 -46948
rect 34724 -47012 34744 -46948
rect 28445 -47028 34744 -47012
rect 28445 -47092 34660 -47028
rect 34724 -47092 34744 -47028
rect 28445 -47108 34744 -47092
rect 28445 -47172 34660 -47108
rect 34724 -47172 34744 -47108
rect 28445 -47200 34744 -47172
rect 34764 -41028 41063 -41000
rect 34764 -41092 40979 -41028
rect 41043 -41092 41063 -41028
rect 34764 -41108 41063 -41092
rect 34764 -41172 40979 -41108
rect 41043 -41172 41063 -41108
rect 34764 -41188 41063 -41172
rect 34764 -41252 40979 -41188
rect 41043 -41252 41063 -41188
rect 34764 -41268 41063 -41252
rect 34764 -41332 40979 -41268
rect 41043 -41332 41063 -41268
rect 34764 -41348 41063 -41332
rect 34764 -41412 40979 -41348
rect 41043 -41412 41063 -41348
rect 34764 -41428 41063 -41412
rect 34764 -41492 40979 -41428
rect 41043 -41492 41063 -41428
rect 34764 -41508 41063 -41492
rect 34764 -41572 40979 -41508
rect 41043 -41572 41063 -41508
rect 34764 -41588 41063 -41572
rect 34764 -41652 40979 -41588
rect 41043 -41652 41063 -41588
rect 34764 -41668 41063 -41652
rect 34764 -41732 40979 -41668
rect 41043 -41732 41063 -41668
rect 34764 -41748 41063 -41732
rect 34764 -41812 40979 -41748
rect 41043 -41812 41063 -41748
rect 34764 -41828 41063 -41812
rect 34764 -41892 40979 -41828
rect 41043 -41892 41063 -41828
rect 34764 -41908 41063 -41892
rect 34764 -41972 40979 -41908
rect 41043 -41972 41063 -41908
rect 34764 -41988 41063 -41972
rect 34764 -42052 40979 -41988
rect 41043 -42052 41063 -41988
rect 34764 -42068 41063 -42052
rect 34764 -42132 40979 -42068
rect 41043 -42132 41063 -42068
rect 34764 -42148 41063 -42132
rect 34764 -42212 40979 -42148
rect 41043 -42212 41063 -42148
rect 34764 -42228 41063 -42212
rect 34764 -42292 40979 -42228
rect 41043 -42292 41063 -42228
rect 34764 -42308 41063 -42292
rect 34764 -42372 40979 -42308
rect 41043 -42372 41063 -42308
rect 34764 -42388 41063 -42372
rect 34764 -42452 40979 -42388
rect 41043 -42452 41063 -42388
rect 34764 -42468 41063 -42452
rect 34764 -42532 40979 -42468
rect 41043 -42532 41063 -42468
rect 34764 -42548 41063 -42532
rect 34764 -42612 40979 -42548
rect 41043 -42612 41063 -42548
rect 34764 -42628 41063 -42612
rect 34764 -42692 40979 -42628
rect 41043 -42692 41063 -42628
rect 34764 -42708 41063 -42692
rect 34764 -42772 40979 -42708
rect 41043 -42772 41063 -42708
rect 34764 -42788 41063 -42772
rect 34764 -42852 40979 -42788
rect 41043 -42852 41063 -42788
rect 34764 -42868 41063 -42852
rect 34764 -42932 40979 -42868
rect 41043 -42932 41063 -42868
rect 34764 -42948 41063 -42932
rect 34764 -43012 40979 -42948
rect 41043 -43012 41063 -42948
rect 34764 -43028 41063 -43012
rect 34764 -43092 40979 -43028
rect 41043 -43092 41063 -43028
rect 34764 -43108 41063 -43092
rect 34764 -43172 40979 -43108
rect 41043 -43172 41063 -43108
rect 34764 -43188 41063 -43172
rect 34764 -43252 40979 -43188
rect 41043 -43252 41063 -43188
rect 34764 -43268 41063 -43252
rect 34764 -43332 40979 -43268
rect 41043 -43332 41063 -43268
rect 34764 -43348 41063 -43332
rect 34764 -43412 40979 -43348
rect 41043 -43412 41063 -43348
rect 34764 -43428 41063 -43412
rect 34764 -43492 40979 -43428
rect 41043 -43492 41063 -43428
rect 34764 -43508 41063 -43492
rect 34764 -43572 40979 -43508
rect 41043 -43572 41063 -43508
rect 34764 -43588 41063 -43572
rect 34764 -43652 40979 -43588
rect 41043 -43652 41063 -43588
rect 34764 -43668 41063 -43652
rect 34764 -43732 40979 -43668
rect 41043 -43732 41063 -43668
rect 34764 -43748 41063 -43732
rect 34764 -43812 40979 -43748
rect 41043 -43812 41063 -43748
rect 34764 -43828 41063 -43812
rect 34764 -43892 40979 -43828
rect 41043 -43892 41063 -43828
rect 34764 -43908 41063 -43892
rect 34764 -43972 40979 -43908
rect 41043 -43972 41063 -43908
rect 34764 -43988 41063 -43972
rect 34764 -44052 40979 -43988
rect 41043 -44052 41063 -43988
rect 34764 -44068 41063 -44052
rect 34764 -44132 40979 -44068
rect 41043 -44132 41063 -44068
rect 34764 -44148 41063 -44132
rect 34764 -44212 40979 -44148
rect 41043 -44212 41063 -44148
rect 34764 -44228 41063 -44212
rect 34764 -44292 40979 -44228
rect 41043 -44292 41063 -44228
rect 34764 -44308 41063 -44292
rect 34764 -44372 40979 -44308
rect 41043 -44372 41063 -44308
rect 34764 -44388 41063 -44372
rect 34764 -44452 40979 -44388
rect 41043 -44452 41063 -44388
rect 34764 -44468 41063 -44452
rect 34764 -44532 40979 -44468
rect 41043 -44532 41063 -44468
rect 34764 -44548 41063 -44532
rect 34764 -44612 40979 -44548
rect 41043 -44612 41063 -44548
rect 34764 -44628 41063 -44612
rect 34764 -44692 40979 -44628
rect 41043 -44692 41063 -44628
rect 34764 -44708 41063 -44692
rect 34764 -44772 40979 -44708
rect 41043 -44772 41063 -44708
rect 34764 -44788 41063 -44772
rect 34764 -44852 40979 -44788
rect 41043 -44852 41063 -44788
rect 34764 -44868 41063 -44852
rect 34764 -44932 40979 -44868
rect 41043 -44932 41063 -44868
rect 34764 -44948 41063 -44932
rect 34764 -45012 40979 -44948
rect 41043 -45012 41063 -44948
rect 34764 -45028 41063 -45012
rect 34764 -45092 40979 -45028
rect 41043 -45092 41063 -45028
rect 34764 -45108 41063 -45092
rect 34764 -45172 40979 -45108
rect 41043 -45172 41063 -45108
rect 34764 -45188 41063 -45172
rect 34764 -45252 40979 -45188
rect 41043 -45252 41063 -45188
rect 34764 -45268 41063 -45252
rect 34764 -45332 40979 -45268
rect 41043 -45332 41063 -45268
rect 34764 -45348 41063 -45332
rect 34764 -45412 40979 -45348
rect 41043 -45412 41063 -45348
rect 34764 -45428 41063 -45412
rect 34764 -45492 40979 -45428
rect 41043 -45492 41063 -45428
rect 34764 -45508 41063 -45492
rect 34764 -45572 40979 -45508
rect 41043 -45572 41063 -45508
rect 34764 -45588 41063 -45572
rect 34764 -45652 40979 -45588
rect 41043 -45652 41063 -45588
rect 34764 -45668 41063 -45652
rect 34764 -45732 40979 -45668
rect 41043 -45732 41063 -45668
rect 34764 -45748 41063 -45732
rect 34764 -45812 40979 -45748
rect 41043 -45812 41063 -45748
rect 34764 -45828 41063 -45812
rect 34764 -45892 40979 -45828
rect 41043 -45892 41063 -45828
rect 34764 -45908 41063 -45892
rect 34764 -45972 40979 -45908
rect 41043 -45972 41063 -45908
rect 34764 -45988 41063 -45972
rect 34764 -46052 40979 -45988
rect 41043 -46052 41063 -45988
rect 34764 -46068 41063 -46052
rect 34764 -46132 40979 -46068
rect 41043 -46132 41063 -46068
rect 34764 -46148 41063 -46132
rect 34764 -46212 40979 -46148
rect 41043 -46212 41063 -46148
rect 34764 -46228 41063 -46212
rect 34764 -46292 40979 -46228
rect 41043 -46292 41063 -46228
rect 34764 -46308 41063 -46292
rect 34764 -46372 40979 -46308
rect 41043 -46372 41063 -46308
rect 34764 -46388 41063 -46372
rect 34764 -46452 40979 -46388
rect 41043 -46452 41063 -46388
rect 34764 -46468 41063 -46452
rect 34764 -46532 40979 -46468
rect 41043 -46532 41063 -46468
rect 34764 -46548 41063 -46532
rect 34764 -46612 40979 -46548
rect 41043 -46612 41063 -46548
rect 34764 -46628 41063 -46612
rect 34764 -46692 40979 -46628
rect 41043 -46692 41063 -46628
rect 34764 -46708 41063 -46692
rect 34764 -46772 40979 -46708
rect 41043 -46772 41063 -46708
rect 34764 -46788 41063 -46772
rect 34764 -46852 40979 -46788
rect 41043 -46852 41063 -46788
rect 34764 -46868 41063 -46852
rect 34764 -46932 40979 -46868
rect 41043 -46932 41063 -46868
rect 34764 -46948 41063 -46932
rect 34764 -47012 40979 -46948
rect 41043 -47012 41063 -46948
rect 34764 -47028 41063 -47012
rect 34764 -47092 40979 -47028
rect 41043 -47092 41063 -47028
rect 34764 -47108 41063 -47092
rect 34764 -47172 40979 -47108
rect 41043 -47172 41063 -47108
rect 34764 -47200 41063 -47172
rect 41083 -41028 47382 -41000
rect 41083 -41092 47298 -41028
rect 47362 -41092 47382 -41028
rect 41083 -41108 47382 -41092
rect 41083 -41172 47298 -41108
rect 47362 -41172 47382 -41108
rect 41083 -41188 47382 -41172
rect 41083 -41252 47298 -41188
rect 47362 -41252 47382 -41188
rect 41083 -41268 47382 -41252
rect 41083 -41332 47298 -41268
rect 47362 -41332 47382 -41268
rect 41083 -41348 47382 -41332
rect 41083 -41412 47298 -41348
rect 47362 -41412 47382 -41348
rect 41083 -41428 47382 -41412
rect 41083 -41492 47298 -41428
rect 47362 -41492 47382 -41428
rect 41083 -41508 47382 -41492
rect 41083 -41572 47298 -41508
rect 47362 -41572 47382 -41508
rect 41083 -41588 47382 -41572
rect 41083 -41652 47298 -41588
rect 47362 -41652 47382 -41588
rect 41083 -41668 47382 -41652
rect 41083 -41732 47298 -41668
rect 47362 -41732 47382 -41668
rect 41083 -41748 47382 -41732
rect 41083 -41812 47298 -41748
rect 47362 -41812 47382 -41748
rect 41083 -41828 47382 -41812
rect 41083 -41892 47298 -41828
rect 47362 -41892 47382 -41828
rect 41083 -41908 47382 -41892
rect 41083 -41972 47298 -41908
rect 47362 -41972 47382 -41908
rect 41083 -41988 47382 -41972
rect 41083 -42052 47298 -41988
rect 47362 -42052 47382 -41988
rect 41083 -42068 47382 -42052
rect 41083 -42132 47298 -42068
rect 47362 -42132 47382 -42068
rect 41083 -42148 47382 -42132
rect 41083 -42212 47298 -42148
rect 47362 -42212 47382 -42148
rect 41083 -42228 47382 -42212
rect 41083 -42292 47298 -42228
rect 47362 -42292 47382 -42228
rect 41083 -42308 47382 -42292
rect 41083 -42372 47298 -42308
rect 47362 -42372 47382 -42308
rect 41083 -42388 47382 -42372
rect 41083 -42452 47298 -42388
rect 47362 -42452 47382 -42388
rect 41083 -42468 47382 -42452
rect 41083 -42532 47298 -42468
rect 47362 -42532 47382 -42468
rect 41083 -42548 47382 -42532
rect 41083 -42612 47298 -42548
rect 47362 -42612 47382 -42548
rect 41083 -42628 47382 -42612
rect 41083 -42692 47298 -42628
rect 47362 -42692 47382 -42628
rect 41083 -42708 47382 -42692
rect 41083 -42772 47298 -42708
rect 47362 -42772 47382 -42708
rect 41083 -42788 47382 -42772
rect 41083 -42852 47298 -42788
rect 47362 -42852 47382 -42788
rect 41083 -42868 47382 -42852
rect 41083 -42932 47298 -42868
rect 47362 -42932 47382 -42868
rect 41083 -42948 47382 -42932
rect 41083 -43012 47298 -42948
rect 47362 -43012 47382 -42948
rect 41083 -43028 47382 -43012
rect 41083 -43092 47298 -43028
rect 47362 -43092 47382 -43028
rect 41083 -43108 47382 -43092
rect 41083 -43172 47298 -43108
rect 47362 -43172 47382 -43108
rect 41083 -43188 47382 -43172
rect 41083 -43252 47298 -43188
rect 47362 -43252 47382 -43188
rect 41083 -43268 47382 -43252
rect 41083 -43332 47298 -43268
rect 47362 -43332 47382 -43268
rect 41083 -43348 47382 -43332
rect 41083 -43412 47298 -43348
rect 47362 -43412 47382 -43348
rect 41083 -43428 47382 -43412
rect 41083 -43492 47298 -43428
rect 47362 -43492 47382 -43428
rect 41083 -43508 47382 -43492
rect 41083 -43572 47298 -43508
rect 47362 -43572 47382 -43508
rect 41083 -43588 47382 -43572
rect 41083 -43652 47298 -43588
rect 47362 -43652 47382 -43588
rect 41083 -43668 47382 -43652
rect 41083 -43732 47298 -43668
rect 47362 -43732 47382 -43668
rect 41083 -43748 47382 -43732
rect 41083 -43812 47298 -43748
rect 47362 -43812 47382 -43748
rect 41083 -43828 47382 -43812
rect 41083 -43892 47298 -43828
rect 47362 -43892 47382 -43828
rect 41083 -43908 47382 -43892
rect 41083 -43972 47298 -43908
rect 47362 -43972 47382 -43908
rect 41083 -43988 47382 -43972
rect 41083 -44052 47298 -43988
rect 47362 -44052 47382 -43988
rect 41083 -44068 47382 -44052
rect 41083 -44132 47298 -44068
rect 47362 -44132 47382 -44068
rect 41083 -44148 47382 -44132
rect 41083 -44212 47298 -44148
rect 47362 -44212 47382 -44148
rect 41083 -44228 47382 -44212
rect 41083 -44292 47298 -44228
rect 47362 -44292 47382 -44228
rect 41083 -44308 47382 -44292
rect 41083 -44372 47298 -44308
rect 47362 -44372 47382 -44308
rect 41083 -44388 47382 -44372
rect 41083 -44452 47298 -44388
rect 47362 -44452 47382 -44388
rect 41083 -44468 47382 -44452
rect 41083 -44532 47298 -44468
rect 47362 -44532 47382 -44468
rect 41083 -44548 47382 -44532
rect 41083 -44612 47298 -44548
rect 47362 -44612 47382 -44548
rect 41083 -44628 47382 -44612
rect 41083 -44692 47298 -44628
rect 47362 -44692 47382 -44628
rect 41083 -44708 47382 -44692
rect 41083 -44772 47298 -44708
rect 47362 -44772 47382 -44708
rect 41083 -44788 47382 -44772
rect 41083 -44852 47298 -44788
rect 47362 -44852 47382 -44788
rect 41083 -44868 47382 -44852
rect 41083 -44932 47298 -44868
rect 47362 -44932 47382 -44868
rect 41083 -44948 47382 -44932
rect 41083 -45012 47298 -44948
rect 47362 -45012 47382 -44948
rect 41083 -45028 47382 -45012
rect 41083 -45092 47298 -45028
rect 47362 -45092 47382 -45028
rect 41083 -45108 47382 -45092
rect 41083 -45172 47298 -45108
rect 47362 -45172 47382 -45108
rect 41083 -45188 47382 -45172
rect 41083 -45252 47298 -45188
rect 47362 -45252 47382 -45188
rect 41083 -45268 47382 -45252
rect 41083 -45332 47298 -45268
rect 47362 -45332 47382 -45268
rect 41083 -45348 47382 -45332
rect 41083 -45412 47298 -45348
rect 47362 -45412 47382 -45348
rect 41083 -45428 47382 -45412
rect 41083 -45492 47298 -45428
rect 47362 -45492 47382 -45428
rect 41083 -45508 47382 -45492
rect 41083 -45572 47298 -45508
rect 47362 -45572 47382 -45508
rect 41083 -45588 47382 -45572
rect 41083 -45652 47298 -45588
rect 47362 -45652 47382 -45588
rect 41083 -45668 47382 -45652
rect 41083 -45732 47298 -45668
rect 47362 -45732 47382 -45668
rect 41083 -45748 47382 -45732
rect 41083 -45812 47298 -45748
rect 47362 -45812 47382 -45748
rect 41083 -45828 47382 -45812
rect 41083 -45892 47298 -45828
rect 47362 -45892 47382 -45828
rect 41083 -45908 47382 -45892
rect 41083 -45972 47298 -45908
rect 47362 -45972 47382 -45908
rect 41083 -45988 47382 -45972
rect 41083 -46052 47298 -45988
rect 47362 -46052 47382 -45988
rect 41083 -46068 47382 -46052
rect 41083 -46132 47298 -46068
rect 47362 -46132 47382 -46068
rect 41083 -46148 47382 -46132
rect 41083 -46212 47298 -46148
rect 47362 -46212 47382 -46148
rect 41083 -46228 47382 -46212
rect 41083 -46292 47298 -46228
rect 47362 -46292 47382 -46228
rect 41083 -46308 47382 -46292
rect 41083 -46372 47298 -46308
rect 47362 -46372 47382 -46308
rect 41083 -46388 47382 -46372
rect 41083 -46452 47298 -46388
rect 47362 -46452 47382 -46388
rect 41083 -46468 47382 -46452
rect 41083 -46532 47298 -46468
rect 47362 -46532 47382 -46468
rect 41083 -46548 47382 -46532
rect 41083 -46612 47298 -46548
rect 47362 -46612 47382 -46548
rect 41083 -46628 47382 -46612
rect 41083 -46692 47298 -46628
rect 47362 -46692 47382 -46628
rect 41083 -46708 47382 -46692
rect 41083 -46772 47298 -46708
rect 47362 -46772 47382 -46708
rect 41083 -46788 47382 -46772
rect 41083 -46852 47298 -46788
rect 47362 -46852 47382 -46788
rect 41083 -46868 47382 -46852
rect 41083 -46932 47298 -46868
rect 47362 -46932 47382 -46868
rect 41083 -46948 47382 -46932
rect 41083 -47012 47298 -46948
rect 47362 -47012 47382 -46948
rect 41083 -47028 47382 -47012
rect 41083 -47092 47298 -47028
rect 47362 -47092 47382 -47028
rect 41083 -47108 47382 -47092
rect 41083 -47172 47298 -47108
rect 47362 -47172 47382 -47108
rect 41083 -47200 47382 -47172
<< via3 >>
rect -41168 47108 -41104 47172
rect -41168 47028 -41104 47092
rect -41168 46948 -41104 47012
rect -41168 46868 -41104 46932
rect -41168 46788 -41104 46852
rect -41168 46708 -41104 46772
rect -41168 46628 -41104 46692
rect -41168 46548 -41104 46612
rect -41168 46468 -41104 46532
rect -41168 46388 -41104 46452
rect -41168 46308 -41104 46372
rect -41168 46228 -41104 46292
rect -41168 46148 -41104 46212
rect -41168 46068 -41104 46132
rect -41168 45988 -41104 46052
rect -41168 45908 -41104 45972
rect -41168 45828 -41104 45892
rect -41168 45748 -41104 45812
rect -41168 45668 -41104 45732
rect -41168 45588 -41104 45652
rect -41168 45508 -41104 45572
rect -41168 45428 -41104 45492
rect -41168 45348 -41104 45412
rect -41168 45268 -41104 45332
rect -41168 45188 -41104 45252
rect -41168 45108 -41104 45172
rect -41168 45028 -41104 45092
rect -41168 44948 -41104 45012
rect -41168 44868 -41104 44932
rect -41168 44788 -41104 44852
rect -41168 44708 -41104 44772
rect -41168 44628 -41104 44692
rect -41168 44548 -41104 44612
rect -41168 44468 -41104 44532
rect -41168 44388 -41104 44452
rect -41168 44308 -41104 44372
rect -41168 44228 -41104 44292
rect -41168 44148 -41104 44212
rect -41168 44068 -41104 44132
rect -41168 43988 -41104 44052
rect -41168 43908 -41104 43972
rect -41168 43828 -41104 43892
rect -41168 43748 -41104 43812
rect -41168 43668 -41104 43732
rect -41168 43588 -41104 43652
rect -41168 43508 -41104 43572
rect -41168 43428 -41104 43492
rect -41168 43348 -41104 43412
rect -41168 43268 -41104 43332
rect -41168 43188 -41104 43252
rect -41168 43108 -41104 43172
rect -41168 43028 -41104 43092
rect -41168 42948 -41104 43012
rect -41168 42868 -41104 42932
rect -41168 42788 -41104 42852
rect -41168 42708 -41104 42772
rect -41168 42628 -41104 42692
rect -41168 42548 -41104 42612
rect -41168 42468 -41104 42532
rect -41168 42388 -41104 42452
rect -41168 42308 -41104 42372
rect -41168 42228 -41104 42292
rect -41168 42148 -41104 42212
rect -41168 42068 -41104 42132
rect -41168 41988 -41104 42052
rect -41168 41908 -41104 41972
rect -41168 41828 -41104 41892
rect -41168 41748 -41104 41812
rect -41168 41668 -41104 41732
rect -41168 41588 -41104 41652
rect -41168 41508 -41104 41572
rect -41168 41428 -41104 41492
rect -41168 41348 -41104 41412
rect -41168 41268 -41104 41332
rect -41168 41188 -41104 41252
rect -41168 41108 -41104 41172
rect -41168 41028 -41104 41092
rect -34849 47108 -34785 47172
rect -34849 47028 -34785 47092
rect -34849 46948 -34785 47012
rect -34849 46868 -34785 46932
rect -34849 46788 -34785 46852
rect -34849 46708 -34785 46772
rect -34849 46628 -34785 46692
rect -34849 46548 -34785 46612
rect -34849 46468 -34785 46532
rect -34849 46388 -34785 46452
rect -34849 46308 -34785 46372
rect -34849 46228 -34785 46292
rect -34849 46148 -34785 46212
rect -34849 46068 -34785 46132
rect -34849 45988 -34785 46052
rect -34849 45908 -34785 45972
rect -34849 45828 -34785 45892
rect -34849 45748 -34785 45812
rect -34849 45668 -34785 45732
rect -34849 45588 -34785 45652
rect -34849 45508 -34785 45572
rect -34849 45428 -34785 45492
rect -34849 45348 -34785 45412
rect -34849 45268 -34785 45332
rect -34849 45188 -34785 45252
rect -34849 45108 -34785 45172
rect -34849 45028 -34785 45092
rect -34849 44948 -34785 45012
rect -34849 44868 -34785 44932
rect -34849 44788 -34785 44852
rect -34849 44708 -34785 44772
rect -34849 44628 -34785 44692
rect -34849 44548 -34785 44612
rect -34849 44468 -34785 44532
rect -34849 44388 -34785 44452
rect -34849 44308 -34785 44372
rect -34849 44228 -34785 44292
rect -34849 44148 -34785 44212
rect -34849 44068 -34785 44132
rect -34849 43988 -34785 44052
rect -34849 43908 -34785 43972
rect -34849 43828 -34785 43892
rect -34849 43748 -34785 43812
rect -34849 43668 -34785 43732
rect -34849 43588 -34785 43652
rect -34849 43508 -34785 43572
rect -34849 43428 -34785 43492
rect -34849 43348 -34785 43412
rect -34849 43268 -34785 43332
rect -34849 43188 -34785 43252
rect -34849 43108 -34785 43172
rect -34849 43028 -34785 43092
rect -34849 42948 -34785 43012
rect -34849 42868 -34785 42932
rect -34849 42788 -34785 42852
rect -34849 42708 -34785 42772
rect -34849 42628 -34785 42692
rect -34849 42548 -34785 42612
rect -34849 42468 -34785 42532
rect -34849 42388 -34785 42452
rect -34849 42308 -34785 42372
rect -34849 42228 -34785 42292
rect -34849 42148 -34785 42212
rect -34849 42068 -34785 42132
rect -34849 41988 -34785 42052
rect -34849 41908 -34785 41972
rect -34849 41828 -34785 41892
rect -34849 41748 -34785 41812
rect -34849 41668 -34785 41732
rect -34849 41588 -34785 41652
rect -34849 41508 -34785 41572
rect -34849 41428 -34785 41492
rect -34849 41348 -34785 41412
rect -34849 41268 -34785 41332
rect -34849 41188 -34785 41252
rect -34849 41108 -34785 41172
rect -34849 41028 -34785 41092
rect -28530 47108 -28466 47172
rect -28530 47028 -28466 47092
rect -28530 46948 -28466 47012
rect -28530 46868 -28466 46932
rect -28530 46788 -28466 46852
rect -28530 46708 -28466 46772
rect -28530 46628 -28466 46692
rect -28530 46548 -28466 46612
rect -28530 46468 -28466 46532
rect -28530 46388 -28466 46452
rect -28530 46308 -28466 46372
rect -28530 46228 -28466 46292
rect -28530 46148 -28466 46212
rect -28530 46068 -28466 46132
rect -28530 45988 -28466 46052
rect -28530 45908 -28466 45972
rect -28530 45828 -28466 45892
rect -28530 45748 -28466 45812
rect -28530 45668 -28466 45732
rect -28530 45588 -28466 45652
rect -28530 45508 -28466 45572
rect -28530 45428 -28466 45492
rect -28530 45348 -28466 45412
rect -28530 45268 -28466 45332
rect -28530 45188 -28466 45252
rect -28530 45108 -28466 45172
rect -28530 45028 -28466 45092
rect -28530 44948 -28466 45012
rect -28530 44868 -28466 44932
rect -28530 44788 -28466 44852
rect -28530 44708 -28466 44772
rect -28530 44628 -28466 44692
rect -28530 44548 -28466 44612
rect -28530 44468 -28466 44532
rect -28530 44388 -28466 44452
rect -28530 44308 -28466 44372
rect -28530 44228 -28466 44292
rect -28530 44148 -28466 44212
rect -28530 44068 -28466 44132
rect -28530 43988 -28466 44052
rect -28530 43908 -28466 43972
rect -28530 43828 -28466 43892
rect -28530 43748 -28466 43812
rect -28530 43668 -28466 43732
rect -28530 43588 -28466 43652
rect -28530 43508 -28466 43572
rect -28530 43428 -28466 43492
rect -28530 43348 -28466 43412
rect -28530 43268 -28466 43332
rect -28530 43188 -28466 43252
rect -28530 43108 -28466 43172
rect -28530 43028 -28466 43092
rect -28530 42948 -28466 43012
rect -28530 42868 -28466 42932
rect -28530 42788 -28466 42852
rect -28530 42708 -28466 42772
rect -28530 42628 -28466 42692
rect -28530 42548 -28466 42612
rect -28530 42468 -28466 42532
rect -28530 42388 -28466 42452
rect -28530 42308 -28466 42372
rect -28530 42228 -28466 42292
rect -28530 42148 -28466 42212
rect -28530 42068 -28466 42132
rect -28530 41988 -28466 42052
rect -28530 41908 -28466 41972
rect -28530 41828 -28466 41892
rect -28530 41748 -28466 41812
rect -28530 41668 -28466 41732
rect -28530 41588 -28466 41652
rect -28530 41508 -28466 41572
rect -28530 41428 -28466 41492
rect -28530 41348 -28466 41412
rect -28530 41268 -28466 41332
rect -28530 41188 -28466 41252
rect -28530 41108 -28466 41172
rect -28530 41028 -28466 41092
rect -22211 47108 -22147 47172
rect -22211 47028 -22147 47092
rect -22211 46948 -22147 47012
rect -22211 46868 -22147 46932
rect -22211 46788 -22147 46852
rect -22211 46708 -22147 46772
rect -22211 46628 -22147 46692
rect -22211 46548 -22147 46612
rect -22211 46468 -22147 46532
rect -22211 46388 -22147 46452
rect -22211 46308 -22147 46372
rect -22211 46228 -22147 46292
rect -22211 46148 -22147 46212
rect -22211 46068 -22147 46132
rect -22211 45988 -22147 46052
rect -22211 45908 -22147 45972
rect -22211 45828 -22147 45892
rect -22211 45748 -22147 45812
rect -22211 45668 -22147 45732
rect -22211 45588 -22147 45652
rect -22211 45508 -22147 45572
rect -22211 45428 -22147 45492
rect -22211 45348 -22147 45412
rect -22211 45268 -22147 45332
rect -22211 45188 -22147 45252
rect -22211 45108 -22147 45172
rect -22211 45028 -22147 45092
rect -22211 44948 -22147 45012
rect -22211 44868 -22147 44932
rect -22211 44788 -22147 44852
rect -22211 44708 -22147 44772
rect -22211 44628 -22147 44692
rect -22211 44548 -22147 44612
rect -22211 44468 -22147 44532
rect -22211 44388 -22147 44452
rect -22211 44308 -22147 44372
rect -22211 44228 -22147 44292
rect -22211 44148 -22147 44212
rect -22211 44068 -22147 44132
rect -22211 43988 -22147 44052
rect -22211 43908 -22147 43972
rect -22211 43828 -22147 43892
rect -22211 43748 -22147 43812
rect -22211 43668 -22147 43732
rect -22211 43588 -22147 43652
rect -22211 43508 -22147 43572
rect -22211 43428 -22147 43492
rect -22211 43348 -22147 43412
rect -22211 43268 -22147 43332
rect -22211 43188 -22147 43252
rect -22211 43108 -22147 43172
rect -22211 43028 -22147 43092
rect -22211 42948 -22147 43012
rect -22211 42868 -22147 42932
rect -22211 42788 -22147 42852
rect -22211 42708 -22147 42772
rect -22211 42628 -22147 42692
rect -22211 42548 -22147 42612
rect -22211 42468 -22147 42532
rect -22211 42388 -22147 42452
rect -22211 42308 -22147 42372
rect -22211 42228 -22147 42292
rect -22211 42148 -22147 42212
rect -22211 42068 -22147 42132
rect -22211 41988 -22147 42052
rect -22211 41908 -22147 41972
rect -22211 41828 -22147 41892
rect -22211 41748 -22147 41812
rect -22211 41668 -22147 41732
rect -22211 41588 -22147 41652
rect -22211 41508 -22147 41572
rect -22211 41428 -22147 41492
rect -22211 41348 -22147 41412
rect -22211 41268 -22147 41332
rect -22211 41188 -22147 41252
rect -22211 41108 -22147 41172
rect -22211 41028 -22147 41092
rect -15892 47108 -15828 47172
rect -15892 47028 -15828 47092
rect -15892 46948 -15828 47012
rect -15892 46868 -15828 46932
rect -15892 46788 -15828 46852
rect -15892 46708 -15828 46772
rect -15892 46628 -15828 46692
rect -15892 46548 -15828 46612
rect -15892 46468 -15828 46532
rect -15892 46388 -15828 46452
rect -15892 46308 -15828 46372
rect -15892 46228 -15828 46292
rect -15892 46148 -15828 46212
rect -15892 46068 -15828 46132
rect -15892 45988 -15828 46052
rect -15892 45908 -15828 45972
rect -15892 45828 -15828 45892
rect -15892 45748 -15828 45812
rect -15892 45668 -15828 45732
rect -15892 45588 -15828 45652
rect -15892 45508 -15828 45572
rect -15892 45428 -15828 45492
rect -15892 45348 -15828 45412
rect -15892 45268 -15828 45332
rect -15892 45188 -15828 45252
rect -15892 45108 -15828 45172
rect -15892 45028 -15828 45092
rect -15892 44948 -15828 45012
rect -15892 44868 -15828 44932
rect -15892 44788 -15828 44852
rect -15892 44708 -15828 44772
rect -15892 44628 -15828 44692
rect -15892 44548 -15828 44612
rect -15892 44468 -15828 44532
rect -15892 44388 -15828 44452
rect -15892 44308 -15828 44372
rect -15892 44228 -15828 44292
rect -15892 44148 -15828 44212
rect -15892 44068 -15828 44132
rect -15892 43988 -15828 44052
rect -15892 43908 -15828 43972
rect -15892 43828 -15828 43892
rect -15892 43748 -15828 43812
rect -15892 43668 -15828 43732
rect -15892 43588 -15828 43652
rect -15892 43508 -15828 43572
rect -15892 43428 -15828 43492
rect -15892 43348 -15828 43412
rect -15892 43268 -15828 43332
rect -15892 43188 -15828 43252
rect -15892 43108 -15828 43172
rect -15892 43028 -15828 43092
rect -15892 42948 -15828 43012
rect -15892 42868 -15828 42932
rect -15892 42788 -15828 42852
rect -15892 42708 -15828 42772
rect -15892 42628 -15828 42692
rect -15892 42548 -15828 42612
rect -15892 42468 -15828 42532
rect -15892 42388 -15828 42452
rect -15892 42308 -15828 42372
rect -15892 42228 -15828 42292
rect -15892 42148 -15828 42212
rect -15892 42068 -15828 42132
rect -15892 41988 -15828 42052
rect -15892 41908 -15828 41972
rect -15892 41828 -15828 41892
rect -15892 41748 -15828 41812
rect -15892 41668 -15828 41732
rect -15892 41588 -15828 41652
rect -15892 41508 -15828 41572
rect -15892 41428 -15828 41492
rect -15892 41348 -15828 41412
rect -15892 41268 -15828 41332
rect -15892 41188 -15828 41252
rect -15892 41108 -15828 41172
rect -15892 41028 -15828 41092
rect -9573 47108 -9509 47172
rect -9573 47028 -9509 47092
rect -9573 46948 -9509 47012
rect -9573 46868 -9509 46932
rect -9573 46788 -9509 46852
rect -9573 46708 -9509 46772
rect -9573 46628 -9509 46692
rect -9573 46548 -9509 46612
rect -9573 46468 -9509 46532
rect -9573 46388 -9509 46452
rect -9573 46308 -9509 46372
rect -9573 46228 -9509 46292
rect -9573 46148 -9509 46212
rect -9573 46068 -9509 46132
rect -9573 45988 -9509 46052
rect -9573 45908 -9509 45972
rect -9573 45828 -9509 45892
rect -9573 45748 -9509 45812
rect -9573 45668 -9509 45732
rect -9573 45588 -9509 45652
rect -9573 45508 -9509 45572
rect -9573 45428 -9509 45492
rect -9573 45348 -9509 45412
rect -9573 45268 -9509 45332
rect -9573 45188 -9509 45252
rect -9573 45108 -9509 45172
rect -9573 45028 -9509 45092
rect -9573 44948 -9509 45012
rect -9573 44868 -9509 44932
rect -9573 44788 -9509 44852
rect -9573 44708 -9509 44772
rect -9573 44628 -9509 44692
rect -9573 44548 -9509 44612
rect -9573 44468 -9509 44532
rect -9573 44388 -9509 44452
rect -9573 44308 -9509 44372
rect -9573 44228 -9509 44292
rect -9573 44148 -9509 44212
rect -9573 44068 -9509 44132
rect -9573 43988 -9509 44052
rect -9573 43908 -9509 43972
rect -9573 43828 -9509 43892
rect -9573 43748 -9509 43812
rect -9573 43668 -9509 43732
rect -9573 43588 -9509 43652
rect -9573 43508 -9509 43572
rect -9573 43428 -9509 43492
rect -9573 43348 -9509 43412
rect -9573 43268 -9509 43332
rect -9573 43188 -9509 43252
rect -9573 43108 -9509 43172
rect -9573 43028 -9509 43092
rect -9573 42948 -9509 43012
rect -9573 42868 -9509 42932
rect -9573 42788 -9509 42852
rect -9573 42708 -9509 42772
rect -9573 42628 -9509 42692
rect -9573 42548 -9509 42612
rect -9573 42468 -9509 42532
rect -9573 42388 -9509 42452
rect -9573 42308 -9509 42372
rect -9573 42228 -9509 42292
rect -9573 42148 -9509 42212
rect -9573 42068 -9509 42132
rect -9573 41988 -9509 42052
rect -9573 41908 -9509 41972
rect -9573 41828 -9509 41892
rect -9573 41748 -9509 41812
rect -9573 41668 -9509 41732
rect -9573 41588 -9509 41652
rect -9573 41508 -9509 41572
rect -9573 41428 -9509 41492
rect -9573 41348 -9509 41412
rect -9573 41268 -9509 41332
rect -9573 41188 -9509 41252
rect -9573 41108 -9509 41172
rect -9573 41028 -9509 41092
rect -3254 47108 -3190 47172
rect -3254 47028 -3190 47092
rect -3254 46948 -3190 47012
rect -3254 46868 -3190 46932
rect -3254 46788 -3190 46852
rect -3254 46708 -3190 46772
rect -3254 46628 -3190 46692
rect -3254 46548 -3190 46612
rect -3254 46468 -3190 46532
rect -3254 46388 -3190 46452
rect -3254 46308 -3190 46372
rect -3254 46228 -3190 46292
rect -3254 46148 -3190 46212
rect -3254 46068 -3190 46132
rect -3254 45988 -3190 46052
rect -3254 45908 -3190 45972
rect -3254 45828 -3190 45892
rect -3254 45748 -3190 45812
rect -3254 45668 -3190 45732
rect -3254 45588 -3190 45652
rect -3254 45508 -3190 45572
rect -3254 45428 -3190 45492
rect -3254 45348 -3190 45412
rect -3254 45268 -3190 45332
rect -3254 45188 -3190 45252
rect -3254 45108 -3190 45172
rect -3254 45028 -3190 45092
rect -3254 44948 -3190 45012
rect -3254 44868 -3190 44932
rect -3254 44788 -3190 44852
rect -3254 44708 -3190 44772
rect -3254 44628 -3190 44692
rect -3254 44548 -3190 44612
rect -3254 44468 -3190 44532
rect -3254 44388 -3190 44452
rect -3254 44308 -3190 44372
rect -3254 44228 -3190 44292
rect -3254 44148 -3190 44212
rect -3254 44068 -3190 44132
rect -3254 43988 -3190 44052
rect -3254 43908 -3190 43972
rect -3254 43828 -3190 43892
rect -3254 43748 -3190 43812
rect -3254 43668 -3190 43732
rect -3254 43588 -3190 43652
rect -3254 43508 -3190 43572
rect -3254 43428 -3190 43492
rect -3254 43348 -3190 43412
rect -3254 43268 -3190 43332
rect -3254 43188 -3190 43252
rect -3254 43108 -3190 43172
rect -3254 43028 -3190 43092
rect -3254 42948 -3190 43012
rect -3254 42868 -3190 42932
rect -3254 42788 -3190 42852
rect -3254 42708 -3190 42772
rect -3254 42628 -3190 42692
rect -3254 42548 -3190 42612
rect -3254 42468 -3190 42532
rect -3254 42388 -3190 42452
rect -3254 42308 -3190 42372
rect -3254 42228 -3190 42292
rect -3254 42148 -3190 42212
rect -3254 42068 -3190 42132
rect -3254 41988 -3190 42052
rect -3254 41908 -3190 41972
rect -3254 41828 -3190 41892
rect -3254 41748 -3190 41812
rect -3254 41668 -3190 41732
rect -3254 41588 -3190 41652
rect -3254 41508 -3190 41572
rect -3254 41428 -3190 41492
rect -3254 41348 -3190 41412
rect -3254 41268 -3190 41332
rect -3254 41188 -3190 41252
rect -3254 41108 -3190 41172
rect -3254 41028 -3190 41092
rect 3065 47108 3129 47172
rect 3065 47028 3129 47092
rect 3065 46948 3129 47012
rect 3065 46868 3129 46932
rect 3065 46788 3129 46852
rect 3065 46708 3129 46772
rect 3065 46628 3129 46692
rect 3065 46548 3129 46612
rect 3065 46468 3129 46532
rect 3065 46388 3129 46452
rect 3065 46308 3129 46372
rect 3065 46228 3129 46292
rect 3065 46148 3129 46212
rect 3065 46068 3129 46132
rect 3065 45988 3129 46052
rect 3065 45908 3129 45972
rect 3065 45828 3129 45892
rect 3065 45748 3129 45812
rect 3065 45668 3129 45732
rect 3065 45588 3129 45652
rect 3065 45508 3129 45572
rect 3065 45428 3129 45492
rect 3065 45348 3129 45412
rect 3065 45268 3129 45332
rect 3065 45188 3129 45252
rect 3065 45108 3129 45172
rect 3065 45028 3129 45092
rect 3065 44948 3129 45012
rect 3065 44868 3129 44932
rect 3065 44788 3129 44852
rect 3065 44708 3129 44772
rect 3065 44628 3129 44692
rect 3065 44548 3129 44612
rect 3065 44468 3129 44532
rect 3065 44388 3129 44452
rect 3065 44308 3129 44372
rect 3065 44228 3129 44292
rect 3065 44148 3129 44212
rect 3065 44068 3129 44132
rect 3065 43988 3129 44052
rect 3065 43908 3129 43972
rect 3065 43828 3129 43892
rect 3065 43748 3129 43812
rect 3065 43668 3129 43732
rect 3065 43588 3129 43652
rect 3065 43508 3129 43572
rect 3065 43428 3129 43492
rect 3065 43348 3129 43412
rect 3065 43268 3129 43332
rect 3065 43188 3129 43252
rect 3065 43108 3129 43172
rect 3065 43028 3129 43092
rect 3065 42948 3129 43012
rect 3065 42868 3129 42932
rect 3065 42788 3129 42852
rect 3065 42708 3129 42772
rect 3065 42628 3129 42692
rect 3065 42548 3129 42612
rect 3065 42468 3129 42532
rect 3065 42388 3129 42452
rect 3065 42308 3129 42372
rect 3065 42228 3129 42292
rect 3065 42148 3129 42212
rect 3065 42068 3129 42132
rect 3065 41988 3129 42052
rect 3065 41908 3129 41972
rect 3065 41828 3129 41892
rect 3065 41748 3129 41812
rect 3065 41668 3129 41732
rect 3065 41588 3129 41652
rect 3065 41508 3129 41572
rect 3065 41428 3129 41492
rect 3065 41348 3129 41412
rect 3065 41268 3129 41332
rect 3065 41188 3129 41252
rect 3065 41108 3129 41172
rect 3065 41028 3129 41092
rect 9384 47108 9448 47172
rect 9384 47028 9448 47092
rect 9384 46948 9448 47012
rect 9384 46868 9448 46932
rect 9384 46788 9448 46852
rect 9384 46708 9448 46772
rect 9384 46628 9448 46692
rect 9384 46548 9448 46612
rect 9384 46468 9448 46532
rect 9384 46388 9448 46452
rect 9384 46308 9448 46372
rect 9384 46228 9448 46292
rect 9384 46148 9448 46212
rect 9384 46068 9448 46132
rect 9384 45988 9448 46052
rect 9384 45908 9448 45972
rect 9384 45828 9448 45892
rect 9384 45748 9448 45812
rect 9384 45668 9448 45732
rect 9384 45588 9448 45652
rect 9384 45508 9448 45572
rect 9384 45428 9448 45492
rect 9384 45348 9448 45412
rect 9384 45268 9448 45332
rect 9384 45188 9448 45252
rect 9384 45108 9448 45172
rect 9384 45028 9448 45092
rect 9384 44948 9448 45012
rect 9384 44868 9448 44932
rect 9384 44788 9448 44852
rect 9384 44708 9448 44772
rect 9384 44628 9448 44692
rect 9384 44548 9448 44612
rect 9384 44468 9448 44532
rect 9384 44388 9448 44452
rect 9384 44308 9448 44372
rect 9384 44228 9448 44292
rect 9384 44148 9448 44212
rect 9384 44068 9448 44132
rect 9384 43988 9448 44052
rect 9384 43908 9448 43972
rect 9384 43828 9448 43892
rect 9384 43748 9448 43812
rect 9384 43668 9448 43732
rect 9384 43588 9448 43652
rect 9384 43508 9448 43572
rect 9384 43428 9448 43492
rect 9384 43348 9448 43412
rect 9384 43268 9448 43332
rect 9384 43188 9448 43252
rect 9384 43108 9448 43172
rect 9384 43028 9448 43092
rect 9384 42948 9448 43012
rect 9384 42868 9448 42932
rect 9384 42788 9448 42852
rect 9384 42708 9448 42772
rect 9384 42628 9448 42692
rect 9384 42548 9448 42612
rect 9384 42468 9448 42532
rect 9384 42388 9448 42452
rect 9384 42308 9448 42372
rect 9384 42228 9448 42292
rect 9384 42148 9448 42212
rect 9384 42068 9448 42132
rect 9384 41988 9448 42052
rect 9384 41908 9448 41972
rect 9384 41828 9448 41892
rect 9384 41748 9448 41812
rect 9384 41668 9448 41732
rect 9384 41588 9448 41652
rect 9384 41508 9448 41572
rect 9384 41428 9448 41492
rect 9384 41348 9448 41412
rect 9384 41268 9448 41332
rect 9384 41188 9448 41252
rect 9384 41108 9448 41172
rect 9384 41028 9448 41092
rect 15703 47108 15767 47172
rect 15703 47028 15767 47092
rect 15703 46948 15767 47012
rect 15703 46868 15767 46932
rect 15703 46788 15767 46852
rect 15703 46708 15767 46772
rect 15703 46628 15767 46692
rect 15703 46548 15767 46612
rect 15703 46468 15767 46532
rect 15703 46388 15767 46452
rect 15703 46308 15767 46372
rect 15703 46228 15767 46292
rect 15703 46148 15767 46212
rect 15703 46068 15767 46132
rect 15703 45988 15767 46052
rect 15703 45908 15767 45972
rect 15703 45828 15767 45892
rect 15703 45748 15767 45812
rect 15703 45668 15767 45732
rect 15703 45588 15767 45652
rect 15703 45508 15767 45572
rect 15703 45428 15767 45492
rect 15703 45348 15767 45412
rect 15703 45268 15767 45332
rect 15703 45188 15767 45252
rect 15703 45108 15767 45172
rect 15703 45028 15767 45092
rect 15703 44948 15767 45012
rect 15703 44868 15767 44932
rect 15703 44788 15767 44852
rect 15703 44708 15767 44772
rect 15703 44628 15767 44692
rect 15703 44548 15767 44612
rect 15703 44468 15767 44532
rect 15703 44388 15767 44452
rect 15703 44308 15767 44372
rect 15703 44228 15767 44292
rect 15703 44148 15767 44212
rect 15703 44068 15767 44132
rect 15703 43988 15767 44052
rect 15703 43908 15767 43972
rect 15703 43828 15767 43892
rect 15703 43748 15767 43812
rect 15703 43668 15767 43732
rect 15703 43588 15767 43652
rect 15703 43508 15767 43572
rect 15703 43428 15767 43492
rect 15703 43348 15767 43412
rect 15703 43268 15767 43332
rect 15703 43188 15767 43252
rect 15703 43108 15767 43172
rect 15703 43028 15767 43092
rect 15703 42948 15767 43012
rect 15703 42868 15767 42932
rect 15703 42788 15767 42852
rect 15703 42708 15767 42772
rect 15703 42628 15767 42692
rect 15703 42548 15767 42612
rect 15703 42468 15767 42532
rect 15703 42388 15767 42452
rect 15703 42308 15767 42372
rect 15703 42228 15767 42292
rect 15703 42148 15767 42212
rect 15703 42068 15767 42132
rect 15703 41988 15767 42052
rect 15703 41908 15767 41972
rect 15703 41828 15767 41892
rect 15703 41748 15767 41812
rect 15703 41668 15767 41732
rect 15703 41588 15767 41652
rect 15703 41508 15767 41572
rect 15703 41428 15767 41492
rect 15703 41348 15767 41412
rect 15703 41268 15767 41332
rect 15703 41188 15767 41252
rect 15703 41108 15767 41172
rect 15703 41028 15767 41092
rect 22022 47108 22086 47172
rect 22022 47028 22086 47092
rect 22022 46948 22086 47012
rect 22022 46868 22086 46932
rect 22022 46788 22086 46852
rect 22022 46708 22086 46772
rect 22022 46628 22086 46692
rect 22022 46548 22086 46612
rect 22022 46468 22086 46532
rect 22022 46388 22086 46452
rect 22022 46308 22086 46372
rect 22022 46228 22086 46292
rect 22022 46148 22086 46212
rect 22022 46068 22086 46132
rect 22022 45988 22086 46052
rect 22022 45908 22086 45972
rect 22022 45828 22086 45892
rect 22022 45748 22086 45812
rect 22022 45668 22086 45732
rect 22022 45588 22086 45652
rect 22022 45508 22086 45572
rect 22022 45428 22086 45492
rect 22022 45348 22086 45412
rect 22022 45268 22086 45332
rect 22022 45188 22086 45252
rect 22022 45108 22086 45172
rect 22022 45028 22086 45092
rect 22022 44948 22086 45012
rect 22022 44868 22086 44932
rect 22022 44788 22086 44852
rect 22022 44708 22086 44772
rect 22022 44628 22086 44692
rect 22022 44548 22086 44612
rect 22022 44468 22086 44532
rect 22022 44388 22086 44452
rect 22022 44308 22086 44372
rect 22022 44228 22086 44292
rect 22022 44148 22086 44212
rect 22022 44068 22086 44132
rect 22022 43988 22086 44052
rect 22022 43908 22086 43972
rect 22022 43828 22086 43892
rect 22022 43748 22086 43812
rect 22022 43668 22086 43732
rect 22022 43588 22086 43652
rect 22022 43508 22086 43572
rect 22022 43428 22086 43492
rect 22022 43348 22086 43412
rect 22022 43268 22086 43332
rect 22022 43188 22086 43252
rect 22022 43108 22086 43172
rect 22022 43028 22086 43092
rect 22022 42948 22086 43012
rect 22022 42868 22086 42932
rect 22022 42788 22086 42852
rect 22022 42708 22086 42772
rect 22022 42628 22086 42692
rect 22022 42548 22086 42612
rect 22022 42468 22086 42532
rect 22022 42388 22086 42452
rect 22022 42308 22086 42372
rect 22022 42228 22086 42292
rect 22022 42148 22086 42212
rect 22022 42068 22086 42132
rect 22022 41988 22086 42052
rect 22022 41908 22086 41972
rect 22022 41828 22086 41892
rect 22022 41748 22086 41812
rect 22022 41668 22086 41732
rect 22022 41588 22086 41652
rect 22022 41508 22086 41572
rect 22022 41428 22086 41492
rect 22022 41348 22086 41412
rect 22022 41268 22086 41332
rect 22022 41188 22086 41252
rect 22022 41108 22086 41172
rect 22022 41028 22086 41092
rect 28341 47108 28405 47172
rect 28341 47028 28405 47092
rect 28341 46948 28405 47012
rect 28341 46868 28405 46932
rect 28341 46788 28405 46852
rect 28341 46708 28405 46772
rect 28341 46628 28405 46692
rect 28341 46548 28405 46612
rect 28341 46468 28405 46532
rect 28341 46388 28405 46452
rect 28341 46308 28405 46372
rect 28341 46228 28405 46292
rect 28341 46148 28405 46212
rect 28341 46068 28405 46132
rect 28341 45988 28405 46052
rect 28341 45908 28405 45972
rect 28341 45828 28405 45892
rect 28341 45748 28405 45812
rect 28341 45668 28405 45732
rect 28341 45588 28405 45652
rect 28341 45508 28405 45572
rect 28341 45428 28405 45492
rect 28341 45348 28405 45412
rect 28341 45268 28405 45332
rect 28341 45188 28405 45252
rect 28341 45108 28405 45172
rect 28341 45028 28405 45092
rect 28341 44948 28405 45012
rect 28341 44868 28405 44932
rect 28341 44788 28405 44852
rect 28341 44708 28405 44772
rect 28341 44628 28405 44692
rect 28341 44548 28405 44612
rect 28341 44468 28405 44532
rect 28341 44388 28405 44452
rect 28341 44308 28405 44372
rect 28341 44228 28405 44292
rect 28341 44148 28405 44212
rect 28341 44068 28405 44132
rect 28341 43988 28405 44052
rect 28341 43908 28405 43972
rect 28341 43828 28405 43892
rect 28341 43748 28405 43812
rect 28341 43668 28405 43732
rect 28341 43588 28405 43652
rect 28341 43508 28405 43572
rect 28341 43428 28405 43492
rect 28341 43348 28405 43412
rect 28341 43268 28405 43332
rect 28341 43188 28405 43252
rect 28341 43108 28405 43172
rect 28341 43028 28405 43092
rect 28341 42948 28405 43012
rect 28341 42868 28405 42932
rect 28341 42788 28405 42852
rect 28341 42708 28405 42772
rect 28341 42628 28405 42692
rect 28341 42548 28405 42612
rect 28341 42468 28405 42532
rect 28341 42388 28405 42452
rect 28341 42308 28405 42372
rect 28341 42228 28405 42292
rect 28341 42148 28405 42212
rect 28341 42068 28405 42132
rect 28341 41988 28405 42052
rect 28341 41908 28405 41972
rect 28341 41828 28405 41892
rect 28341 41748 28405 41812
rect 28341 41668 28405 41732
rect 28341 41588 28405 41652
rect 28341 41508 28405 41572
rect 28341 41428 28405 41492
rect 28341 41348 28405 41412
rect 28341 41268 28405 41332
rect 28341 41188 28405 41252
rect 28341 41108 28405 41172
rect 28341 41028 28405 41092
rect 34660 47108 34724 47172
rect 34660 47028 34724 47092
rect 34660 46948 34724 47012
rect 34660 46868 34724 46932
rect 34660 46788 34724 46852
rect 34660 46708 34724 46772
rect 34660 46628 34724 46692
rect 34660 46548 34724 46612
rect 34660 46468 34724 46532
rect 34660 46388 34724 46452
rect 34660 46308 34724 46372
rect 34660 46228 34724 46292
rect 34660 46148 34724 46212
rect 34660 46068 34724 46132
rect 34660 45988 34724 46052
rect 34660 45908 34724 45972
rect 34660 45828 34724 45892
rect 34660 45748 34724 45812
rect 34660 45668 34724 45732
rect 34660 45588 34724 45652
rect 34660 45508 34724 45572
rect 34660 45428 34724 45492
rect 34660 45348 34724 45412
rect 34660 45268 34724 45332
rect 34660 45188 34724 45252
rect 34660 45108 34724 45172
rect 34660 45028 34724 45092
rect 34660 44948 34724 45012
rect 34660 44868 34724 44932
rect 34660 44788 34724 44852
rect 34660 44708 34724 44772
rect 34660 44628 34724 44692
rect 34660 44548 34724 44612
rect 34660 44468 34724 44532
rect 34660 44388 34724 44452
rect 34660 44308 34724 44372
rect 34660 44228 34724 44292
rect 34660 44148 34724 44212
rect 34660 44068 34724 44132
rect 34660 43988 34724 44052
rect 34660 43908 34724 43972
rect 34660 43828 34724 43892
rect 34660 43748 34724 43812
rect 34660 43668 34724 43732
rect 34660 43588 34724 43652
rect 34660 43508 34724 43572
rect 34660 43428 34724 43492
rect 34660 43348 34724 43412
rect 34660 43268 34724 43332
rect 34660 43188 34724 43252
rect 34660 43108 34724 43172
rect 34660 43028 34724 43092
rect 34660 42948 34724 43012
rect 34660 42868 34724 42932
rect 34660 42788 34724 42852
rect 34660 42708 34724 42772
rect 34660 42628 34724 42692
rect 34660 42548 34724 42612
rect 34660 42468 34724 42532
rect 34660 42388 34724 42452
rect 34660 42308 34724 42372
rect 34660 42228 34724 42292
rect 34660 42148 34724 42212
rect 34660 42068 34724 42132
rect 34660 41988 34724 42052
rect 34660 41908 34724 41972
rect 34660 41828 34724 41892
rect 34660 41748 34724 41812
rect 34660 41668 34724 41732
rect 34660 41588 34724 41652
rect 34660 41508 34724 41572
rect 34660 41428 34724 41492
rect 34660 41348 34724 41412
rect 34660 41268 34724 41332
rect 34660 41188 34724 41252
rect 34660 41108 34724 41172
rect 34660 41028 34724 41092
rect 40979 47108 41043 47172
rect 40979 47028 41043 47092
rect 40979 46948 41043 47012
rect 40979 46868 41043 46932
rect 40979 46788 41043 46852
rect 40979 46708 41043 46772
rect 40979 46628 41043 46692
rect 40979 46548 41043 46612
rect 40979 46468 41043 46532
rect 40979 46388 41043 46452
rect 40979 46308 41043 46372
rect 40979 46228 41043 46292
rect 40979 46148 41043 46212
rect 40979 46068 41043 46132
rect 40979 45988 41043 46052
rect 40979 45908 41043 45972
rect 40979 45828 41043 45892
rect 40979 45748 41043 45812
rect 40979 45668 41043 45732
rect 40979 45588 41043 45652
rect 40979 45508 41043 45572
rect 40979 45428 41043 45492
rect 40979 45348 41043 45412
rect 40979 45268 41043 45332
rect 40979 45188 41043 45252
rect 40979 45108 41043 45172
rect 40979 45028 41043 45092
rect 40979 44948 41043 45012
rect 40979 44868 41043 44932
rect 40979 44788 41043 44852
rect 40979 44708 41043 44772
rect 40979 44628 41043 44692
rect 40979 44548 41043 44612
rect 40979 44468 41043 44532
rect 40979 44388 41043 44452
rect 40979 44308 41043 44372
rect 40979 44228 41043 44292
rect 40979 44148 41043 44212
rect 40979 44068 41043 44132
rect 40979 43988 41043 44052
rect 40979 43908 41043 43972
rect 40979 43828 41043 43892
rect 40979 43748 41043 43812
rect 40979 43668 41043 43732
rect 40979 43588 41043 43652
rect 40979 43508 41043 43572
rect 40979 43428 41043 43492
rect 40979 43348 41043 43412
rect 40979 43268 41043 43332
rect 40979 43188 41043 43252
rect 40979 43108 41043 43172
rect 40979 43028 41043 43092
rect 40979 42948 41043 43012
rect 40979 42868 41043 42932
rect 40979 42788 41043 42852
rect 40979 42708 41043 42772
rect 40979 42628 41043 42692
rect 40979 42548 41043 42612
rect 40979 42468 41043 42532
rect 40979 42388 41043 42452
rect 40979 42308 41043 42372
rect 40979 42228 41043 42292
rect 40979 42148 41043 42212
rect 40979 42068 41043 42132
rect 40979 41988 41043 42052
rect 40979 41908 41043 41972
rect 40979 41828 41043 41892
rect 40979 41748 41043 41812
rect 40979 41668 41043 41732
rect 40979 41588 41043 41652
rect 40979 41508 41043 41572
rect 40979 41428 41043 41492
rect 40979 41348 41043 41412
rect 40979 41268 41043 41332
rect 40979 41188 41043 41252
rect 40979 41108 41043 41172
rect 40979 41028 41043 41092
rect 47298 47108 47362 47172
rect 47298 47028 47362 47092
rect 47298 46948 47362 47012
rect 47298 46868 47362 46932
rect 47298 46788 47362 46852
rect 47298 46708 47362 46772
rect 47298 46628 47362 46692
rect 47298 46548 47362 46612
rect 47298 46468 47362 46532
rect 47298 46388 47362 46452
rect 47298 46308 47362 46372
rect 47298 46228 47362 46292
rect 47298 46148 47362 46212
rect 47298 46068 47362 46132
rect 47298 45988 47362 46052
rect 47298 45908 47362 45972
rect 47298 45828 47362 45892
rect 47298 45748 47362 45812
rect 47298 45668 47362 45732
rect 47298 45588 47362 45652
rect 47298 45508 47362 45572
rect 47298 45428 47362 45492
rect 47298 45348 47362 45412
rect 47298 45268 47362 45332
rect 47298 45188 47362 45252
rect 47298 45108 47362 45172
rect 47298 45028 47362 45092
rect 47298 44948 47362 45012
rect 47298 44868 47362 44932
rect 47298 44788 47362 44852
rect 47298 44708 47362 44772
rect 47298 44628 47362 44692
rect 47298 44548 47362 44612
rect 47298 44468 47362 44532
rect 47298 44388 47362 44452
rect 47298 44308 47362 44372
rect 47298 44228 47362 44292
rect 47298 44148 47362 44212
rect 47298 44068 47362 44132
rect 47298 43988 47362 44052
rect 47298 43908 47362 43972
rect 47298 43828 47362 43892
rect 47298 43748 47362 43812
rect 47298 43668 47362 43732
rect 47298 43588 47362 43652
rect 47298 43508 47362 43572
rect 47298 43428 47362 43492
rect 47298 43348 47362 43412
rect 47298 43268 47362 43332
rect 47298 43188 47362 43252
rect 47298 43108 47362 43172
rect 47298 43028 47362 43092
rect 47298 42948 47362 43012
rect 47298 42868 47362 42932
rect 47298 42788 47362 42852
rect 47298 42708 47362 42772
rect 47298 42628 47362 42692
rect 47298 42548 47362 42612
rect 47298 42468 47362 42532
rect 47298 42388 47362 42452
rect 47298 42308 47362 42372
rect 47298 42228 47362 42292
rect 47298 42148 47362 42212
rect 47298 42068 47362 42132
rect 47298 41988 47362 42052
rect 47298 41908 47362 41972
rect 47298 41828 47362 41892
rect 47298 41748 47362 41812
rect 47298 41668 47362 41732
rect 47298 41588 47362 41652
rect 47298 41508 47362 41572
rect 47298 41428 47362 41492
rect 47298 41348 47362 41412
rect 47298 41268 47362 41332
rect 47298 41188 47362 41252
rect 47298 41108 47362 41172
rect 47298 41028 47362 41092
rect -41168 40808 -41104 40872
rect -41168 40728 -41104 40792
rect -41168 40648 -41104 40712
rect -41168 40568 -41104 40632
rect -41168 40488 -41104 40552
rect -41168 40408 -41104 40472
rect -41168 40328 -41104 40392
rect -41168 40248 -41104 40312
rect -41168 40168 -41104 40232
rect -41168 40088 -41104 40152
rect -41168 40008 -41104 40072
rect -41168 39928 -41104 39992
rect -41168 39848 -41104 39912
rect -41168 39768 -41104 39832
rect -41168 39688 -41104 39752
rect -41168 39608 -41104 39672
rect -41168 39528 -41104 39592
rect -41168 39448 -41104 39512
rect -41168 39368 -41104 39432
rect -41168 39288 -41104 39352
rect -41168 39208 -41104 39272
rect -41168 39128 -41104 39192
rect -41168 39048 -41104 39112
rect -41168 38968 -41104 39032
rect -41168 38888 -41104 38952
rect -41168 38808 -41104 38872
rect -41168 38728 -41104 38792
rect -41168 38648 -41104 38712
rect -41168 38568 -41104 38632
rect -41168 38488 -41104 38552
rect -41168 38408 -41104 38472
rect -41168 38328 -41104 38392
rect -41168 38248 -41104 38312
rect -41168 38168 -41104 38232
rect -41168 38088 -41104 38152
rect -41168 38008 -41104 38072
rect -41168 37928 -41104 37992
rect -41168 37848 -41104 37912
rect -41168 37768 -41104 37832
rect -41168 37688 -41104 37752
rect -41168 37608 -41104 37672
rect -41168 37528 -41104 37592
rect -41168 37448 -41104 37512
rect -41168 37368 -41104 37432
rect -41168 37288 -41104 37352
rect -41168 37208 -41104 37272
rect -41168 37128 -41104 37192
rect -41168 37048 -41104 37112
rect -41168 36968 -41104 37032
rect -41168 36888 -41104 36952
rect -41168 36808 -41104 36872
rect -41168 36728 -41104 36792
rect -41168 36648 -41104 36712
rect -41168 36568 -41104 36632
rect -41168 36488 -41104 36552
rect -41168 36408 -41104 36472
rect -41168 36328 -41104 36392
rect -41168 36248 -41104 36312
rect -41168 36168 -41104 36232
rect -41168 36088 -41104 36152
rect -41168 36008 -41104 36072
rect -41168 35928 -41104 35992
rect -41168 35848 -41104 35912
rect -41168 35768 -41104 35832
rect -41168 35688 -41104 35752
rect -41168 35608 -41104 35672
rect -41168 35528 -41104 35592
rect -41168 35448 -41104 35512
rect -41168 35368 -41104 35432
rect -41168 35288 -41104 35352
rect -41168 35208 -41104 35272
rect -41168 35128 -41104 35192
rect -41168 35048 -41104 35112
rect -41168 34968 -41104 35032
rect -41168 34888 -41104 34952
rect -41168 34808 -41104 34872
rect -41168 34728 -41104 34792
rect -34849 40808 -34785 40872
rect -34849 40728 -34785 40792
rect -34849 40648 -34785 40712
rect -34849 40568 -34785 40632
rect -34849 40488 -34785 40552
rect -34849 40408 -34785 40472
rect -34849 40328 -34785 40392
rect -34849 40248 -34785 40312
rect -34849 40168 -34785 40232
rect -34849 40088 -34785 40152
rect -34849 40008 -34785 40072
rect -34849 39928 -34785 39992
rect -34849 39848 -34785 39912
rect -34849 39768 -34785 39832
rect -34849 39688 -34785 39752
rect -34849 39608 -34785 39672
rect -34849 39528 -34785 39592
rect -34849 39448 -34785 39512
rect -34849 39368 -34785 39432
rect -34849 39288 -34785 39352
rect -34849 39208 -34785 39272
rect -34849 39128 -34785 39192
rect -34849 39048 -34785 39112
rect -34849 38968 -34785 39032
rect -34849 38888 -34785 38952
rect -34849 38808 -34785 38872
rect -34849 38728 -34785 38792
rect -34849 38648 -34785 38712
rect -34849 38568 -34785 38632
rect -34849 38488 -34785 38552
rect -34849 38408 -34785 38472
rect -34849 38328 -34785 38392
rect -34849 38248 -34785 38312
rect -34849 38168 -34785 38232
rect -34849 38088 -34785 38152
rect -34849 38008 -34785 38072
rect -34849 37928 -34785 37992
rect -34849 37848 -34785 37912
rect -34849 37768 -34785 37832
rect -34849 37688 -34785 37752
rect -34849 37608 -34785 37672
rect -34849 37528 -34785 37592
rect -34849 37448 -34785 37512
rect -34849 37368 -34785 37432
rect -34849 37288 -34785 37352
rect -34849 37208 -34785 37272
rect -34849 37128 -34785 37192
rect -34849 37048 -34785 37112
rect -34849 36968 -34785 37032
rect -34849 36888 -34785 36952
rect -34849 36808 -34785 36872
rect -34849 36728 -34785 36792
rect -34849 36648 -34785 36712
rect -34849 36568 -34785 36632
rect -34849 36488 -34785 36552
rect -34849 36408 -34785 36472
rect -34849 36328 -34785 36392
rect -34849 36248 -34785 36312
rect -34849 36168 -34785 36232
rect -34849 36088 -34785 36152
rect -34849 36008 -34785 36072
rect -34849 35928 -34785 35992
rect -34849 35848 -34785 35912
rect -34849 35768 -34785 35832
rect -34849 35688 -34785 35752
rect -34849 35608 -34785 35672
rect -34849 35528 -34785 35592
rect -34849 35448 -34785 35512
rect -34849 35368 -34785 35432
rect -34849 35288 -34785 35352
rect -34849 35208 -34785 35272
rect -34849 35128 -34785 35192
rect -34849 35048 -34785 35112
rect -34849 34968 -34785 35032
rect -34849 34888 -34785 34952
rect -34849 34808 -34785 34872
rect -34849 34728 -34785 34792
rect -28530 40808 -28466 40872
rect -28530 40728 -28466 40792
rect -28530 40648 -28466 40712
rect -28530 40568 -28466 40632
rect -28530 40488 -28466 40552
rect -28530 40408 -28466 40472
rect -28530 40328 -28466 40392
rect -28530 40248 -28466 40312
rect -28530 40168 -28466 40232
rect -28530 40088 -28466 40152
rect -28530 40008 -28466 40072
rect -28530 39928 -28466 39992
rect -28530 39848 -28466 39912
rect -28530 39768 -28466 39832
rect -28530 39688 -28466 39752
rect -28530 39608 -28466 39672
rect -28530 39528 -28466 39592
rect -28530 39448 -28466 39512
rect -28530 39368 -28466 39432
rect -28530 39288 -28466 39352
rect -28530 39208 -28466 39272
rect -28530 39128 -28466 39192
rect -28530 39048 -28466 39112
rect -28530 38968 -28466 39032
rect -28530 38888 -28466 38952
rect -28530 38808 -28466 38872
rect -28530 38728 -28466 38792
rect -28530 38648 -28466 38712
rect -28530 38568 -28466 38632
rect -28530 38488 -28466 38552
rect -28530 38408 -28466 38472
rect -28530 38328 -28466 38392
rect -28530 38248 -28466 38312
rect -28530 38168 -28466 38232
rect -28530 38088 -28466 38152
rect -28530 38008 -28466 38072
rect -28530 37928 -28466 37992
rect -28530 37848 -28466 37912
rect -28530 37768 -28466 37832
rect -28530 37688 -28466 37752
rect -28530 37608 -28466 37672
rect -28530 37528 -28466 37592
rect -28530 37448 -28466 37512
rect -28530 37368 -28466 37432
rect -28530 37288 -28466 37352
rect -28530 37208 -28466 37272
rect -28530 37128 -28466 37192
rect -28530 37048 -28466 37112
rect -28530 36968 -28466 37032
rect -28530 36888 -28466 36952
rect -28530 36808 -28466 36872
rect -28530 36728 -28466 36792
rect -28530 36648 -28466 36712
rect -28530 36568 -28466 36632
rect -28530 36488 -28466 36552
rect -28530 36408 -28466 36472
rect -28530 36328 -28466 36392
rect -28530 36248 -28466 36312
rect -28530 36168 -28466 36232
rect -28530 36088 -28466 36152
rect -28530 36008 -28466 36072
rect -28530 35928 -28466 35992
rect -28530 35848 -28466 35912
rect -28530 35768 -28466 35832
rect -28530 35688 -28466 35752
rect -28530 35608 -28466 35672
rect -28530 35528 -28466 35592
rect -28530 35448 -28466 35512
rect -28530 35368 -28466 35432
rect -28530 35288 -28466 35352
rect -28530 35208 -28466 35272
rect -28530 35128 -28466 35192
rect -28530 35048 -28466 35112
rect -28530 34968 -28466 35032
rect -28530 34888 -28466 34952
rect -28530 34808 -28466 34872
rect -28530 34728 -28466 34792
rect -22211 40808 -22147 40872
rect -22211 40728 -22147 40792
rect -22211 40648 -22147 40712
rect -22211 40568 -22147 40632
rect -22211 40488 -22147 40552
rect -22211 40408 -22147 40472
rect -22211 40328 -22147 40392
rect -22211 40248 -22147 40312
rect -22211 40168 -22147 40232
rect -22211 40088 -22147 40152
rect -22211 40008 -22147 40072
rect -22211 39928 -22147 39992
rect -22211 39848 -22147 39912
rect -22211 39768 -22147 39832
rect -22211 39688 -22147 39752
rect -22211 39608 -22147 39672
rect -22211 39528 -22147 39592
rect -22211 39448 -22147 39512
rect -22211 39368 -22147 39432
rect -22211 39288 -22147 39352
rect -22211 39208 -22147 39272
rect -22211 39128 -22147 39192
rect -22211 39048 -22147 39112
rect -22211 38968 -22147 39032
rect -22211 38888 -22147 38952
rect -22211 38808 -22147 38872
rect -22211 38728 -22147 38792
rect -22211 38648 -22147 38712
rect -22211 38568 -22147 38632
rect -22211 38488 -22147 38552
rect -22211 38408 -22147 38472
rect -22211 38328 -22147 38392
rect -22211 38248 -22147 38312
rect -22211 38168 -22147 38232
rect -22211 38088 -22147 38152
rect -22211 38008 -22147 38072
rect -22211 37928 -22147 37992
rect -22211 37848 -22147 37912
rect -22211 37768 -22147 37832
rect -22211 37688 -22147 37752
rect -22211 37608 -22147 37672
rect -22211 37528 -22147 37592
rect -22211 37448 -22147 37512
rect -22211 37368 -22147 37432
rect -22211 37288 -22147 37352
rect -22211 37208 -22147 37272
rect -22211 37128 -22147 37192
rect -22211 37048 -22147 37112
rect -22211 36968 -22147 37032
rect -22211 36888 -22147 36952
rect -22211 36808 -22147 36872
rect -22211 36728 -22147 36792
rect -22211 36648 -22147 36712
rect -22211 36568 -22147 36632
rect -22211 36488 -22147 36552
rect -22211 36408 -22147 36472
rect -22211 36328 -22147 36392
rect -22211 36248 -22147 36312
rect -22211 36168 -22147 36232
rect -22211 36088 -22147 36152
rect -22211 36008 -22147 36072
rect -22211 35928 -22147 35992
rect -22211 35848 -22147 35912
rect -22211 35768 -22147 35832
rect -22211 35688 -22147 35752
rect -22211 35608 -22147 35672
rect -22211 35528 -22147 35592
rect -22211 35448 -22147 35512
rect -22211 35368 -22147 35432
rect -22211 35288 -22147 35352
rect -22211 35208 -22147 35272
rect -22211 35128 -22147 35192
rect -22211 35048 -22147 35112
rect -22211 34968 -22147 35032
rect -22211 34888 -22147 34952
rect -22211 34808 -22147 34872
rect -22211 34728 -22147 34792
rect -15892 40808 -15828 40872
rect -15892 40728 -15828 40792
rect -15892 40648 -15828 40712
rect -15892 40568 -15828 40632
rect -15892 40488 -15828 40552
rect -15892 40408 -15828 40472
rect -15892 40328 -15828 40392
rect -15892 40248 -15828 40312
rect -15892 40168 -15828 40232
rect -15892 40088 -15828 40152
rect -15892 40008 -15828 40072
rect -15892 39928 -15828 39992
rect -15892 39848 -15828 39912
rect -15892 39768 -15828 39832
rect -15892 39688 -15828 39752
rect -15892 39608 -15828 39672
rect -15892 39528 -15828 39592
rect -15892 39448 -15828 39512
rect -15892 39368 -15828 39432
rect -15892 39288 -15828 39352
rect -15892 39208 -15828 39272
rect -15892 39128 -15828 39192
rect -15892 39048 -15828 39112
rect -15892 38968 -15828 39032
rect -15892 38888 -15828 38952
rect -15892 38808 -15828 38872
rect -15892 38728 -15828 38792
rect -15892 38648 -15828 38712
rect -15892 38568 -15828 38632
rect -15892 38488 -15828 38552
rect -15892 38408 -15828 38472
rect -15892 38328 -15828 38392
rect -15892 38248 -15828 38312
rect -15892 38168 -15828 38232
rect -15892 38088 -15828 38152
rect -15892 38008 -15828 38072
rect -15892 37928 -15828 37992
rect -15892 37848 -15828 37912
rect -15892 37768 -15828 37832
rect -15892 37688 -15828 37752
rect -15892 37608 -15828 37672
rect -15892 37528 -15828 37592
rect -15892 37448 -15828 37512
rect -15892 37368 -15828 37432
rect -15892 37288 -15828 37352
rect -15892 37208 -15828 37272
rect -15892 37128 -15828 37192
rect -15892 37048 -15828 37112
rect -15892 36968 -15828 37032
rect -15892 36888 -15828 36952
rect -15892 36808 -15828 36872
rect -15892 36728 -15828 36792
rect -15892 36648 -15828 36712
rect -15892 36568 -15828 36632
rect -15892 36488 -15828 36552
rect -15892 36408 -15828 36472
rect -15892 36328 -15828 36392
rect -15892 36248 -15828 36312
rect -15892 36168 -15828 36232
rect -15892 36088 -15828 36152
rect -15892 36008 -15828 36072
rect -15892 35928 -15828 35992
rect -15892 35848 -15828 35912
rect -15892 35768 -15828 35832
rect -15892 35688 -15828 35752
rect -15892 35608 -15828 35672
rect -15892 35528 -15828 35592
rect -15892 35448 -15828 35512
rect -15892 35368 -15828 35432
rect -15892 35288 -15828 35352
rect -15892 35208 -15828 35272
rect -15892 35128 -15828 35192
rect -15892 35048 -15828 35112
rect -15892 34968 -15828 35032
rect -15892 34888 -15828 34952
rect -15892 34808 -15828 34872
rect -15892 34728 -15828 34792
rect -9573 40808 -9509 40872
rect -9573 40728 -9509 40792
rect -9573 40648 -9509 40712
rect -9573 40568 -9509 40632
rect -9573 40488 -9509 40552
rect -9573 40408 -9509 40472
rect -9573 40328 -9509 40392
rect -9573 40248 -9509 40312
rect -9573 40168 -9509 40232
rect -9573 40088 -9509 40152
rect -9573 40008 -9509 40072
rect -9573 39928 -9509 39992
rect -9573 39848 -9509 39912
rect -9573 39768 -9509 39832
rect -9573 39688 -9509 39752
rect -9573 39608 -9509 39672
rect -9573 39528 -9509 39592
rect -9573 39448 -9509 39512
rect -9573 39368 -9509 39432
rect -9573 39288 -9509 39352
rect -9573 39208 -9509 39272
rect -9573 39128 -9509 39192
rect -9573 39048 -9509 39112
rect -9573 38968 -9509 39032
rect -9573 38888 -9509 38952
rect -9573 38808 -9509 38872
rect -9573 38728 -9509 38792
rect -9573 38648 -9509 38712
rect -9573 38568 -9509 38632
rect -9573 38488 -9509 38552
rect -9573 38408 -9509 38472
rect -9573 38328 -9509 38392
rect -9573 38248 -9509 38312
rect -9573 38168 -9509 38232
rect -9573 38088 -9509 38152
rect -9573 38008 -9509 38072
rect -9573 37928 -9509 37992
rect -9573 37848 -9509 37912
rect -9573 37768 -9509 37832
rect -9573 37688 -9509 37752
rect -9573 37608 -9509 37672
rect -9573 37528 -9509 37592
rect -9573 37448 -9509 37512
rect -9573 37368 -9509 37432
rect -9573 37288 -9509 37352
rect -9573 37208 -9509 37272
rect -9573 37128 -9509 37192
rect -9573 37048 -9509 37112
rect -9573 36968 -9509 37032
rect -9573 36888 -9509 36952
rect -9573 36808 -9509 36872
rect -9573 36728 -9509 36792
rect -9573 36648 -9509 36712
rect -9573 36568 -9509 36632
rect -9573 36488 -9509 36552
rect -9573 36408 -9509 36472
rect -9573 36328 -9509 36392
rect -9573 36248 -9509 36312
rect -9573 36168 -9509 36232
rect -9573 36088 -9509 36152
rect -9573 36008 -9509 36072
rect -9573 35928 -9509 35992
rect -9573 35848 -9509 35912
rect -9573 35768 -9509 35832
rect -9573 35688 -9509 35752
rect -9573 35608 -9509 35672
rect -9573 35528 -9509 35592
rect -9573 35448 -9509 35512
rect -9573 35368 -9509 35432
rect -9573 35288 -9509 35352
rect -9573 35208 -9509 35272
rect -9573 35128 -9509 35192
rect -9573 35048 -9509 35112
rect -9573 34968 -9509 35032
rect -9573 34888 -9509 34952
rect -9573 34808 -9509 34872
rect -9573 34728 -9509 34792
rect -3254 40808 -3190 40872
rect -3254 40728 -3190 40792
rect -3254 40648 -3190 40712
rect -3254 40568 -3190 40632
rect -3254 40488 -3190 40552
rect -3254 40408 -3190 40472
rect -3254 40328 -3190 40392
rect -3254 40248 -3190 40312
rect -3254 40168 -3190 40232
rect -3254 40088 -3190 40152
rect -3254 40008 -3190 40072
rect -3254 39928 -3190 39992
rect -3254 39848 -3190 39912
rect -3254 39768 -3190 39832
rect -3254 39688 -3190 39752
rect -3254 39608 -3190 39672
rect -3254 39528 -3190 39592
rect -3254 39448 -3190 39512
rect -3254 39368 -3190 39432
rect -3254 39288 -3190 39352
rect -3254 39208 -3190 39272
rect -3254 39128 -3190 39192
rect -3254 39048 -3190 39112
rect -3254 38968 -3190 39032
rect -3254 38888 -3190 38952
rect -3254 38808 -3190 38872
rect -3254 38728 -3190 38792
rect -3254 38648 -3190 38712
rect -3254 38568 -3190 38632
rect -3254 38488 -3190 38552
rect -3254 38408 -3190 38472
rect -3254 38328 -3190 38392
rect -3254 38248 -3190 38312
rect -3254 38168 -3190 38232
rect -3254 38088 -3190 38152
rect -3254 38008 -3190 38072
rect -3254 37928 -3190 37992
rect -3254 37848 -3190 37912
rect -3254 37768 -3190 37832
rect -3254 37688 -3190 37752
rect -3254 37608 -3190 37672
rect -3254 37528 -3190 37592
rect -3254 37448 -3190 37512
rect -3254 37368 -3190 37432
rect -3254 37288 -3190 37352
rect -3254 37208 -3190 37272
rect -3254 37128 -3190 37192
rect -3254 37048 -3190 37112
rect -3254 36968 -3190 37032
rect -3254 36888 -3190 36952
rect -3254 36808 -3190 36872
rect -3254 36728 -3190 36792
rect -3254 36648 -3190 36712
rect -3254 36568 -3190 36632
rect -3254 36488 -3190 36552
rect -3254 36408 -3190 36472
rect -3254 36328 -3190 36392
rect -3254 36248 -3190 36312
rect -3254 36168 -3190 36232
rect -3254 36088 -3190 36152
rect -3254 36008 -3190 36072
rect -3254 35928 -3190 35992
rect -3254 35848 -3190 35912
rect -3254 35768 -3190 35832
rect -3254 35688 -3190 35752
rect -3254 35608 -3190 35672
rect -3254 35528 -3190 35592
rect -3254 35448 -3190 35512
rect -3254 35368 -3190 35432
rect -3254 35288 -3190 35352
rect -3254 35208 -3190 35272
rect -3254 35128 -3190 35192
rect -3254 35048 -3190 35112
rect -3254 34968 -3190 35032
rect -3254 34888 -3190 34952
rect -3254 34808 -3190 34872
rect -3254 34728 -3190 34792
rect 3065 40808 3129 40872
rect 3065 40728 3129 40792
rect 3065 40648 3129 40712
rect 3065 40568 3129 40632
rect 3065 40488 3129 40552
rect 3065 40408 3129 40472
rect 3065 40328 3129 40392
rect 3065 40248 3129 40312
rect 3065 40168 3129 40232
rect 3065 40088 3129 40152
rect 3065 40008 3129 40072
rect 3065 39928 3129 39992
rect 3065 39848 3129 39912
rect 3065 39768 3129 39832
rect 3065 39688 3129 39752
rect 3065 39608 3129 39672
rect 3065 39528 3129 39592
rect 3065 39448 3129 39512
rect 3065 39368 3129 39432
rect 3065 39288 3129 39352
rect 3065 39208 3129 39272
rect 3065 39128 3129 39192
rect 3065 39048 3129 39112
rect 3065 38968 3129 39032
rect 3065 38888 3129 38952
rect 3065 38808 3129 38872
rect 3065 38728 3129 38792
rect 3065 38648 3129 38712
rect 3065 38568 3129 38632
rect 3065 38488 3129 38552
rect 3065 38408 3129 38472
rect 3065 38328 3129 38392
rect 3065 38248 3129 38312
rect 3065 38168 3129 38232
rect 3065 38088 3129 38152
rect 3065 38008 3129 38072
rect 3065 37928 3129 37992
rect 3065 37848 3129 37912
rect 3065 37768 3129 37832
rect 3065 37688 3129 37752
rect 3065 37608 3129 37672
rect 3065 37528 3129 37592
rect 3065 37448 3129 37512
rect 3065 37368 3129 37432
rect 3065 37288 3129 37352
rect 3065 37208 3129 37272
rect 3065 37128 3129 37192
rect 3065 37048 3129 37112
rect 3065 36968 3129 37032
rect 3065 36888 3129 36952
rect 3065 36808 3129 36872
rect 3065 36728 3129 36792
rect 3065 36648 3129 36712
rect 3065 36568 3129 36632
rect 3065 36488 3129 36552
rect 3065 36408 3129 36472
rect 3065 36328 3129 36392
rect 3065 36248 3129 36312
rect 3065 36168 3129 36232
rect 3065 36088 3129 36152
rect 3065 36008 3129 36072
rect 3065 35928 3129 35992
rect 3065 35848 3129 35912
rect 3065 35768 3129 35832
rect 3065 35688 3129 35752
rect 3065 35608 3129 35672
rect 3065 35528 3129 35592
rect 3065 35448 3129 35512
rect 3065 35368 3129 35432
rect 3065 35288 3129 35352
rect 3065 35208 3129 35272
rect 3065 35128 3129 35192
rect 3065 35048 3129 35112
rect 3065 34968 3129 35032
rect 3065 34888 3129 34952
rect 3065 34808 3129 34872
rect 3065 34728 3129 34792
rect 9384 40808 9448 40872
rect 9384 40728 9448 40792
rect 9384 40648 9448 40712
rect 9384 40568 9448 40632
rect 9384 40488 9448 40552
rect 9384 40408 9448 40472
rect 9384 40328 9448 40392
rect 9384 40248 9448 40312
rect 9384 40168 9448 40232
rect 9384 40088 9448 40152
rect 9384 40008 9448 40072
rect 9384 39928 9448 39992
rect 9384 39848 9448 39912
rect 9384 39768 9448 39832
rect 9384 39688 9448 39752
rect 9384 39608 9448 39672
rect 9384 39528 9448 39592
rect 9384 39448 9448 39512
rect 9384 39368 9448 39432
rect 9384 39288 9448 39352
rect 9384 39208 9448 39272
rect 9384 39128 9448 39192
rect 9384 39048 9448 39112
rect 9384 38968 9448 39032
rect 9384 38888 9448 38952
rect 9384 38808 9448 38872
rect 9384 38728 9448 38792
rect 9384 38648 9448 38712
rect 9384 38568 9448 38632
rect 9384 38488 9448 38552
rect 9384 38408 9448 38472
rect 9384 38328 9448 38392
rect 9384 38248 9448 38312
rect 9384 38168 9448 38232
rect 9384 38088 9448 38152
rect 9384 38008 9448 38072
rect 9384 37928 9448 37992
rect 9384 37848 9448 37912
rect 9384 37768 9448 37832
rect 9384 37688 9448 37752
rect 9384 37608 9448 37672
rect 9384 37528 9448 37592
rect 9384 37448 9448 37512
rect 9384 37368 9448 37432
rect 9384 37288 9448 37352
rect 9384 37208 9448 37272
rect 9384 37128 9448 37192
rect 9384 37048 9448 37112
rect 9384 36968 9448 37032
rect 9384 36888 9448 36952
rect 9384 36808 9448 36872
rect 9384 36728 9448 36792
rect 9384 36648 9448 36712
rect 9384 36568 9448 36632
rect 9384 36488 9448 36552
rect 9384 36408 9448 36472
rect 9384 36328 9448 36392
rect 9384 36248 9448 36312
rect 9384 36168 9448 36232
rect 9384 36088 9448 36152
rect 9384 36008 9448 36072
rect 9384 35928 9448 35992
rect 9384 35848 9448 35912
rect 9384 35768 9448 35832
rect 9384 35688 9448 35752
rect 9384 35608 9448 35672
rect 9384 35528 9448 35592
rect 9384 35448 9448 35512
rect 9384 35368 9448 35432
rect 9384 35288 9448 35352
rect 9384 35208 9448 35272
rect 9384 35128 9448 35192
rect 9384 35048 9448 35112
rect 9384 34968 9448 35032
rect 9384 34888 9448 34952
rect 9384 34808 9448 34872
rect 9384 34728 9448 34792
rect 15703 40808 15767 40872
rect 15703 40728 15767 40792
rect 15703 40648 15767 40712
rect 15703 40568 15767 40632
rect 15703 40488 15767 40552
rect 15703 40408 15767 40472
rect 15703 40328 15767 40392
rect 15703 40248 15767 40312
rect 15703 40168 15767 40232
rect 15703 40088 15767 40152
rect 15703 40008 15767 40072
rect 15703 39928 15767 39992
rect 15703 39848 15767 39912
rect 15703 39768 15767 39832
rect 15703 39688 15767 39752
rect 15703 39608 15767 39672
rect 15703 39528 15767 39592
rect 15703 39448 15767 39512
rect 15703 39368 15767 39432
rect 15703 39288 15767 39352
rect 15703 39208 15767 39272
rect 15703 39128 15767 39192
rect 15703 39048 15767 39112
rect 15703 38968 15767 39032
rect 15703 38888 15767 38952
rect 15703 38808 15767 38872
rect 15703 38728 15767 38792
rect 15703 38648 15767 38712
rect 15703 38568 15767 38632
rect 15703 38488 15767 38552
rect 15703 38408 15767 38472
rect 15703 38328 15767 38392
rect 15703 38248 15767 38312
rect 15703 38168 15767 38232
rect 15703 38088 15767 38152
rect 15703 38008 15767 38072
rect 15703 37928 15767 37992
rect 15703 37848 15767 37912
rect 15703 37768 15767 37832
rect 15703 37688 15767 37752
rect 15703 37608 15767 37672
rect 15703 37528 15767 37592
rect 15703 37448 15767 37512
rect 15703 37368 15767 37432
rect 15703 37288 15767 37352
rect 15703 37208 15767 37272
rect 15703 37128 15767 37192
rect 15703 37048 15767 37112
rect 15703 36968 15767 37032
rect 15703 36888 15767 36952
rect 15703 36808 15767 36872
rect 15703 36728 15767 36792
rect 15703 36648 15767 36712
rect 15703 36568 15767 36632
rect 15703 36488 15767 36552
rect 15703 36408 15767 36472
rect 15703 36328 15767 36392
rect 15703 36248 15767 36312
rect 15703 36168 15767 36232
rect 15703 36088 15767 36152
rect 15703 36008 15767 36072
rect 15703 35928 15767 35992
rect 15703 35848 15767 35912
rect 15703 35768 15767 35832
rect 15703 35688 15767 35752
rect 15703 35608 15767 35672
rect 15703 35528 15767 35592
rect 15703 35448 15767 35512
rect 15703 35368 15767 35432
rect 15703 35288 15767 35352
rect 15703 35208 15767 35272
rect 15703 35128 15767 35192
rect 15703 35048 15767 35112
rect 15703 34968 15767 35032
rect 15703 34888 15767 34952
rect 15703 34808 15767 34872
rect 15703 34728 15767 34792
rect 22022 40808 22086 40872
rect 22022 40728 22086 40792
rect 22022 40648 22086 40712
rect 22022 40568 22086 40632
rect 22022 40488 22086 40552
rect 22022 40408 22086 40472
rect 22022 40328 22086 40392
rect 22022 40248 22086 40312
rect 22022 40168 22086 40232
rect 22022 40088 22086 40152
rect 22022 40008 22086 40072
rect 22022 39928 22086 39992
rect 22022 39848 22086 39912
rect 22022 39768 22086 39832
rect 22022 39688 22086 39752
rect 22022 39608 22086 39672
rect 22022 39528 22086 39592
rect 22022 39448 22086 39512
rect 22022 39368 22086 39432
rect 22022 39288 22086 39352
rect 22022 39208 22086 39272
rect 22022 39128 22086 39192
rect 22022 39048 22086 39112
rect 22022 38968 22086 39032
rect 22022 38888 22086 38952
rect 22022 38808 22086 38872
rect 22022 38728 22086 38792
rect 22022 38648 22086 38712
rect 22022 38568 22086 38632
rect 22022 38488 22086 38552
rect 22022 38408 22086 38472
rect 22022 38328 22086 38392
rect 22022 38248 22086 38312
rect 22022 38168 22086 38232
rect 22022 38088 22086 38152
rect 22022 38008 22086 38072
rect 22022 37928 22086 37992
rect 22022 37848 22086 37912
rect 22022 37768 22086 37832
rect 22022 37688 22086 37752
rect 22022 37608 22086 37672
rect 22022 37528 22086 37592
rect 22022 37448 22086 37512
rect 22022 37368 22086 37432
rect 22022 37288 22086 37352
rect 22022 37208 22086 37272
rect 22022 37128 22086 37192
rect 22022 37048 22086 37112
rect 22022 36968 22086 37032
rect 22022 36888 22086 36952
rect 22022 36808 22086 36872
rect 22022 36728 22086 36792
rect 22022 36648 22086 36712
rect 22022 36568 22086 36632
rect 22022 36488 22086 36552
rect 22022 36408 22086 36472
rect 22022 36328 22086 36392
rect 22022 36248 22086 36312
rect 22022 36168 22086 36232
rect 22022 36088 22086 36152
rect 22022 36008 22086 36072
rect 22022 35928 22086 35992
rect 22022 35848 22086 35912
rect 22022 35768 22086 35832
rect 22022 35688 22086 35752
rect 22022 35608 22086 35672
rect 22022 35528 22086 35592
rect 22022 35448 22086 35512
rect 22022 35368 22086 35432
rect 22022 35288 22086 35352
rect 22022 35208 22086 35272
rect 22022 35128 22086 35192
rect 22022 35048 22086 35112
rect 22022 34968 22086 35032
rect 22022 34888 22086 34952
rect 22022 34808 22086 34872
rect 22022 34728 22086 34792
rect 28341 40808 28405 40872
rect 28341 40728 28405 40792
rect 28341 40648 28405 40712
rect 28341 40568 28405 40632
rect 28341 40488 28405 40552
rect 28341 40408 28405 40472
rect 28341 40328 28405 40392
rect 28341 40248 28405 40312
rect 28341 40168 28405 40232
rect 28341 40088 28405 40152
rect 28341 40008 28405 40072
rect 28341 39928 28405 39992
rect 28341 39848 28405 39912
rect 28341 39768 28405 39832
rect 28341 39688 28405 39752
rect 28341 39608 28405 39672
rect 28341 39528 28405 39592
rect 28341 39448 28405 39512
rect 28341 39368 28405 39432
rect 28341 39288 28405 39352
rect 28341 39208 28405 39272
rect 28341 39128 28405 39192
rect 28341 39048 28405 39112
rect 28341 38968 28405 39032
rect 28341 38888 28405 38952
rect 28341 38808 28405 38872
rect 28341 38728 28405 38792
rect 28341 38648 28405 38712
rect 28341 38568 28405 38632
rect 28341 38488 28405 38552
rect 28341 38408 28405 38472
rect 28341 38328 28405 38392
rect 28341 38248 28405 38312
rect 28341 38168 28405 38232
rect 28341 38088 28405 38152
rect 28341 38008 28405 38072
rect 28341 37928 28405 37992
rect 28341 37848 28405 37912
rect 28341 37768 28405 37832
rect 28341 37688 28405 37752
rect 28341 37608 28405 37672
rect 28341 37528 28405 37592
rect 28341 37448 28405 37512
rect 28341 37368 28405 37432
rect 28341 37288 28405 37352
rect 28341 37208 28405 37272
rect 28341 37128 28405 37192
rect 28341 37048 28405 37112
rect 28341 36968 28405 37032
rect 28341 36888 28405 36952
rect 28341 36808 28405 36872
rect 28341 36728 28405 36792
rect 28341 36648 28405 36712
rect 28341 36568 28405 36632
rect 28341 36488 28405 36552
rect 28341 36408 28405 36472
rect 28341 36328 28405 36392
rect 28341 36248 28405 36312
rect 28341 36168 28405 36232
rect 28341 36088 28405 36152
rect 28341 36008 28405 36072
rect 28341 35928 28405 35992
rect 28341 35848 28405 35912
rect 28341 35768 28405 35832
rect 28341 35688 28405 35752
rect 28341 35608 28405 35672
rect 28341 35528 28405 35592
rect 28341 35448 28405 35512
rect 28341 35368 28405 35432
rect 28341 35288 28405 35352
rect 28341 35208 28405 35272
rect 28341 35128 28405 35192
rect 28341 35048 28405 35112
rect 28341 34968 28405 35032
rect 28341 34888 28405 34952
rect 28341 34808 28405 34872
rect 28341 34728 28405 34792
rect 34660 40808 34724 40872
rect 34660 40728 34724 40792
rect 34660 40648 34724 40712
rect 34660 40568 34724 40632
rect 34660 40488 34724 40552
rect 34660 40408 34724 40472
rect 34660 40328 34724 40392
rect 34660 40248 34724 40312
rect 34660 40168 34724 40232
rect 34660 40088 34724 40152
rect 34660 40008 34724 40072
rect 34660 39928 34724 39992
rect 34660 39848 34724 39912
rect 34660 39768 34724 39832
rect 34660 39688 34724 39752
rect 34660 39608 34724 39672
rect 34660 39528 34724 39592
rect 34660 39448 34724 39512
rect 34660 39368 34724 39432
rect 34660 39288 34724 39352
rect 34660 39208 34724 39272
rect 34660 39128 34724 39192
rect 34660 39048 34724 39112
rect 34660 38968 34724 39032
rect 34660 38888 34724 38952
rect 34660 38808 34724 38872
rect 34660 38728 34724 38792
rect 34660 38648 34724 38712
rect 34660 38568 34724 38632
rect 34660 38488 34724 38552
rect 34660 38408 34724 38472
rect 34660 38328 34724 38392
rect 34660 38248 34724 38312
rect 34660 38168 34724 38232
rect 34660 38088 34724 38152
rect 34660 38008 34724 38072
rect 34660 37928 34724 37992
rect 34660 37848 34724 37912
rect 34660 37768 34724 37832
rect 34660 37688 34724 37752
rect 34660 37608 34724 37672
rect 34660 37528 34724 37592
rect 34660 37448 34724 37512
rect 34660 37368 34724 37432
rect 34660 37288 34724 37352
rect 34660 37208 34724 37272
rect 34660 37128 34724 37192
rect 34660 37048 34724 37112
rect 34660 36968 34724 37032
rect 34660 36888 34724 36952
rect 34660 36808 34724 36872
rect 34660 36728 34724 36792
rect 34660 36648 34724 36712
rect 34660 36568 34724 36632
rect 34660 36488 34724 36552
rect 34660 36408 34724 36472
rect 34660 36328 34724 36392
rect 34660 36248 34724 36312
rect 34660 36168 34724 36232
rect 34660 36088 34724 36152
rect 34660 36008 34724 36072
rect 34660 35928 34724 35992
rect 34660 35848 34724 35912
rect 34660 35768 34724 35832
rect 34660 35688 34724 35752
rect 34660 35608 34724 35672
rect 34660 35528 34724 35592
rect 34660 35448 34724 35512
rect 34660 35368 34724 35432
rect 34660 35288 34724 35352
rect 34660 35208 34724 35272
rect 34660 35128 34724 35192
rect 34660 35048 34724 35112
rect 34660 34968 34724 35032
rect 34660 34888 34724 34952
rect 34660 34808 34724 34872
rect 34660 34728 34724 34792
rect 40979 40808 41043 40872
rect 40979 40728 41043 40792
rect 40979 40648 41043 40712
rect 40979 40568 41043 40632
rect 40979 40488 41043 40552
rect 40979 40408 41043 40472
rect 40979 40328 41043 40392
rect 40979 40248 41043 40312
rect 40979 40168 41043 40232
rect 40979 40088 41043 40152
rect 40979 40008 41043 40072
rect 40979 39928 41043 39992
rect 40979 39848 41043 39912
rect 40979 39768 41043 39832
rect 40979 39688 41043 39752
rect 40979 39608 41043 39672
rect 40979 39528 41043 39592
rect 40979 39448 41043 39512
rect 40979 39368 41043 39432
rect 40979 39288 41043 39352
rect 40979 39208 41043 39272
rect 40979 39128 41043 39192
rect 40979 39048 41043 39112
rect 40979 38968 41043 39032
rect 40979 38888 41043 38952
rect 40979 38808 41043 38872
rect 40979 38728 41043 38792
rect 40979 38648 41043 38712
rect 40979 38568 41043 38632
rect 40979 38488 41043 38552
rect 40979 38408 41043 38472
rect 40979 38328 41043 38392
rect 40979 38248 41043 38312
rect 40979 38168 41043 38232
rect 40979 38088 41043 38152
rect 40979 38008 41043 38072
rect 40979 37928 41043 37992
rect 40979 37848 41043 37912
rect 40979 37768 41043 37832
rect 40979 37688 41043 37752
rect 40979 37608 41043 37672
rect 40979 37528 41043 37592
rect 40979 37448 41043 37512
rect 40979 37368 41043 37432
rect 40979 37288 41043 37352
rect 40979 37208 41043 37272
rect 40979 37128 41043 37192
rect 40979 37048 41043 37112
rect 40979 36968 41043 37032
rect 40979 36888 41043 36952
rect 40979 36808 41043 36872
rect 40979 36728 41043 36792
rect 40979 36648 41043 36712
rect 40979 36568 41043 36632
rect 40979 36488 41043 36552
rect 40979 36408 41043 36472
rect 40979 36328 41043 36392
rect 40979 36248 41043 36312
rect 40979 36168 41043 36232
rect 40979 36088 41043 36152
rect 40979 36008 41043 36072
rect 40979 35928 41043 35992
rect 40979 35848 41043 35912
rect 40979 35768 41043 35832
rect 40979 35688 41043 35752
rect 40979 35608 41043 35672
rect 40979 35528 41043 35592
rect 40979 35448 41043 35512
rect 40979 35368 41043 35432
rect 40979 35288 41043 35352
rect 40979 35208 41043 35272
rect 40979 35128 41043 35192
rect 40979 35048 41043 35112
rect 40979 34968 41043 35032
rect 40979 34888 41043 34952
rect 40979 34808 41043 34872
rect 40979 34728 41043 34792
rect 47298 40808 47362 40872
rect 47298 40728 47362 40792
rect 47298 40648 47362 40712
rect 47298 40568 47362 40632
rect 47298 40488 47362 40552
rect 47298 40408 47362 40472
rect 47298 40328 47362 40392
rect 47298 40248 47362 40312
rect 47298 40168 47362 40232
rect 47298 40088 47362 40152
rect 47298 40008 47362 40072
rect 47298 39928 47362 39992
rect 47298 39848 47362 39912
rect 47298 39768 47362 39832
rect 47298 39688 47362 39752
rect 47298 39608 47362 39672
rect 47298 39528 47362 39592
rect 47298 39448 47362 39512
rect 47298 39368 47362 39432
rect 47298 39288 47362 39352
rect 47298 39208 47362 39272
rect 47298 39128 47362 39192
rect 47298 39048 47362 39112
rect 47298 38968 47362 39032
rect 47298 38888 47362 38952
rect 47298 38808 47362 38872
rect 47298 38728 47362 38792
rect 47298 38648 47362 38712
rect 47298 38568 47362 38632
rect 47298 38488 47362 38552
rect 47298 38408 47362 38472
rect 47298 38328 47362 38392
rect 47298 38248 47362 38312
rect 47298 38168 47362 38232
rect 47298 38088 47362 38152
rect 47298 38008 47362 38072
rect 47298 37928 47362 37992
rect 47298 37848 47362 37912
rect 47298 37768 47362 37832
rect 47298 37688 47362 37752
rect 47298 37608 47362 37672
rect 47298 37528 47362 37592
rect 47298 37448 47362 37512
rect 47298 37368 47362 37432
rect 47298 37288 47362 37352
rect 47298 37208 47362 37272
rect 47298 37128 47362 37192
rect 47298 37048 47362 37112
rect 47298 36968 47362 37032
rect 47298 36888 47362 36952
rect 47298 36808 47362 36872
rect 47298 36728 47362 36792
rect 47298 36648 47362 36712
rect 47298 36568 47362 36632
rect 47298 36488 47362 36552
rect 47298 36408 47362 36472
rect 47298 36328 47362 36392
rect 47298 36248 47362 36312
rect 47298 36168 47362 36232
rect 47298 36088 47362 36152
rect 47298 36008 47362 36072
rect 47298 35928 47362 35992
rect 47298 35848 47362 35912
rect 47298 35768 47362 35832
rect 47298 35688 47362 35752
rect 47298 35608 47362 35672
rect 47298 35528 47362 35592
rect 47298 35448 47362 35512
rect 47298 35368 47362 35432
rect 47298 35288 47362 35352
rect 47298 35208 47362 35272
rect 47298 35128 47362 35192
rect 47298 35048 47362 35112
rect 47298 34968 47362 35032
rect 47298 34888 47362 34952
rect 47298 34808 47362 34872
rect 47298 34728 47362 34792
rect -41168 34508 -41104 34572
rect -41168 34428 -41104 34492
rect -41168 34348 -41104 34412
rect -41168 34268 -41104 34332
rect -41168 34188 -41104 34252
rect -41168 34108 -41104 34172
rect -41168 34028 -41104 34092
rect -41168 33948 -41104 34012
rect -41168 33868 -41104 33932
rect -41168 33788 -41104 33852
rect -41168 33708 -41104 33772
rect -41168 33628 -41104 33692
rect -41168 33548 -41104 33612
rect -41168 33468 -41104 33532
rect -41168 33388 -41104 33452
rect -41168 33308 -41104 33372
rect -41168 33228 -41104 33292
rect -41168 33148 -41104 33212
rect -41168 33068 -41104 33132
rect -41168 32988 -41104 33052
rect -41168 32908 -41104 32972
rect -41168 32828 -41104 32892
rect -41168 32748 -41104 32812
rect -41168 32668 -41104 32732
rect -41168 32588 -41104 32652
rect -41168 32508 -41104 32572
rect -41168 32428 -41104 32492
rect -41168 32348 -41104 32412
rect -41168 32268 -41104 32332
rect -41168 32188 -41104 32252
rect -41168 32108 -41104 32172
rect -41168 32028 -41104 32092
rect -41168 31948 -41104 32012
rect -41168 31868 -41104 31932
rect -41168 31788 -41104 31852
rect -41168 31708 -41104 31772
rect -41168 31628 -41104 31692
rect -41168 31548 -41104 31612
rect -41168 31468 -41104 31532
rect -41168 31388 -41104 31452
rect -41168 31308 -41104 31372
rect -41168 31228 -41104 31292
rect -41168 31148 -41104 31212
rect -41168 31068 -41104 31132
rect -41168 30988 -41104 31052
rect -41168 30908 -41104 30972
rect -41168 30828 -41104 30892
rect -41168 30748 -41104 30812
rect -41168 30668 -41104 30732
rect -41168 30588 -41104 30652
rect -41168 30508 -41104 30572
rect -41168 30428 -41104 30492
rect -41168 30348 -41104 30412
rect -41168 30268 -41104 30332
rect -41168 30188 -41104 30252
rect -41168 30108 -41104 30172
rect -41168 30028 -41104 30092
rect -41168 29948 -41104 30012
rect -41168 29868 -41104 29932
rect -41168 29788 -41104 29852
rect -41168 29708 -41104 29772
rect -41168 29628 -41104 29692
rect -41168 29548 -41104 29612
rect -41168 29468 -41104 29532
rect -41168 29388 -41104 29452
rect -41168 29308 -41104 29372
rect -41168 29228 -41104 29292
rect -41168 29148 -41104 29212
rect -41168 29068 -41104 29132
rect -41168 28988 -41104 29052
rect -41168 28908 -41104 28972
rect -41168 28828 -41104 28892
rect -41168 28748 -41104 28812
rect -41168 28668 -41104 28732
rect -41168 28588 -41104 28652
rect -41168 28508 -41104 28572
rect -41168 28428 -41104 28492
rect -34849 34508 -34785 34572
rect -34849 34428 -34785 34492
rect -34849 34348 -34785 34412
rect -34849 34268 -34785 34332
rect -34849 34188 -34785 34252
rect -34849 34108 -34785 34172
rect -34849 34028 -34785 34092
rect -34849 33948 -34785 34012
rect -34849 33868 -34785 33932
rect -34849 33788 -34785 33852
rect -34849 33708 -34785 33772
rect -34849 33628 -34785 33692
rect -34849 33548 -34785 33612
rect -34849 33468 -34785 33532
rect -34849 33388 -34785 33452
rect -34849 33308 -34785 33372
rect -34849 33228 -34785 33292
rect -34849 33148 -34785 33212
rect -34849 33068 -34785 33132
rect -34849 32988 -34785 33052
rect -34849 32908 -34785 32972
rect -34849 32828 -34785 32892
rect -34849 32748 -34785 32812
rect -34849 32668 -34785 32732
rect -34849 32588 -34785 32652
rect -34849 32508 -34785 32572
rect -34849 32428 -34785 32492
rect -34849 32348 -34785 32412
rect -34849 32268 -34785 32332
rect -34849 32188 -34785 32252
rect -34849 32108 -34785 32172
rect -34849 32028 -34785 32092
rect -34849 31948 -34785 32012
rect -34849 31868 -34785 31932
rect -34849 31788 -34785 31852
rect -34849 31708 -34785 31772
rect -34849 31628 -34785 31692
rect -34849 31548 -34785 31612
rect -34849 31468 -34785 31532
rect -34849 31388 -34785 31452
rect -34849 31308 -34785 31372
rect -34849 31228 -34785 31292
rect -34849 31148 -34785 31212
rect -34849 31068 -34785 31132
rect -34849 30988 -34785 31052
rect -34849 30908 -34785 30972
rect -34849 30828 -34785 30892
rect -34849 30748 -34785 30812
rect -34849 30668 -34785 30732
rect -34849 30588 -34785 30652
rect -34849 30508 -34785 30572
rect -34849 30428 -34785 30492
rect -34849 30348 -34785 30412
rect -34849 30268 -34785 30332
rect -34849 30188 -34785 30252
rect -34849 30108 -34785 30172
rect -34849 30028 -34785 30092
rect -34849 29948 -34785 30012
rect -34849 29868 -34785 29932
rect -34849 29788 -34785 29852
rect -34849 29708 -34785 29772
rect -34849 29628 -34785 29692
rect -34849 29548 -34785 29612
rect -34849 29468 -34785 29532
rect -34849 29388 -34785 29452
rect -34849 29308 -34785 29372
rect -34849 29228 -34785 29292
rect -34849 29148 -34785 29212
rect -34849 29068 -34785 29132
rect -34849 28988 -34785 29052
rect -34849 28908 -34785 28972
rect -34849 28828 -34785 28892
rect -34849 28748 -34785 28812
rect -34849 28668 -34785 28732
rect -34849 28588 -34785 28652
rect -34849 28508 -34785 28572
rect -34849 28428 -34785 28492
rect -28530 34508 -28466 34572
rect -28530 34428 -28466 34492
rect -28530 34348 -28466 34412
rect -28530 34268 -28466 34332
rect -28530 34188 -28466 34252
rect -28530 34108 -28466 34172
rect -28530 34028 -28466 34092
rect -28530 33948 -28466 34012
rect -28530 33868 -28466 33932
rect -28530 33788 -28466 33852
rect -28530 33708 -28466 33772
rect -28530 33628 -28466 33692
rect -28530 33548 -28466 33612
rect -28530 33468 -28466 33532
rect -28530 33388 -28466 33452
rect -28530 33308 -28466 33372
rect -28530 33228 -28466 33292
rect -28530 33148 -28466 33212
rect -28530 33068 -28466 33132
rect -28530 32988 -28466 33052
rect -28530 32908 -28466 32972
rect -28530 32828 -28466 32892
rect -28530 32748 -28466 32812
rect -28530 32668 -28466 32732
rect -28530 32588 -28466 32652
rect -28530 32508 -28466 32572
rect -28530 32428 -28466 32492
rect -28530 32348 -28466 32412
rect -28530 32268 -28466 32332
rect -28530 32188 -28466 32252
rect -28530 32108 -28466 32172
rect -28530 32028 -28466 32092
rect -28530 31948 -28466 32012
rect -28530 31868 -28466 31932
rect -28530 31788 -28466 31852
rect -28530 31708 -28466 31772
rect -28530 31628 -28466 31692
rect -28530 31548 -28466 31612
rect -28530 31468 -28466 31532
rect -28530 31388 -28466 31452
rect -28530 31308 -28466 31372
rect -28530 31228 -28466 31292
rect -28530 31148 -28466 31212
rect -28530 31068 -28466 31132
rect -28530 30988 -28466 31052
rect -28530 30908 -28466 30972
rect -28530 30828 -28466 30892
rect -28530 30748 -28466 30812
rect -28530 30668 -28466 30732
rect -28530 30588 -28466 30652
rect -28530 30508 -28466 30572
rect -28530 30428 -28466 30492
rect -28530 30348 -28466 30412
rect -28530 30268 -28466 30332
rect -28530 30188 -28466 30252
rect -28530 30108 -28466 30172
rect -28530 30028 -28466 30092
rect -28530 29948 -28466 30012
rect -28530 29868 -28466 29932
rect -28530 29788 -28466 29852
rect -28530 29708 -28466 29772
rect -28530 29628 -28466 29692
rect -28530 29548 -28466 29612
rect -28530 29468 -28466 29532
rect -28530 29388 -28466 29452
rect -28530 29308 -28466 29372
rect -28530 29228 -28466 29292
rect -28530 29148 -28466 29212
rect -28530 29068 -28466 29132
rect -28530 28988 -28466 29052
rect -28530 28908 -28466 28972
rect -28530 28828 -28466 28892
rect -28530 28748 -28466 28812
rect -28530 28668 -28466 28732
rect -28530 28588 -28466 28652
rect -28530 28508 -28466 28572
rect -28530 28428 -28466 28492
rect -22211 34508 -22147 34572
rect -22211 34428 -22147 34492
rect -22211 34348 -22147 34412
rect -22211 34268 -22147 34332
rect -22211 34188 -22147 34252
rect -22211 34108 -22147 34172
rect -22211 34028 -22147 34092
rect -22211 33948 -22147 34012
rect -22211 33868 -22147 33932
rect -22211 33788 -22147 33852
rect -22211 33708 -22147 33772
rect -22211 33628 -22147 33692
rect -22211 33548 -22147 33612
rect -22211 33468 -22147 33532
rect -22211 33388 -22147 33452
rect -22211 33308 -22147 33372
rect -22211 33228 -22147 33292
rect -22211 33148 -22147 33212
rect -22211 33068 -22147 33132
rect -22211 32988 -22147 33052
rect -22211 32908 -22147 32972
rect -22211 32828 -22147 32892
rect -22211 32748 -22147 32812
rect -22211 32668 -22147 32732
rect -22211 32588 -22147 32652
rect -22211 32508 -22147 32572
rect -22211 32428 -22147 32492
rect -22211 32348 -22147 32412
rect -22211 32268 -22147 32332
rect -22211 32188 -22147 32252
rect -22211 32108 -22147 32172
rect -22211 32028 -22147 32092
rect -22211 31948 -22147 32012
rect -22211 31868 -22147 31932
rect -22211 31788 -22147 31852
rect -22211 31708 -22147 31772
rect -22211 31628 -22147 31692
rect -22211 31548 -22147 31612
rect -22211 31468 -22147 31532
rect -22211 31388 -22147 31452
rect -22211 31308 -22147 31372
rect -22211 31228 -22147 31292
rect -22211 31148 -22147 31212
rect -22211 31068 -22147 31132
rect -22211 30988 -22147 31052
rect -22211 30908 -22147 30972
rect -22211 30828 -22147 30892
rect -22211 30748 -22147 30812
rect -22211 30668 -22147 30732
rect -22211 30588 -22147 30652
rect -22211 30508 -22147 30572
rect -22211 30428 -22147 30492
rect -22211 30348 -22147 30412
rect -22211 30268 -22147 30332
rect -22211 30188 -22147 30252
rect -22211 30108 -22147 30172
rect -22211 30028 -22147 30092
rect -22211 29948 -22147 30012
rect -22211 29868 -22147 29932
rect -22211 29788 -22147 29852
rect -22211 29708 -22147 29772
rect -22211 29628 -22147 29692
rect -22211 29548 -22147 29612
rect -22211 29468 -22147 29532
rect -22211 29388 -22147 29452
rect -22211 29308 -22147 29372
rect -22211 29228 -22147 29292
rect -22211 29148 -22147 29212
rect -22211 29068 -22147 29132
rect -22211 28988 -22147 29052
rect -22211 28908 -22147 28972
rect -22211 28828 -22147 28892
rect -22211 28748 -22147 28812
rect -22211 28668 -22147 28732
rect -22211 28588 -22147 28652
rect -22211 28508 -22147 28572
rect -22211 28428 -22147 28492
rect -15892 34508 -15828 34572
rect -15892 34428 -15828 34492
rect -15892 34348 -15828 34412
rect -15892 34268 -15828 34332
rect -15892 34188 -15828 34252
rect -15892 34108 -15828 34172
rect -15892 34028 -15828 34092
rect -15892 33948 -15828 34012
rect -15892 33868 -15828 33932
rect -15892 33788 -15828 33852
rect -15892 33708 -15828 33772
rect -15892 33628 -15828 33692
rect -15892 33548 -15828 33612
rect -15892 33468 -15828 33532
rect -15892 33388 -15828 33452
rect -15892 33308 -15828 33372
rect -15892 33228 -15828 33292
rect -15892 33148 -15828 33212
rect -15892 33068 -15828 33132
rect -15892 32988 -15828 33052
rect -15892 32908 -15828 32972
rect -15892 32828 -15828 32892
rect -15892 32748 -15828 32812
rect -15892 32668 -15828 32732
rect -15892 32588 -15828 32652
rect -15892 32508 -15828 32572
rect -15892 32428 -15828 32492
rect -15892 32348 -15828 32412
rect -15892 32268 -15828 32332
rect -15892 32188 -15828 32252
rect -15892 32108 -15828 32172
rect -15892 32028 -15828 32092
rect -15892 31948 -15828 32012
rect -15892 31868 -15828 31932
rect -15892 31788 -15828 31852
rect -15892 31708 -15828 31772
rect -15892 31628 -15828 31692
rect -15892 31548 -15828 31612
rect -15892 31468 -15828 31532
rect -15892 31388 -15828 31452
rect -15892 31308 -15828 31372
rect -15892 31228 -15828 31292
rect -15892 31148 -15828 31212
rect -15892 31068 -15828 31132
rect -15892 30988 -15828 31052
rect -15892 30908 -15828 30972
rect -15892 30828 -15828 30892
rect -15892 30748 -15828 30812
rect -15892 30668 -15828 30732
rect -15892 30588 -15828 30652
rect -15892 30508 -15828 30572
rect -15892 30428 -15828 30492
rect -15892 30348 -15828 30412
rect -15892 30268 -15828 30332
rect -15892 30188 -15828 30252
rect -15892 30108 -15828 30172
rect -15892 30028 -15828 30092
rect -15892 29948 -15828 30012
rect -15892 29868 -15828 29932
rect -15892 29788 -15828 29852
rect -15892 29708 -15828 29772
rect -15892 29628 -15828 29692
rect -15892 29548 -15828 29612
rect -15892 29468 -15828 29532
rect -15892 29388 -15828 29452
rect -15892 29308 -15828 29372
rect -15892 29228 -15828 29292
rect -15892 29148 -15828 29212
rect -15892 29068 -15828 29132
rect -15892 28988 -15828 29052
rect -15892 28908 -15828 28972
rect -15892 28828 -15828 28892
rect -15892 28748 -15828 28812
rect -15892 28668 -15828 28732
rect -15892 28588 -15828 28652
rect -15892 28508 -15828 28572
rect -15892 28428 -15828 28492
rect -9573 34508 -9509 34572
rect -9573 34428 -9509 34492
rect -9573 34348 -9509 34412
rect -9573 34268 -9509 34332
rect -9573 34188 -9509 34252
rect -9573 34108 -9509 34172
rect -9573 34028 -9509 34092
rect -9573 33948 -9509 34012
rect -9573 33868 -9509 33932
rect -9573 33788 -9509 33852
rect -9573 33708 -9509 33772
rect -9573 33628 -9509 33692
rect -9573 33548 -9509 33612
rect -9573 33468 -9509 33532
rect -9573 33388 -9509 33452
rect -9573 33308 -9509 33372
rect -9573 33228 -9509 33292
rect -9573 33148 -9509 33212
rect -9573 33068 -9509 33132
rect -9573 32988 -9509 33052
rect -9573 32908 -9509 32972
rect -9573 32828 -9509 32892
rect -9573 32748 -9509 32812
rect -9573 32668 -9509 32732
rect -9573 32588 -9509 32652
rect -9573 32508 -9509 32572
rect -9573 32428 -9509 32492
rect -9573 32348 -9509 32412
rect -9573 32268 -9509 32332
rect -9573 32188 -9509 32252
rect -9573 32108 -9509 32172
rect -9573 32028 -9509 32092
rect -9573 31948 -9509 32012
rect -9573 31868 -9509 31932
rect -9573 31788 -9509 31852
rect -9573 31708 -9509 31772
rect -9573 31628 -9509 31692
rect -9573 31548 -9509 31612
rect -9573 31468 -9509 31532
rect -9573 31388 -9509 31452
rect -9573 31308 -9509 31372
rect -9573 31228 -9509 31292
rect -9573 31148 -9509 31212
rect -9573 31068 -9509 31132
rect -9573 30988 -9509 31052
rect -9573 30908 -9509 30972
rect -9573 30828 -9509 30892
rect -9573 30748 -9509 30812
rect -9573 30668 -9509 30732
rect -9573 30588 -9509 30652
rect -9573 30508 -9509 30572
rect -9573 30428 -9509 30492
rect -9573 30348 -9509 30412
rect -9573 30268 -9509 30332
rect -9573 30188 -9509 30252
rect -9573 30108 -9509 30172
rect -9573 30028 -9509 30092
rect -9573 29948 -9509 30012
rect -9573 29868 -9509 29932
rect -9573 29788 -9509 29852
rect -9573 29708 -9509 29772
rect -9573 29628 -9509 29692
rect -9573 29548 -9509 29612
rect -9573 29468 -9509 29532
rect -9573 29388 -9509 29452
rect -9573 29308 -9509 29372
rect -9573 29228 -9509 29292
rect -9573 29148 -9509 29212
rect -9573 29068 -9509 29132
rect -9573 28988 -9509 29052
rect -9573 28908 -9509 28972
rect -9573 28828 -9509 28892
rect -9573 28748 -9509 28812
rect -9573 28668 -9509 28732
rect -9573 28588 -9509 28652
rect -9573 28508 -9509 28572
rect -9573 28428 -9509 28492
rect -3254 34508 -3190 34572
rect -3254 34428 -3190 34492
rect -3254 34348 -3190 34412
rect -3254 34268 -3190 34332
rect -3254 34188 -3190 34252
rect -3254 34108 -3190 34172
rect -3254 34028 -3190 34092
rect -3254 33948 -3190 34012
rect -3254 33868 -3190 33932
rect -3254 33788 -3190 33852
rect -3254 33708 -3190 33772
rect -3254 33628 -3190 33692
rect -3254 33548 -3190 33612
rect -3254 33468 -3190 33532
rect -3254 33388 -3190 33452
rect -3254 33308 -3190 33372
rect -3254 33228 -3190 33292
rect -3254 33148 -3190 33212
rect -3254 33068 -3190 33132
rect -3254 32988 -3190 33052
rect -3254 32908 -3190 32972
rect -3254 32828 -3190 32892
rect -3254 32748 -3190 32812
rect -3254 32668 -3190 32732
rect -3254 32588 -3190 32652
rect -3254 32508 -3190 32572
rect -3254 32428 -3190 32492
rect -3254 32348 -3190 32412
rect -3254 32268 -3190 32332
rect -3254 32188 -3190 32252
rect -3254 32108 -3190 32172
rect -3254 32028 -3190 32092
rect -3254 31948 -3190 32012
rect -3254 31868 -3190 31932
rect -3254 31788 -3190 31852
rect -3254 31708 -3190 31772
rect -3254 31628 -3190 31692
rect -3254 31548 -3190 31612
rect -3254 31468 -3190 31532
rect -3254 31388 -3190 31452
rect -3254 31308 -3190 31372
rect -3254 31228 -3190 31292
rect -3254 31148 -3190 31212
rect -3254 31068 -3190 31132
rect -3254 30988 -3190 31052
rect -3254 30908 -3190 30972
rect -3254 30828 -3190 30892
rect -3254 30748 -3190 30812
rect -3254 30668 -3190 30732
rect -3254 30588 -3190 30652
rect -3254 30508 -3190 30572
rect -3254 30428 -3190 30492
rect -3254 30348 -3190 30412
rect -3254 30268 -3190 30332
rect -3254 30188 -3190 30252
rect -3254 30108 -3190 30172
rect -3254 30028 -3190 30092
rect -3254 29948 -3190 30012
rect -3254 29868 -3190 29932
rect -3254 29788 -3190 29852
rect -3254 29708 -3190 29772
rect -3254 29628 -3190 29692
rect -3254 29548 -3190 29612
rect -3254 29468 -3190 29532
rect -3254 29388 -3190 29452
rect -3254 29308 -3190 29372
rect -3254 29228 -3190 29292
rect -3254 29148 -3190 29212
rect -3254 29068 -3190 29132
rect -3254 28988 -3190 29052
rect -3254 28908 -3190 28972
rect -3254 28828 -3190 28892
rect -3254 28748 -3190 28812
rect -3254 28668 -3190 28732
rect -3254 28588 -3190 28652
rect -3254 28508 -3190 28572
rect -3254 28428 -3190 28492
rect 3065 34508 3129 34572
rect 3065 34428 3129 34492
rect 3065 34348 3129 34412
rect 3065 34268 3129 34332
rect 3065 34188 3129 34252
rect 3065 34108 3129 34172
rect 3065 34028 3129 34092
rect 3065 33948 3129 34012
rect 3065 33868 3129 33932
rect 3065 33788 3129 33852
rect 3065 33708 3129 33772
rect 3065 33628 3129 33692
rect 3065 33548 3129 33612
rect 3065 33468 3129 33532
rect 3065 33388 3129 33452
rect 3065 33308 3129 33372
rect 3065 33228 3129 33292
rect 3065 33148 3129 33212
rect 3065 33068 3129 33132
rect 3065 32988 3129 33052
rect 3065 32908 3129 32972
rect 3065 32828 3129 32892
rect 3065 32748 3129 32812
rect 3065 32668 3129 32732
rect 3065 32588 3129 32652
rect 3065 32508 3129 32572
rect 3065 32428 3129 32492
rect 3065 32348 3129 32412
rect 3065 32268 3129 32332
rect 3065 32188 3129 32252
rect 3065 32108 3129 32172
rect 3065 32028 3129 32092
rect 3065 31948 3129 32012
rect 3065 31868 3129 31932
rect 3065 31788 3129 31852
rect 3065 31708 3129 31772
rect 3065 31628 3129 31692
rect 3065 31548 3129 31612
rect 3065 31468 3129 31532
rect 3065 31388 3129 31452
rect 3065 31308 3129 31372
rect 3065 31228 3129 31292
rect 3065 31148 3129 31212
rect 3065 31068 3129 31132
rect 3065 30988 3129 31052
rect 3065 30908 3129 30972
rect 3065 30828 3129 30892
rect 3065 30748 3129 30812
rect 3065 30668 3129 30732
rect 3065 30588 3129 30652
rect 3065 30508 3129 30572
rect 3065 30428 3129 30492
rect 3065 30348 3129 30412
rect 3065 30268 3129 30332
rect 3065 30188 3129 30252
rect 3065 30108 3129 30172
rect 3065 30028 3129 30092
rect 3065 29948 3129 30012
rect 3065 29868 3129 29932
rect 3065 29788 3129 29852
rect 3065 29708 3129 29772
rect 3065 29628 3129 29692
rect 3065 29548 3129 29612
rect 3065 29468 3129 29532
rect 3065 29388 3129 29452
rect 3065 29308 3129 29372
rect 3065 29228 3129 29292
rect 3065 29148 3129 29212
rect 3065 29068 3129 29132
rect 3065 28988 3129 29052
rect 3065 28908 3129 28972
rect 3065 28828 3129 28892
rect 3065 28748 3129 28812
rect 3065 28668 3129 28732
rect 3065 28588 3129 28652
rect 3065 28508 3129 28572
rect 3065 28428 3129 28492
rect 9384 34508 9448 34572
rect 9384 34428 9448 34492
rect 9384 34348 9448 34412
rect 9384 34268 9448 34332
rect 9384 34188 9448 34252
rect 9384 34108 9448 34172
rect 9384 34028 9448 34092
rect 9384 33948 9448 34012
rect 9384 33868 9448 33932
rect 9384 33788 9448 33852
rect 9384 33708 9448 33772
rect 9384 33628 9448 33692
rect 9384 33548 9448 33612
rect 9384 33468 9448 33532
rect 9384 33388 9448 33452
rect 9384 33308 9448 33372
rect 9384 33228 9448 33292
rect 9384 33148 9448 33212
rect 9384 33068 9448 33132
rect 9384 32988 9448 33052
rect 9384 32908 9448 32972
rect 9384 32828 9448 32892
rect 9384 32748 9448 32812
rect 9384 32668 9448 32732
rect 9384 32588 9448 32652
rect 9384 32508 9448 32572
rect 9384 32428 9448 32492
rect 9384 32348 9448 32412
rect 9384 32268 9448 32332
rect 9384 32188 9448 32252
rect 9384 32108 9448 32172
rect 9384 32028 9448 32092
rect 9384 31948 9448 32012
rect 9384 31868 9448 31932
rect 9384 31788 9448 31852
rect 9384 31708 9448 31772
rect 9384 31628 9448 31692
rect 9384 31548 9448 31612
rect 9384 31468 9448 31532
rect 9384 31388 9448 31452
rect 9384 31308 9448 31372
rect 9384 31228 9448 31292
rect 9384 31148 9448 31212
rect 9384 31068 9448 31132
rect 9384 30988 9448 31052
rect 9384 30908 9448 30972
rect 9384 30828 9448 30892
rect 9384 30748 9448 30812
rect 9384 30668 9448 30732
rect 9384 30588 9448 30652
rect 9384 30508 9448 30572
rect 9384 30428 9448 30492
rect 9384 30348 9448 30412
rect 9384 30268 9448 30332
rect 9384 30188 9448 30252
rect 9384 30108 9448 30172
rect 9384 30028 9448 30092
rect 9384 29948 9448 30012
rect 9384 29868 9448 29932
rect 9384 29788 9448 29852
rect 9384 29708 9448 29772
rect 9384 29628 9448 29692
rect 9384 29548 9448 29612
rect 9384 29468 9448 29532
rect 9384 29388 9448 29452
rect 9384 29308 9448 29372
rect 9384 29228 9448 29292
rect 9384 29148 9448 29212
rect 9384 29068 9448 29132
rect 9384 28988 9448 29052
rect 9384 28908 9448 28972
rect 9384 28828 9448 28892
rect 9384 28748 9448 28812
rect 9384 28668 9448 28732
rect 9384 28588 9448 28652
rect 9384 28508 9448 28572
rect 9384 28428 9448 28492
rect 15703 34508 15767 34572
rect 15703 34428 15767 34492
rect 15703 34348 15767 34412
rect 15703 34268 15767 34332
rect 15703 34188 15767 34252
rect 15703 34108 15767 34172
rect 15703 34028 15767 34092
rect 15703 33948 15767 34012
rect 15703 33868 15767 33932
rect 15703 33788 15767 33852
rect 15703 33708 15767 33772
rect 15703 33628 15767 33692
rect 15703 33548 15767 33612
rect 15703 33468 15767 33532
rect 15703 33388 15767 33452
rect 15703 33308 15767 33372
rect 15703 33228 15767 33292
rect 15703 33148 15767 33212
rect 15703 33068 15767 33132
rect 15703 32988 15767 33052
rect 15703 32908 15767 32972
rect 15703 32828 15767 32892
rect 15703 32748 15767 32812
rect 15703 32668 15767 32732
rect 15703 32588 15767 32652
rect 15703 32508 15767 32572
rect 15703 32428 15767 32492
rect 15703 32348 15767 32412
rect 15703 32268 15767 32332
rect 15703 32188 15767 32252
rect 15703 32108 15767 32172
rect 15703 32028 15767 32092
rect 15703 31948 15767 32012
rect 15703 31868 15767 31932
rect 15703 31788 15767 31852
rect 15703 31708 15767 31772
rect 15703 31628 15767 31692
rect 15703 31548 15767 31612
rect 15703 31468 15767 31532
rect 15703 31388 15767 31452
rect 15703 31308 15767 31372
rect 15703 31228 15767 31292
rect 15703 31148 15767 31212
rect 15703 31068 15767 31132
rect 15703 30988 15767 31052
rect 15703 30908 15767 30972
rect 15703 30828 15767 30892
rect 15703 30748 15767 30812
rect 15703 30668 15767 30732
rect 15703 30588 15767 30652
rect 15703 30508 15767 30572
rect 15703 30428 15767 30492
rect 15703 30348 15767 30412
rect 15703 30268 15767 30332
rect 15703 30188 15767 30252
rect 15703 30108 15767 30172
rect 15703 30028 15767 30092
rect 15703 29948 15767 30012
rect 15703 29868 15767 29932
rect 15703 29788 15767 29852
rect 15703 29708 15767 29772
rect 15703 29628 15767 29692
rect 15703 29548 15767 29612
rect 15703 29468 15767 29532
rect 15703 29388 15767 29452
rect 15703 29308 15767 29372
rect 15703 29228 15767 29292
rect 15703 29148 15767 29212
rect 15703 29068 15767 29132
rect 15703 28988 15767 29052
rect 15703 28908 15767 28972
rect 15703 28828 15767 28892
rect 15703 28748 15767 28812
rect 15703 28668 15767 28732
rect 15703 28588 15767 28652
rect 15703 28508 15767 28572
rect 15703 28428 15767 28492
rect 22022 34508 22086 34572
rect 22022 34428 22086 34492
rect 22022 34348 22086 34412
rect 22022 34268 22086 34332
rect 22022 34188 22086 34252
rect 22022 34108 22086 34172
rect 22022 34028 22086 34092
rect 22022 33948 22086 34012
rect 22022 33868 22086 33932
rect 22022 33788 22086 33852
rect 22022 33708 22086 33772
rect 22022 33628 22086 33692
rect 22022 33548 22086 33612
rect 22022 33468 22086 33532
rect 22022 33388 22086 33452
rect 22022 33308 22086 33372
rect 22022 33228 22086 33292
rect 22022 33148 22086 33212
rect 22022 33068 22086 33132
rect 22022 32988 22086 33052
rect 22022 32908 22086 32972
rect 22022 32828 22086 32892
rect 22022 32748 22086 32812
rect 22022 32668 22086 32732
rect 22022 32588 22086 32652
rect 22022 32508 22086 32572
rect 22022 32428 22086 32492
rect 22022 32348 22086 32412
rect 22022 32268 22086 32332
rect 22022 32188 22086 32252
rect 22022 32108 22086 32172
rect 22022 32028 22086 32092
rect 22022 31948 22086 32012
rect 22022 31868 22086 31932
rect 22022 31788 22086 31852
rect 22022 31708 22086 31772
rect 22022 31628 22086 31692
rect 22022 31548 22086 31612
rect 22022 31468 22086 31532
rect 22022 31388 22086 31452
rect 22022 31308 22086 31372
rect 22022 31228 22086 31292
rect 22022 31148 22086 31212
rect 22022 31068 22086 31132
rect 22022 30988 22086 31052
rect 22022 30908 22086 30972
rect 22022 30828 22086 30892
rect 22022 30748 22086 30812
rect 22022 30668 22086 30732
rect 22022 30588 22086 30652
rect 22022 30508 22086 30572
rect 22022 30428 22086 30492
rect 22022 30348 22086 30412
rect 22022 30268 22086 30332
rect 22022 30188 22086 30252
rect 22022 30108 22086 30172
rect 22022 30028 22086 30092
rect 22022 29948 22086 30012
rect 22022 29868 22086 29932
rect 22022 29788 22086 29852
rect 22022 29708 22086 29772
rect 22022 29628 22086 29692
rect 22022 29548 22086 29612
rect 22022 29468 22086 29532
rect 22022 29388 22086 29452
rect 22022 29308 22086 29372
rect 22022 29228 22086 29292
rect 22022 29148 22086 29212
rect 22022 29068 22086 29132
rect 22022 28988 22086 29052
rect 22022 28908 22086 28972
rect 22022 28828 22086 28892
rect 22022 28748 22086 28812
rect 22022 28668 22086 28732
rect 22022 28588 22086 28652
rect 22022 28508 22086 28572
rect 22022 28428 22086 28492
rect 28341 34508 28405 34572
rect 28341 34428 28405 34492
rect 28341 34348 28405 34412
rect 28341 34268 28405 34332
rect 28341 34188 28405 34252
rect 28341 34108 28405 34172
rect 28341 34028 28405 34092
rect 28341 33948 28405 34012
rect 28341 33868 28405 33932
rect 28341 33788 28405 33852
rect 28341 33708 28405 33772
rect 28341 33628 28405 33692
rect 28341 33548 28405 33612
rect 28341 33468 28405 33532
rect 28341 33388 28405 33452
rect 28341 33308 28405 33372
rect 28341 33228 28405 33292
rect 28341 33148 28405 33212
rect 28341 33068 28405 33132
rect 28341 32988 28405 33052
rect 28341 32908 28405 32972
rect 28341 32828 28405 32892
rect 28341 32748 28405 32812
rect 28341 32668 28405 32732
rect 28341 32588 28405 32652
rect 28341 32508 28405 32572
rect 28341 32428 28405 32492
rect 28341 32348 28405 32412
rect 28341 32268 28405 32332
rect 28341 32188 28405 32252
rect 28341 32108 28405 32172
rect 28341 32028 28405 32092
rect 28341 31948 28405 32012
rect 28341 31868 28405 31932
rect 28341 31788 28405 31852
rect 28341 31708 28405 31772
rect 28341 31628 28405 31692
rect 28341 31548 28405 31612
rect 28341 31468 28405 31532
rect 28341 31388 28405 31452
rect 28341 31308 28405 31372
rect 28341 31228 28405 31292
rect 28341 31148 28405 31212
rect 28341 31068 28405 31132
rect 28341 30988 28405 31052
rect 28341 30908 28405 30972
rect 28341 30828 28405 30892
rect 28341 30748 28405 30812
rect 28341 30668 28405 30732
rect 28341 30588 28405 30652
rect 28341 30508 28405 30572
rect 28341 30428 28405 30492
rect 28341 30348 28405 30412
rect 28341 30268 28405 30332
rect 28341 30188 28405 30252
rect 28341 30108 28405 30172
rect 28341 30028 28405 30092
rect 28341 29948 28405 30012
rect 28341 29868 28405 29932
rect 28341 29788 28405 29852
rect 28341 29708 28405 29772
rect 28341 29628 28405 29692
rect 28341 29548 28405 29612
rect 28341 29468 28405 29532
rect 28341 29388 28405 29452
rect 28341 29308 28405 29372
rect 28341 29228 28405 29292
rect 28341 29148 28405 29212
rect 28341 29068 28405 29132
rect 28341 28988 28405 29052
rect 28341 28908 28405 28972
rect 28341 28828 28405 28892
rect 28341 28748 28405 28812
rect 28341 28668 28405 28732
rect 28341 28588 28405 28652
rect 28341 28508 28405 28572
rect 28341 28428 28405 28492
rect 34660 34508 34724 34572
rect 34660 34428 34724 34492
rect 34660 34348 34724 34412
rect 34660 34268 34724 34332
rect 34660 34188 34724 34252
rect 34660 34108 34724 34172
rect 34660 34028 34724 34092
rect 34660 33948 34724 34012
rect 34660 33868 34724 33932
rect 34660 33788 34724 33852
rect 34660 33708 34724 33772
rect 34660 33628 34724 33692
rect 34660 33548 34724 33612
rect 34660 33468 34724 33532
rect 34660 33388 34724 33452
rect 34660 33308 34724 33372
rect 34660 33228 34724 33292
rect 34660 33148 34724 33212
rect 34660 33068 34724 33132
rect 34660 32988 34724 33052
rect 34660 32908 34724 32972
rect 34660 32828 34724 32892
rect 34660 32748 34724 32812
rect 34660 32668 34724 32732
rect 34660 32588 34724 32652
rect 34660 32508 34724 32572
rect 34660 32428 34724 32492
rect 34660 32348 34724 32412
rect 34660 32268 34724 32332
rect 34660 32188 34724 32252
rect 34660 32108 34724 32172
rect 34660 32028 34724 32092
rect 34660 31948 34724 32012
rect 34660 31868 34724 31932
rect 34660 31788 34724 31852
rect 34660 31708 34724 31772
rect 34660 31628 34724 31692
rect 34660 31548 34724 31612
rect 34660 31468 34724 31532
rect 34660 31388 34724 31452
rect 34660 31308 34724 31372
rect 34660 31228 34724 31292
rect 34660 31148 34724 31212
rect 34660 31068 34724 31132
rect 34660 30988 34724 31052
rect 34660 30908 34724 30972
rect 34660 30828 34724 30892
rect 34660 30748 34724 30812
rect 34660 30668 34724 30732
rect 34660 30588 34724 30652
rect 34660 30508 34724 30572
rect 34660 30428 34724 30492
rect 34660 30348 34724 30412
rect 34660 30268 34724 30332
rect 34660 30188 34724 30252
rect 34660 30108 34724 30172
rect 34660 30028 34724 30092
rect 34660 29948 34724 30012
rect 34660 29868 34724 29932
rect 34660 29788 34724 29852
rect 34660 29708 34724 29772
rect 34660 29628 34724 29692
rect 34660 29548 34724 29612
rect 34660 29468 34724 29532
rect 34660 29388 34724 29452
rect 34660 29308 34724 29372
rect 34660 29228 34724 29292
rect 34660 29148 34724 29212
rect 34660 29068 34724 29132
rect 34660 28988 34724 29052
rect 34660 28908 34724 28972
rect 34660 28828 34724 28892
rect 34660 28748 34724 28812
rect 34660 28668 34724 28732
rect 34660 28588 34724 28652
rect 34660 28508 34724 28572
rect 34660 28428 34724 28492
rect 40979 34508 41043 34572
rect 40979 34428 41043 34492
rect 40979 34348 41043 34412
rect 40979 34268 41043 34332
rect 40979 34188 41043 34252
rect 40979 34108 41043 34172
rect 40979 34028 41043 34092
rect 40979 33948 41043 34012
rect 40979 33868 41043 33932
rect 40979 33788 41043 33852
rect 40979 33708 41043 33772
rect 40979 33628 41043 33692
rect 40979 33548 41043 33612
rect 40979 33468 41043 33532
rect 40979 33388 41043 33452
rect 40979 33308 41043 33372
rect 40979 33228 41043 33292
rect 40979 33148 41043 33212
rect 40979 33068 41043 33132
rect 40979 32988 41043 33052
rect 40979 32908 41043 32972
rect 40979 32828 41043 32892
rect 40979 32748 41043 32812
rect 40979 32668 41043 32732
rect 40979 32588 41043 32652
rect 40979 32508 41043 32572
rect 40979 32428 41043 32492
rect 40979 32348 41043 32412
rect 40979 32268 41043 32332
rect 40979 32188 41043 32252
rect 40979 32108 41043 32172
rect 40979 32028 41043 32092
rect 40979 31948 41043 32012
rect 40979 31868 41043 31932
rect 40979 31788 41043 31852
rect 40979 31708 41043 31772
rect 40979 31628 41043 31692
rect 40979 31548 41043 31612
rect 40979 31468 41043 31532
rect 40979 31388 41043 31452
rect 40979 31308 41043 31372
rect 40979 31228 41043 31292
rect 40979 31148 41043 31212
rect 40979 31068 41043 31132
rect 40979 30988 41043 31052
rect 40979 30908 41043 30972
rect 40979 30828 41043 30892
rect 40979 30748 41043 30812
rect 40979 30668 41043 30732
rect 40979 30588 41043 30652
rect 40979 30508 41043 30572
rect 40979 30428 41043 30492
rect 40979 30348 41043 30412
rect 40979 30268 41043 30332
rect 40979 30188 41043 30252
rect 40979 30108 41043 30172
rect 40979 30028 41043 30092
rect 40979 29948 41043 30012
rect 40979 29868 41043 29932
rect 40979 29788 41043 29852
rect 40979 29708 41043 29772
rect 40979 29628 41043 29692
rect 40979 29548 41043 29612
rect 40979 29468 41043 29532
rect 40979 29388 41043 29452
rect 40979 29308 41043 29372
rect 40979 29228 41043 29292
rect 40979 29148 41043 29212
rect 40979 29068 41043 29132
rect 40979 28988 41043 29052
rect 40979 28908 41043 28972
rect 40979 28828 41043 28892
rect 40979 28748 41043 28812
rect 40979 28668 41043 28732
rect 40979 28588 41043 28652
rect 40979 28508 41043 28572
rect 40979 28428 41043 28492
rect 47298 34508 47362 34572
rect 47298 34428 47362 34492
rect 47298 34348 47362 34412
rect 47298 34268 47362 34332
rect 47298 34188 47362 34252
rect 47298 34108 47362 34172
rect 47298 34028 47362 34092
rect 47298 33948 47362 34012
rect 47298 33868 47362 33932
rect 47298 33788 47362 33852
rect 47298 33708 47362 33772
rect 47298 33628 47362 33692
rect 47298 33548 47362 33612
rect 47298 33468 47362 33532
rect 47298 33388 47362 33452
rect 47298 33308 47362 33372
rect 47298 33228 47362 33292
rect 47298 33148 47362 33212
rect 47298 33068 47362 33132
rect 47298 32988 47362 33052
rect 47298 32908 47362 32972
rect 47298 32828 47362 32892
rect 47298 32748 47362 32812
rect 47298 32668 47362 32732
rect 47298 32588 47362 32652
rect 47298 32508 47362 32572
rect 47298 32428 47362 32492
rect 47298 32348 47362 32412
rect 47298 32268 47362 32332
rect 47298 32188 47362 32252
rect 47298 32108 47362 32172
rect 47298 32028 47362 32092
rect 47298 31948 47362 32012
rect 47298 31868 47362 31932
rect 47298 31788 47362 31852
rect 47298 31708 47362 31772
rect 47298 31628 47362 31692
rect 47298 31548 47362 31612
rect 47298 31468 47362 31532
rect 47298 31388 47362 31452
rect 47298 31308 47362 31372
rect 47298 31228 47362 31292
rect 47298 31148 47362 31212
rect 47298 31068 47362 31132
rect 47298 30988 47362 31052
rect 47298 30908 47362 30972
rect 47298 30828 47362 30892
rect 47298 30748 47362 30812
rect 47298 30668 47362 30732
rect 47298 30588 47362 30652
rect 47298 30508 47362 30572
rect 47298 30428 47362 30492
rect 47298 30348 47362 30412
rect 47298 30268 47362 30332
rect 47298 30188 47362 30252
rect 47298 30108 47362 30172
rect 47298 30028 47362 30092
rect 47298 29948 47362 30012
rect 47298 29868 47362 29932
rect 47298 29788 47362 29852
rect 47298 29708 47362 29772
rect 47298 29628 47362 29692
rect 47298 29548 47362 29612
rect 47298 29468 47362 29532
rect 47298 29388 47362 29452
rect 47298 29308 47362 29372
rect 47298 29228 47362 29292
rect 47298 29148 47362 29212
rect 47298 29068 47362 29132
rect 47298 28988 47362 29052
rect 47298 28908 47362 28972
rect 47298 28828 47362 28892
rect 47298 28748 47362 28812
rect 47298 28668 47362 28732
rect 47298 28588 47362 28652
rect 47298 28508 47362 28572
rect 47298 28428 47362 28492
rect -41168 28208 -41104 28272
rect -41168 28128 -41104 28192
rect -41168 28048 -41104 28112
rect -41168 27968 -41104 28032
rect -41168 27888 -41104 27952
rect -41168 27808 -41104 27872
rect -41168 27728 -41104 27792
rect -41168 27648 -41104 27712
rect -41168 27568 -41104 27632
rect -41168 27488 -41104 27552
rect -41168 27408 -41104 27472
rect -41168 27328 -41104 27392
rect -41168 27248 -41104 27312
rect -41168 27168 -41104 27232
rect -41168 27088 -41104 27152
rect -41168 27008 -41104 27072
rect -41168 26928 -41104 26992
rect -41168 26848 -41104 26912
rect -41168 26768 -41104 26832
rect -41168 26688 -41104 26752
rect -41168 26608 -41104 26672
rect -41168 26528 -41104 26592
rect -41168 26448 -41104 26512
rect -41168 26368 -41104 26432
rect -41168 26288 -41104 26352
rect -41168 26208 -41104 26272
rect -41168 26128 -41104 26192
rect -41168 26048 -41104 26112
rect -41168 25968 -41104 26032
rect -41168 25888 -41104 25952
rect -41168 25808 -41104 25872
rect -41168 25728 -41104 25792
rect -41168 25648 -41104 25712
rect -41168 25568 -41104 25632
rect -41168 25488 -41104 25552
rect -41168 25408 -41104 25472
rect -41168 25328 -41104 25392
rect -41168 25248 -41104 25312
rect -41168 25168 -41104 25232
rect -41168 25088 -41104 25152
rect -41168 25008 -41104 25072
rect -41168 24928 -41104 24992
rect -41168 24848 -41104 24912
rect -41168 24768 -41104 24832
rect -41168 24688 -41104 24752
rect -41168 24608 -41104 24672
rect -41168 24528 -41104 24592
rect -41168 24448 -41104 24512
rect -41168 24368 -41104 24432
rect -41168 24288 -41104 24352
rect -41168 24208 -41104 24272
rect -41168 24128 -41104 24192
rect -41168 24048 -41104 24112
rect -41168 23968 -41104 24032
rect -41168 23888 -41104 23952
rect -41168 23808 -41104 23872
rect -41168 23728 -41104 23792
rect -41168 23648 -41104 23712
rect -41168 23568 -41104 23632
rect -41168 23488 -41104 23552
rect -41168 23408 -41104 23472
rect -41168 23328 -41104 23392
rect -41168 23248 -41104 23312
rect -41168 23168 -41104 23232
rect -41168 23088 -41104 23152
rect -41168 23008 -41104 23072
rect -41168 22928 -41104 22992
rect -41168 22848 -41104 22912
rect -41168 22768 -41104 22832
rect -41168 22688 -41104 22752
rect -41168 22608 -41104 22672
rect -41168 22528 -41104 22592
rect -41168 22448 -41104 22512
rect -41168 22368 -41104 22432
rect -41168 22288 -41104 22352
rect -41168 22208 -41104 22272
rect -41168 22128 -41104 22192
rect -34849 28208 -34785 28272
rect -34849 28128 -34785 28192
rect -34849 28048 -34785 28112
rect -34849 27968 -34785 28032
rect -34849 27888 -34785 27952
rect -34849 27808 -34785 27872
rect -34849 27728 -34785 27792
rect -34849 27648 -34785 27712
rect -34849 27568 -34785 27632
rect -34849 27488 -34785 27552
rect -34849 27408 -34785 27472
rect -34849 27328 -34785 27392
rect -34849 27248 -34785 27312
rect -34849 27168 -34785 27232
rect -34849 27088 -34785 27152
rect -34849 27008 -34785 27072
rect -34849 26928 -34785 26992
rect -34849 26848 -34785 26912
rect -34849 26768 -34785 26832
rect -34849 26688 -34785 26752
rect -34849 26608 -34785 26672
rect -34849 26528 -34785 26592
rect -34849 26448 -34785 26512
rect -34849 26368 -34785 26432
rect -34849 26288 -34785 26352
rect -34849 26208 -34785 26272
rect -34849 26128 -34785 26192
rect -34849 26048 -34785 26112
rect -34849 25968 -34785 26032
rect -34849 25888 -34785 25952
rect -34849 25808 -34785 25872
rect -34849 25728 -34785 25792
rect -34849 25648 -34785 25712
rect -34849 25568 -34785 25632
rect -34849 25488 -34785 25552
rect -34849 25408 -34785 25472
rect -34849 25328 -34785 25392
rect -34849 25248 -34785 25312
rect -34849 25168 -34785 25232
rect -34849 25088 -34785 25152
rect -34849 25008 -34785 25072
rect -34849 24928 -34785 24992
rect -34849 24848 -34785 24912
rect -34849 24768 -34785 24832
rect -34849 24688 -34785 24752
rect -34849 24608 -34785 24672
rect -34849 24528 -34785 24592
rect -34849 24448 -34785 24512
rect -34849 24368 -34785 24432
rect -34849 24288 -34785 24352
rect -34849 24208 -34785 24272
rect -34849 24128 -34785 24192
rect -34849 24048 -34785 24112
rect -34849 23968 -34785 24032
rect -34849 23888 -34785 23952
rect -34849 23808 -34785 23872
rect -34849 23728 -34785 23792
rect -34849 23648 -34785 23712
rect -34849 23568 -34785 23632
rect -34849 23488 -34785 23552
rect -34849 23408 -34785 23472
rect -34849 23328 -34785 23392
rect -34849 23248 -34785 23312
rect -34849 23168 -34785 23232
rect -34849 23088 -34785 23152
rect -34849 23008 -34785 23072
rect -34849 22928 -34785 22992
rect -34849 22848 -34785 22912
rect -34849 22768 -34785 22832
rect -34849 22688 -34785 22752
rect -34849 22608 -34785 22672
rect -34849 22528 -34785 22592
rect -34849 22448 -34785 22512
rect -34849 22368 -34785 22432
rect -34849 22288 -34785 22352
rect -34849 22208 -34785 22272
rect -34849 22128 -34785 22192
rect -28530 28208 -28466 28272
rect -28530 28128 -28466 28192
rect -28530 28048 -28466 28112
rect -28530 27968 -28466 28032
rect -28530 27888 -28466 27952
rect -28530 27808 -28466 27872
rect -28530 27728 -28466 27792
rect -28530 27648 -28466 27712
rect -28530 27568 -28466 27632
rect -28530 27488 -28466 27552
rect -28530 27408 -28466 27472
rect -28530 27328 -28466 27392
rect -28530 27248 -28466 27312
rect -28530 27168 -28466 27232
rect -28530 27088 -28466 27152
rect -28530 27008 -28466 27072
rect -28530 26928 -28466 26992
rect -28530 26848 -28466 26912
rect -28530 26768 -28466 26832
rect -28530 26688 -28466 26752
rect -28530 26608 -28466 26672
rect -28530 26528 -28466 26592
rect -28530 26448 -28466 26512
rect -28530 26368 -28466 26432
rect -28530 26288 -28466 26352
rect -28530 26208 -28466 26272
rect -28530 26128 -28466 26192
rect -28530 26048 -28466 26112
rect -28530 25968 -28466 26032
rect -28530 25888 -28466 25952
rect -28530 25808 -28466 25872
rect -28530 25728 -28466 25792
rect -28530 25648 -28466 25712
rect -28530 25568 -28466 25632
rect -28530 25488 -28466 25552
rect -28530 25408 -28466 25472
rect -28530 25328 -28466 25392
rect -28530 25248 -28466 25312
rect -28530 25168 -28466 25232
rect -28530 25088 -28466 25152
rect -28530 25008 -28466 25072
rect -28530 24928 -28466 24992
rect -28530 24848 -28466 24912
rect -28530 24768 -28466 24832
rect -28530 24688 -28466 24752
rect -28530 24608 -28466 24672
rect -28530 24528 -28466 24592
rect -28530 24448 -28466 24512
rect -28530 24368 -28466 24432
rect -28530 24288 -28466 24352
rect -28530 24208 -28466 24272
rect -28530 24128 -28466 24192
rect -28530 24048 -28466 24112
rect -28530 23968 -28466 24032
rect -28530 23888 -28466 23952
rect -28530 23808 -28466 23872
rect -28530 23728 -28466 23792
rect -28530 23648 -28466 23712
rect -28530 23568 -28466 23632
rect -28530 23488 -28466 23552
rect -28530 23408 -28466 23472
rect -28530 23328 -28466 23392
rect -28530 23248 -28466 23312
rect -28530 23168 -28466 23232
rect -28530 23088 -28466 23152
rect -28530 23008 -28466 23072
rect -28530 22928 -28466 22992
rect -28530 22848 -28466 22912
rect -28530 22768 -28466 22832
rect -28530 22688 -28466 22752
rect -28530 22608 -28466 22672
rect -28530 22528 -28466 22592
rect -28530 22448 -28466 22512
rect -28530 22368 -28466 22432
rect -28530 22288 -28466 22352
rect -28530 22208 -28466 22272
rect -28530 22128 -28466 22192
rect -22211 28208 -22147 28272
rect -22211 28128 -22147 28192
rect -22211 28048 -22147 28112
rect -22211 27968 -22147 28032
rect -22211 27888 -22147 27952
rect -22211 27808 -22147 27872
rect -22211 27728 -22147 27792
rect -22211 27648 -22147 27712
rect -22211 27568 -22147 27632
rect -22211 27488 -22147 27552
rect -22211 27408 -22147 27472
rect -22211 27328 -22147 27392
rect -22211 27248 -22147 27312
rect -22211 27168 -22147 27232
rect -22211 27088 -22147 27152
rect -22211 27008 -22147 27072
rect -22211 26928 -22147 26992
rect -22211 26848 -22147 26912
rect -22211 26768 -22147 26832
rect -22211 26688 -22147 26752
rect -22211 26608 -22147 26672
rect -22211 26528 -22147 26592
rect -22211 26448 -22147 26512
rect -22211 26368 -22147 26432
rect -22211 26288 -22147 26352
rect -22211 26208 -22147 26272
rect -22211 26128 -22147 26192
rect -22211 26048 -22147 26112
rect -22211 25968 -22147 26032
rect -22211 25888 -22147 25952
rect -22211 25808 -22147 25872
rect -22211 25728 -22147 25792
rect -22211 25648 -22147 25712
rect -22211 25568 -22147 25632
rect -22211 25488 -22147 25552
rect -22211 25408 -22147 25472
rect -22211 25328 -22147 25392
rect -22211 25248 -22147 25312
rect -22211 25168 -22147 25232
rect -22211 25088 -22147 25152
rect -22211 25008 -22147 25072
rect -22211 24928 -22147 24992
rect -22211 24848 -22147 24912
rect -22211 24768 -22147 24832
rect -22211 24688 -22147 24752
rect -22211 24608 -22147 24672
rect -22211 24528 -22147 24592
rect -22211 24448 -22147 24512
rect -22211 24368 -22147 24432
rect -22211 24288 -22147 24352
rect -22211 24208 -22147 24272
rect -22211 24128 -22147 24192
rect -22211 24048 -22147 24112
rect -22211 23968 -22147 24032
rect -22211 23888 -22147 23952
rect -22211 23808 -22147 23872
rect -22211 23728 -22147 23792
rect -22211 23648 -22147 23712
rect -22211 23568 -22147 23632
rect -22211 23488 -22147 23552
rect -22211 23408 -22147 23472
rect -22211 23328 -22147 23392
rect -22211 23248 -22147 23312
rect -22211 23168 -22147 23232
rect -22211 23088 -22147 23152
rect -22211 23008 -22147 23072
rect -22211 22928 -22147 22992
rect -22211 22848 -22147 22912
rect -22211 22768 -22147 22832
rect -22211 22688 -22147 22752
rect -22211 22608 -22147 22672
rect -22211 22528 -22147 22592
rect -22211 22448 -22147 22512
rect -22211 22368 -22147 22432
rect -22211 22288 -22147 22352
rect -22211 22208 -22147 22272
rect -22211 22128 -22147 22192
rect -15892 28208 -15828 28272
rect -15892 28128 -15828 28192
rect -15892 28048 -15828 28112
rect -15892 27968 -15828 28032
rect -15892 27888 -15828 27952
rect -15892 27808 -15828 27872
rect -15892 27728 -15828 27792
rect -15892 27648 -15828 27712
rect -15892 27568 -15828 27632
rect -15892 27488 -15828 27552
rect -15892 27408 -15828 27472
rect -15892 27328 -15828 27392
rect -15892 27248 -15828 27312
rect -15892 27168 -15828 27232
rect -15892 27088 -15828 27152
rect -15892 27008 -15828 27072
rect -15892 26928 -15828 26992
rect -15892 26848 -15828 26912
rect -15892 26768 -15828 26832
rect -15892 26688 -15828 26752
rect -15892 26608 -15828 26672
rect -15892 26528 -15828 26592
rect -15892 26448 -15828 26512
rect -15892 26368 -15828 26432
rect -15892 26288 -15828 26352
rect -15892 26208 -15828 26272
rect -15892 26128 -15828 26192
rect -15892 26048 -15828 26112
rect -15892 25968 -15828 26032
rect -15892 25888 -15828 25952
rect -15892 25808 -15828 25872
rect -15892 25728 -15828 25792
rect -15892 25648 -15828 25712
rect -15892 25568 -15828 25632
rect -15892 25488 -15828 25552
rect -15892 25408 -15828 25472
rect -15892 25328 -15828 25392
rect -15892 25248 -15828 25312
rect -15892 25168 -15828 25232
rect -15892 25088 -15828 25152
rect -15892 25008 -15828 25072
rect -15892 24928 -15828 24992
rect -15892 24848 -15828 24912
rect -15892 24768 -15828 24832
rect -15892 24688 -15828 24752
rect -15892 24608 -15828 24672
rect -15892 24528 -15828 24592
rect -15892 24448 -15828 24512
rect -15892 24368 -15828 24432
rect -15892 24288 -15828 24352
rect -15892 24208 -15828 24272
rect -15892 24128 -15828 24192
rect -15892 24048 -15828 24112
rect -15892 23968 -15828 24032
rect -15892 23888 -15828 23952
rect -15892 23808 -15828 23872
rect -15892 23728 -15828 23792
rect -15892 23648 -15828 23712
rect -15892 23568 -15828 23632
rect -15892 23488 -15828 23552
rect -15892 23408 -15828 23472
rect -15892 23328 -15828 23392
rect -15892 23248 -15828 23312
rect -15892 23168 -15828 23232
rect -15892 23088 -15828 23152
rect -15892 23008 -15828 23072
rect -15892 22928 -15828 22992
rect -15892 22848 -15828 22912
rect -15892 22768 -15828 22832
rect -15892 22688 -15828 22752
rect -15892 22608 -15828 22672
rect -15892 22528 -15828 22592
rect -15892 22448 -15828 22512
rect -15892 22368 -15828 22432
rect -15892 22288 -15828 22352
rect -15892 22208 -15828 22272
rect -15892 22128 -15828 22192
rect -9573 28208 -9509 28272
rect -9573 28128 -9509 28192
rect -9573 28048 -9509 28112
rect -9573 27968 -9509 28032
rect -9573 27888 -9509 27952
rect -9573 27808 -9509 27872
rect -9573 27728 -9509 27792
rect -9573 27648 -9509 27712
rect -9573 27568 -9509 27632
rect -9573 27488 -9509 27552
rect -9573 27408 -9509 27472
rect -9573 27328 -9509 27392
rect -9573 27248 -9509 27312
rect -9573 27168 -9509 27232
rect -9573 27088 -9509 27152
rect -9573 27008 -9509 27072
rect -9573 26928 -9509 26992
rect -9573 26848 -9509 26912
rect -9573 26768 -9509 26832
rect -9573 26688 -9509 26752
rect -9573 26608 -9509 26672
rect -9573 26528 -9509 26592
rect -9573 26448 -9509 26512
rect -9573 26368 -9509 26432
rect -9573 26288 -9509 26352
rect -9573 26208 -9509 26272
rect -9573 26128 -9509 26192
rect -9573 26048 -9509 26112
rect -9573 25968 -9509 26032
rect -9573 25888 -9509 25952
rect -9573 25808 -9509 25872
rect -9573 25728 -9509 25792
rect -9573 25648 -9509 25712
rect -9573 25568 -9509 25632
rect -9573 25488 -9509 25552
rect -9573 25408 -9509 25472
rect -9573 25328 -9509 25392
rect -9573 25248 -9509 25312
rect -9573 25168 -9509 25232
rect -9573 25088 -9509 25152
rect -9573 25008 -9509 25072
rect -9573 24928 -9509 24992
rect -9573 24848 -9509 24912
rect -9573 24768 -9509 24832
rect -9573 24688 -9509 24752
rect -9573 24608 -9509 24672
rect -9573 24528 -9509 24592
rect -9573 24448 -9509 24512
rect -9573 24368 -9509 24432
rect -9573 24288 -9509 24352
rect -9573 24208 -9509 24272
rect -9573 24128 -9509 24192
rect -9573 24048 -9509 24112
rect -9573 23968 -9509 24032
rect -9573 23888 -9509 23952
rect -9573 23808 -9509 23872
rect -9573 23728 -9509 23792
rect -9573 23648 -9509 23712
rect -9573 23568 -9509 23632
rect -9573 23488 -9509 23552
rect -9573 23408 -9509 23472
rect -9573 23328 -9509 23392
rect -9573 23248 -9509 23312
rect -9573 23168 -9509 23232
rect -9573 23088 -9509 23152
rect -9573 23008 -9509 23072
rect -9573 22928 -9509 22992
rect -9573 22848 -9509 22912
rect -9573 22768 -9509 22832
rect -9573 22688 -9509 22752
rect -9573 22608 -9509 22672
rect -9573 22528 -9509 22592
rect -9573 22448 -9509 22512
rect -9573 22368 -9509 22432
rect -9573 22288 -9509 22352
rect -9573 22208 -9509 22272
rect -9573 22128 -9509 22192
rect -3254 28208 -3190 28272
rect -3254 28128 -3190 28192
rect -3254 28048 -3190 28112
rect -3254 27968 -3190 28032
rect -3254 27888 -3190 27952
rect -3254 27808 -3190 27872
rect -3254 27728 -3190 27792
rect -3254 27648 -3190 27712
rect -3254 27568 -3190 27632
rect -3254 27488 -3190 27552
rect -3254 27408 -3190 27472
rect -3254 27328 -3190 27392
rect -3254 27248 -3190 27312
rect -3254 27168 -3190 27232
rect -3254 27088 -3190 27152
rect -3254 27008 -3190 27072
rect -3254 26928 -3190 26992
rect -3254 26848 -3190 26912
rect -3254 26768 -3190 26832
rect -3254 26688 -3190 26752
rect -3254 26608 -3190 26672
rect -3254 26528 -3190 26592
rect -3254 26448 -3190 26512
rect -3254 26368 -3190 26432
rect -3254 26288 -3190 26352
rect -3254 26208 -3190 26272
rect -3254 26128 -3190 26192
rect -3254 26048 -3190 26112
rect -3254 25968 -3190 26032
rect -3254 25888 -3190 25952
rect -3254 25808 -3190 25872
rect -3254 25728 -3190 25792
rect -3254 25648 -3190 25712
rect -3254 25568 -3190 25632
rect -3254 25488 -3190 25552
rect -3254 25408 -3190 25472
rect -3254 25328 -3190 25392
rect -3254 25248 -3190 25312
rect -3254 25168 -3190 25232
rect -3254 25088 -3190 25152
rect -3254 25008 -3190 25072
rect -3254 24928 -3190 24992
rect -3254 24848 -3190 24912
rect -3254 24768 -3190 24832
rect -3254 24688 -3190 24752
rect -3254 24608 -3190 24672
rect -3254 24528 -3190 24592
rect -3254 24448 -3190 24512
rect -3254 24368 -3190 24432
rect -3254 24288 -3190 24352
rect -3254 24208 -3190 24272
rect -3254 24128 -3190 24192
rect -3254 24048 -3190 24112
rect -3254 23968 -3190 24032
rect -3254 23888 -3190 23952
rect -3254 23808 -3190 23872
rect -3254 23728 -3190 23792
rect -3254 23648 -3190 23712
rect -3254 23568 -3190 23632
rect -3254 23488 -3190 23552
rect -3254 23408 -3190 23472
rect -3254 23328 -3190 23392
rect -3254 23248 -3190 23312
rect -3254 23168 -3190 23232
rect -3254 23088 -3190 23152
rect -3254 23008 -3190 23072
rect -3254 22928 -3190 22992
rect -3254 22848 -3190 22912
rect -3254 22768 -3190 22832
rect -3254 22688 -3190 22752
rect -3254 22608 -3190 22672
rect -3254 22528 -3190 22592
rect -3254 22448 -3190 22512
rect -3254 22368 -3190 22432
rect -3254 22288 -3190 22352
rect -3254 22208 -3190 22272
rect -3254 22128 -3190 22192
rect 3065 28208 3129 28272
rect 3065 28128 3129 28192
rect 3065 28048 3129 28112
rect 3065 27968 3129 28032
rect 3065 27888 3129 27952
rect 3065 27808 3129 27872
rect 3065 27728 3129 27792
rect 3065 27648 3129 27712
rect 3065 27568 3129 27632
rect 3065 27488 3129 27552
rect 3065 27408 3129 27472
rect 3065 27328 3129 27392
rect 3065 27248 3129 27312
rect 3065 27168 3129 27232
rect 3065 27088 3129 27152
rect 3065 27008 3129 27072
rect 3065 26928 3129 26992
rect 3065 26848 3129 26912
rect 3065 26768 3129 26832
rect 3065 26688 3129 26752
rect 3065 26608 3129 26672
rect 3065 26528 3129 26592
rect 3065 26448 3129 26512
rect 3065 26368 3129 26432
rect 3065 26288 3129 26352
rect 3065 26208 3129 26272
rect 3065 26128 3129 26192
rect 3065 26048 3129 26112
rect 3065 25968 3129 26032
rect 3065 25888 3129 25952
rect 3065 25808 3129 25872
rect 3065 25728 3129 25792
rect 3065 25648 3129 25712
rect 3065 25568 3129 25632
rect 3065 25488 3129 25552
rect 3065 25408 3129 25472
rect 3065 25328 3129 25392
rect 3065 25248 3129 25312
rect 3065 25168 3129 25232
rect 3065 25088 3129 25152
rect 3065 25008 3129 25072
rect 3065 24928 3129 24992
rect 3065 24848 3129 24912
rect 3065 24768 3129 24832
rect 3065 24688 3129 24752
rect 3065 24608 3129 24672
rect 3065 24528 3129 24592
rect 3065 24448 3129 24512
rect 3065 24368 3129 24432
rect 3065 24288 3129 24352
rect 3065 24208 3129 24272
rect 3065 24128 3129 24192
rect 3065 24048 3129 24112
rect 3065 23968 3129 24032
rect 3065 23888 3129 23952
rect 3065 23808 3129 23872
rect 3065 23728 3129 23792
rect 3065 23648 3129 23712
rect 3065 23568 3129 23632
rect 3065 23488 3129 23552
rect 3065 23408 3129 23472
rect 3065 23328 3129 23392
rect 3065 23248 3129 23312
rect 3065 23168 3129 23232
rect 3065 23088 3129 23152
rect 3065 23008 3129 23072
rect 3065 22928 3129 22992
rect 3065 22848 3129 22912
rect 3065 22768 3129 22832
rect 3065 22688 3129 22752
rect 3065 22608 3129 22672
rect 3065 22528 3129 22592
rect 3065 22448 3129 22512
rect 3065 22368 3129 22432
rect 3065 22288 3129 22352
rect 3065 22208 3129 22272
rect 3065 22128 3129 22192
rect 9384 28208 9448 28272
rect 9384 28128 9448 28192
rect 9384 28048 9448 28112
rect 9384 27968 9448 28032
rect 9384 27888 9448 27952
rect 9384 27808 9448 27872
rect 9384 27728 9448 27792
rect 9384 27648 9448 27712
rect 9384 27568 9448 27632
rect 9384 27488 9448 27552
rect 9384 27408 9448 27472
rect 9384 27328 9448 27392
rect 9384 27248 9448 27312
rect 9384 27168 9448 27232
rect 9384 27088 9448 27152
rect 9384 27008 9448 27072
rect 9384 26928 9448 26992
rect 9384 26848 9448 26912
rect 9384 26768 9448 26832
rect 9384 26688 9448 26752
rect 9384 26608 9448 26672
rect 9384 26528 9448 26592
rect 9384 26448 9448 26512
rect 9384 26368 9448 26432
rect 9384 26288 9448 26352
rect 9384 26208 9448 26272
rect 9384 26128 9448 26192
rect 9384 26048 9448 26112
rect 9384 25968 9448 26032
rect 9384 25888 9448 25952
rect 9384 25808 9448 25872
rect 9384 25728 9448 25792
rect 9384 25648 9448 25712
rect 9384 25568 9448 25632
rect 9384 25488 9448 25552
rect 9384 25408 9448 25472
rect 9384 25328 9448 25392
rect 9384 25248 9448 25312
rect 9384 25168 9448 25232
rect 9384 25088 9448 25152
rect 9384 25008 9448 25072
rect 9384 24928 9448 24992
rect 9384 24848 9448 24912
rect 9384 24768 9448 24832
rect 9384 24688 9448 24752
rect 9384 24608 9448 24672
rect 9384 24528 9448 24592
rect 9384 24448 9448 24512
rect 9384 24368 9448 24432
rect 9384 24288 9448 24352
rect 9384 24208 9448 24272
rect 9384 24128 9448 24192
rect 9384 24048 9448 24112
rect 9384 23968 9448 24032
rect 9384 23888 9448 23952
rect 9384 23808 9448 23872
rect 9384 23728 9448 23792
rect 9384 23648 9448 23712
rect 9384 23568 9448 23632
rect 9384 23488 9448 23552
rect 9384 23408 9448 23472
rect 9384 23328 9448 23392
rect 9384 23248 9448 23312
rect 9384 23168 9448 23232
rect 9384 23088 9448 23152
rect 9384 23008 9448 23072
rect 9384 22928 9448 22992
rect 9384 22848 9448 22912
rect 9384 22768 9448 22832
rect 9384 22688 9448 22752
rect 9384 22608 9448 22672
rect 9384 22528 9448 22592
rect 9384 22448 9448 22512
rect 9384 22368 9448 22432
rect 9384 22288 9448 22352
rect 9384 22208 9448 22272
rect 9384 22128 9448 22192
rect 15703 28208 15767 28272
rect 15703 28128 15767 28192
rect 15703 28048 15767 28112
rect 15703 27968 15767 28032
rect 15703 27888 15767 27952
rect 15703 27808 15767 27872
rect 15703 27728 15767 27792
rect 15703 27648 15767 27712
rect 15703 27568 15767 27632
rect 15703 27488 15767 27552
rect 15703 27408 15767 27472
rect 15703 27328 15767 27392
rect 15703 27248 15767 27312
rect 15703 27168 15767 27232
rect 15703 27088 15767 27152
rect 15703 27008 15767 27072
rect 15703 26928 15767 26992
rect 15703 26848 15767 26912
rect 15703 26768 15767 26832
rect 15703 26688 15767 26752
rect 15703 26608 15767 26672
rect 15703 26528 15767 26592
rect 15703 26448 15767 26512
rect 15703 26368 15767 26432
rect 15703 26288 15767 26352
rect 15703 26208 15767 26272
rect 15703 26128 15767 26192
rect 15703 26048 15767 26112
rect 15703 25968 15767 26032
rect 15703 25888 15767 25952
rect 15703 25808 15767 25872
rect 15703 25728 15767 25792
rect 15703 25648 15767 25712
rect 15703 25568 15767 25632
rect 15703 25488 15767 25552
rect 15703 25408 15767 25472
rect 15703 25328 15767 25392
rect 15703 25248 15767 25312
rect 15703 25168 15767 25232
rect 15703 25088 15767 25152
rect 15703 25008 15767 25072
rect 15703 24928 15767 24992
rect 15703 24848 15767 24912
rect 15703 24768 15767 24832
rect 15703 24688 15767 24752
rect 15703 24608 15767 24672
rect 15703 24528 15767 24592
rect 15703 24448 15767 24512
rect 15703 24368 15767 24432
rect 15703 24288 15767 24352
rect 15703 24208 15767 24272
rect 15703 24128 15767 24192
rect 15703 24048 15767 24112
rect 15703 23968 15767 24032
rect 15703 23888 15767 23952
rect 15703 23808 15767 23872
rect 15703 23728 15767 23792
rect 15703 23648 15767 23712
rect 15703 23568 15767 23632
rect 15703 23488 15767 23552
rect 15703 23408 15767 23472
rect 15703 23328 15767 23392
rect 15703 23248 15767 23312
rect 15703 23168 15767 23232
rect 15703 23088 15767 23152
rect 15703 23008 15767 23072
rect 15703 22928 15767 22992
rect 15703 22848 15767 22912
rect 15703 22768 15767 22832
rect 15703 22688 15767 22752
rect 15703 22608 15767 22672
rect 15703 22528 15767 22592
rect 15703 22448 15767 22512
rect 15703 22368 15767 22432
rect 15703 22288 15767 22352
rect 15703 22208 15767 22272
rect 15703 22128 15767 22192
rect 22022 28208 22086 28272
rect 22022 28128 22086 28192
rect 22022 28048 22086 28112
rect 22022 27968 22086 28032
rect 22022 27888 22086 27952
rect 22022 27808 22086 27872
rect 22022 27728 22086 27792
rect 22022 27648 22086 27712
rect 22022 27568 22086 27632
rect 22022 27488 22086 27552
rect 22022 27408 22086 27472
rect 22022 27328 22086 27392
rect 22022 27248 22086 27312
rect 22022 27168 22086 27232
rect 22022 27088 22086 27152
rect 22022 27008 22086 27072
rect 22022 26928 22086 26992
rect 22022 26848 22086 26912
rect 22022 26768 22086 26832
rect 22022 26688 22086 26752
rect 22022 26608 22086 26672
rect 22022 26528 22086 26592
rect 22022 26448 22086 26512
rect 22022 26368 22086 26432
rect 22022 26288 22086 26352
rect 22022 26208 22086 26272
rect 22022 26128 22086 26192
rect 22022 26048 22086 26112
rect 22022 25968 22086 26032
rect 22022 25888 22086 25952
rect 22022 25808 22086 25872
rect 22022 25728 22086 25792
rect 22022 25648 22086 25712
rect 22022 25568 22086 25632
rect 22022 25488 22086 25552
rect 22022 25408 22086 25472
rect 22022 25328 22086 25392
rect 22022 25248 22086 25312
rect 22022 25168 22086 25232
rect 22022 25088 22086 25152
rect 22022 25008 22086 25072
rect 22022 24928 22086 24992
rect 22022 24848 22086 24912
rect 22022 24768 22086 24832
rect 22022 24688 22086 24752
rect 22022 24608 22086 24672
rect 22022 24528 22086 24592
rect 22022 24448 22086 24512
rect 22022 24368 22086 24432
rect 22022 24288 22086 24352
rect 22022 24208 22086 24272
rect 22022 24128 22086 24192
rect 22022 24048 22086 24112
rect 22022 23968 22086 24032
rect 22022 23888 22086 23952
rect 22022 23808 22086 23872
rect 22022 23728 22086 23792
rect 22022 23648 22086 23712
rect 22022 23568 22086 23632
rect 22022 23488 22086 23552
rect 22022 23408 22086 23472
rect 22022 23328 22086 23392
rect 22022 23248 22086 23312
rect 22022 23168 22086 23232
rect 22022 23088 22086 23152
rect 22022 23008 22086 23072
rect 22022 22928 22086 22992
rect 22022 22848 22086 22912
rect 22022 22768 22086 22832
rect 22022 22688 22086 22752
rect 22022 22608 22086 22672
rect 22022 22528 22086 22592
rect 22022 22448 22086 22512
rect 22022 22368 22086 22432
rect 22022 22288 22086 22352
rect 22022 22208 22086 22272
rect 22022 22128 22086 22192
rect 28341 28208 28405 28272
rect 28341 28128 28405 28192
rect 28341 28048 28405 28112
rect 28341 27968 28405 28032
rect 28341 27888 28405 27952
rect 28341 27808 28405 27872
rect 28341 27728 28405 27792
rect 28341 27648 28405 27712
rect 28341 27568 28405 27632
rect 28341 27488 28405 27552
rect 28341 27408 28405 27472
rect 28341 27328 28405 27392
rect 28341 27248 28405 27312
rect 28341 27168 28405 27232
rect 28341 27088 28405 27152
rect 28341 27008 28405 27072
rect 28341 26928 28405 26992
rect 28341 26848 28405 26912
rect 28341 26768 28405 26832
rect 28341 26688 28405 26752
rect 28341 26608 28405 26672
rect 28341 26528 28405 26592
rect 28341 26448 28405 26512
rect 28341 26368 28405 26432
rect 28341 26288 28405 26352
rect 28341 26208 28405 26272
rect 28341 26128 28405 26192
rect 28341 26048 28405 26112
rect 28341 25968 28405 26032
rect 28341 25888 28405 25952
rect 28341 25808 28405 25872
rect 28341 25728 28405 25792
rect 28341 25648 28405 25712
rect 28341 25568 28405 25632
rect 28341 25488 28405 25552
rect 28341 25408 28405 25472
rect 28341 25328 28405 25392
rect 28341 25248 28405 25312
rect 28341 25168 28405 25232
rect 28341 25088 28405 25152
rect 28341 25008 28405 25072
rect 28341 24928 28405 24992
rect 28341 24848 28405 24912
rect 28341 24768 28405 24832
rect 28341 24688 28405 24752
rect 28341 24608 28405 24672
rect 28341 24528 28405 24592
rect 28341 24448 28405 24512
rect 28341 24368 28405 24432
rect 28341 24288 28405 24352
rect 28341 24208 28405 24272
rect 28341 24128 28405 24192
rect 28341 24048 28405 24112
rect 28341 23968 28405 24032
rect 28341 23888 28405 23952
rect 28341 23808 28405 23872
rect 28341 23728 28405 23792
rect 28341 23648 28405 23712
rect 28341 23568 28405 23632
rect 28341 23488 28405 23552
rect 28341 23408 28405 23472
rect 28341 23328 28405 23392
rect 28341 23248 28405 23312
rect 28341 23168 28405 23232
rect 28341 23088 28405 23152
rect 28341 23008 28405 23072
rect 28341 22928 28405 22992
rect 28341 22848 28405 22912
rect 28341 22768 28405 22832
rect 28341 22688 28405 22752
rect 28341 22608 28405 22672
rect 28341 22528 28405 22592
rect 28341 22448 28405 22512
rect 28341 22368 28405 22432
rect 28341 22288 28405 22352
rect 28341 22208 28405 22272
rect 28341 22128 28405 22192
rect 34660 28208 34724 28272
rect 34660 28128 34724 28192
rect 34660 28048 34724 28112
rect 34660 27968 34724 28032
rect 34660 27888 34724 27952
rect 34660 27808 34724 27872
rect 34660 27728 34724 27792
rect 34660 27648 34724 27712
rect 34660 27568 34724 27632
rect 34660 27488 34724 27552
rect 34660 27408 34724 27472
rect 34660 27328 34724 27392
rect 34660 27248 34724 27312
rect 34660 27168 34724 27232
rect 34660 27088 34724 27152
rect 34660 27008 34724 27072
rect 34660 26928 34724 26992
rect 34660 26848 34724 26912
rect 34660 26768 34724 26832
rect 34660 26688 34724 26752
rect 34660 26608 34724 26672
rect 34660 26528 34724 26592
rect 34660 26448 34724 26512
rect 34660 26368 34724 26432
rect 34660 26288 34724 26352
rect 34660 26208 34724 26272
rect 34660 26128 34724 26192
rect 34660 26048 34724 26112
rect 34660 25968 34724 26032
rect 34660 25888 34724 25952
rect 34660 25808 34724 25872
rect 34660 25728 34724 25792
rect 34660 25648 34724 25712
rect 34660 25568 34724 25632
rect 34660 25488 34724 25552
rect 34660 25408 34724 25472
rect 34660 25328 34724 25392
rect 34660 25248 34724 25312
rect 34660 25168 34724 25232
rect 34660 25088 34724 25152
rect 34660 25008 34724 25072
rect 34660 24928 34724 24992
rect 34660 24848 34724 24912
rect 34660 24768 34724 24832
rect 34660 24688 34724 24752
rect 34660 24608 34724 24672
rect 34660 24528 34724 24592
rect 34660 24448 34724 24512
rect 34660 24368 34724 24432
rect 34660 24288 34724 24352
rect 34660 24208 34724 24272
rect 34660 24128 34724 24192
rect 34660 24048 34724 24112
rect 34660 23968 34724 24032
rect 34660 23888 34724 23952
rect 34660 23808 34724 23872
rect 34660 23728 34724 23792
rect 34660 23648 34724 23712
rect 34660 23568 34724 23632
rect 34660 23488 34724 23552
rect 34660 23408 34724 23472
rect 34660 23328 34724 23392
rect 34660 23248 34724 23312
rect 34660 23168 34724 23232
rect 34660 23088 34724 23152
rect 34660 23008 34724 23072
rect 34660 22928 34724 22992
rect 34660 22848 34724 22912
rect 34660 22768 34724 22832
rect 34660 22688 34724 22752
rect 34660 22608 34724 22672
rect 34660 22528 34724 22592
rect 34660 22448 34724 22512
rect 34660 22368 34724 22432
rect 34660 22288 34724 22352
rect 34660 22208 34724 22272
rect 34660 22128 34724 22192
rect 40979 28208 41043 28272
rect 40979 28128 41043 28192
rect 40979 28048 41043 28112
rect 40979 27968 41043 28032
rect 40979 27888 41043 27952
rect 40979 27808 41043 27872
rect 40979 27728 41043 27792
rect 40979 27648 41043 27712
rect 40979 27568 41043 27632
rect 40979 27488 41043 27552
rect 40979 27408 41043 27472
rect 40979 27328 41043 27392
rect 40979 27248 41043 27312
rect 40979 27168 41043 27232
rect 40979 27088 41043 27152
rect 40979 27008 41043 27072
rect 40979 26928 41043 26992
rect 40979 26848 41043 26912
rect 40979 26768 41043 26832
rect 40979 26688 41043 26752
rect 40979 26608 41043 26672
rect 40979 26528 41043 26592
rect 40979 26448 41043 26512
rect 40979 26368 41043 26432
rect 40979 26288 41043 26352
rect 40979 26208 41043 26272
rect 40979 26128 41043 26192
rect 40979 26048 41043 26112
rect 40979 25968 41043 26032
rect 40979 25888 41043 25952
rect 40979 25808 41043 25872
rect 40979 25728 41043 25792
rect 40979 25648 41043 25712
rect 40979 25568 41043 25632
rect 40979 25488 41043 25552
rect 40979 25408 41043 25472
rect 40979 25328 41043 25392
rect 40979 25248 41043 25312
rect 40979 25168 41043 25232
rect 40979 25088 41043 25152
rect 40979 25008 41043 25072
rect 40979 24928 41043 24992
rect 40979 24848 41043 24912
rect 40979 24768 41043 24832
rect 40979 24688 41043 24752
rect 40979 24608 41043 24672
rect 40979 24528 41043 24592
rect 40979 24448 41043 24512
rect 40979 24368 41043 24432
rect 40979 24288 41043 24352
rect 40979 24208 41043 24272
rect 40979 24128 41043 24192
rect 40979 24048 41043 24112
rect 40979 23968 41043 24032
rect 40979 23888 41043 23952
rect 40979 23808 41043 23872
rect 40979 23728 41043 23792
rect 40979 23648 41043 23712
rect 40979 23568 41043 23632
rect 40979 23488 41043 23552
rect 40979 23408 41043 23472
rect 40979 23328 41043 23392
rect 40979 23248 41043 23312
rect 40979 23168 41043 23232
rect 40979 23088 41043 23152
rect 40979 23008 41043 23072
rect 40979 22928 41043 22992
rect 40979 22848 41043 22912
rect 40979 22768 41043 22832
rect 40979 22688 41043 22752
rect 40979 22608 41043 22672
rect 40979 22528 41043 22592
rect 40979 22448 41043 22512
rect 40979 22368 41043 22432
rect 40979 22288 41043 22352
rect 40979 22208 41043 22272
rect 40979 22128 41043 22192
rect 47298 28208 47362 28272
rect 47298 28128 47362 28192
rect 47298 28048 47362 28112
rect 47298 27968 47362 28032
rect 47298 27888 47362 27952
rect 47298 27808 47362 27872
rect 47298 27728 47362 27792
rect 47298 27648 47362 27712
rect 47298 27568 47362 27632
rect 47298 27488 47362 27552
rect 47298 27408 47362 27472
rect 47298 27328 47362 27392
rect 47298 27248 47362 27312
rect 47298 27168 47362 27232
rect 47298 27088 47362 27152
rect 47298 27008 47362 27072
rect 47298 26928 47362 26992
rect 47298 26848 47362 26912
rect 47298 26768 47362 26832
rect 47298 26688 47362 26752
rect 47298 26608 47362 26672
rect 47298 26528 47362 26592
rect 47298 26448 47362 26512
rect 47298 26368 47362 26432
rect 47298 26288 47362 26352
rect 47298 26208 47362 26272
rect 47298 26128 47362 26192
rect 47298 26048 47362 26112
rect 47298 25968 47362 26032
rect 47298 25888 47362 25952
rect 47298 25808 47362 25872
rect 47298 25728 47362 25792
rect 47298 25648 47362 25712
rect 47298 25568 47362 25632
rect 47298 25488 47362 25552
rect 47298 25408 47362 25472
rect 47298 25328 47362 25392
rect 47298 25248 47362 25312
rect 47298 25168 47362 25232
rect 47298 25088 47362 25152
rect 47298 25008 47362 25072
rect 47298 24928 47362 24992
rect 47298 24848 47362 24912
rect 47298 24768 47362 24832
rect 47298 24688 47362 24752
rect 47298 24608 47362 24672
rect 47298 24528 47362 24592
rect 47298 24448 47362 24512
rect 47298 24368 47362 24432
rect 47298 24288 47362 24352
rect 47298 24208 47362 24272
rect 47298 24128 47362 24192
rect 47298 24048 47362 24112
rect 47298 23968 47362 24032
rect 47298 23888 47362 23952
rect 47298 23808 47362 23872
rect 47298 23728 47362 23792
rect 47298 23648 47362 23712
rect 47298 23568 47362 23632
rect 47298 23488 47362 23552
rect 47298 23408 47362 23472
rect 47298 23328 47362 23392
rect 47298 23248 47362 23312
rect 47298 23168 47362 23232
rect 47298 23088 47362 23152
rect 47298 23008 47362 23072
rect 47298 22928 47362 22992
rect 47298 22848 47362 22912
rect 47298 22768 47362 22832
rect 47298 22688 47362 22752
rect 47298 22608 47362 22672
rect 47298 22528 47362 22592
rect 47298 22448 47362 22512
rect 47298 22368 47362 22432
rect 47298 22288 47362 22352
rect 47298 22208 47362 22272
rect 47298 22128 47362 22192
rect -41168 21908 -41104 21972
rect -41168 21828 -41104 21892
rect -41168 21748 -41104 21812
rect -41168 21668 -41104 21732
rect -41168 21588 -41104 21652
rect -41168 21508 -41104 21572
rect -41168 21428 -41104 21492
rect -41168 21348 -41104 21412
rect -41168 21268 -41104 21332
rect -41168 21188 -41104 21252
rect -41168 21108 -41104 21172
rect -41168 21028 -41104 21092
rect -41168 20948 -41104 21012
rect -41168 20868 -41104 20932
rect -41168 20788 -41104 20852
rect -41168 20708 -41104 20772
rect -41168 20628 -41104 20692
rect -41168 20548 -41104 20612
rect -41168 20468 -41104 20532
rect -41168 20388 -41104 20452
rect -41168 20308 -41104 20372
rect -41168 20228 -41104 20292
rect -41168 20148 -41104 20212
rect -41168 20068 -41104 20132
rect -41168 19988 -41104 20052
rect -41168 19908 -41104 19972
rect -41168 19828 -41104 19892
rect -41168 19748 -41104 19812
rect -41168 19668 -41104 19732
rect -41168 19588 -41104 19652
rect -41168 19508 -41104 19572
rect -41168 19428 -41104 19492
rect -41168 19348 -41104 19412
rect -41168 19268 -41104 19332
rect -41168 19188 -41104 19252
rect -41168 19108 -41104 19172
rect -41168 19028 -41104 19092
rect -41168 18948 -41104 19012
rect -41168 18868 -41104 18932
rect -41168 18788 -41104 18852
rect -41168 18708 -41104 18772
rect -41168 18628 -41104 18692
rect -41168 18548 -41104 18612
rect -41168 18468 -41104 18532
rect -41168 18388 -41104 18452
rect -41168 18308 -41104 18372
rect -41168 18228 -41104 18292
rect -41168 18148 -41104 18212
rect -41168 18068 -41104 18132
rect -41168 17988 -41104 18052
rect -41168 17908 -41104 17972
rect -41168 17828 -41104 17892
rect -41168 17748 -41104 17812
rect -41168 17668 -41104 17732
rect -41168 17588 -41104 17652
rect -41168 17508 -41104 17572
rect -41168 17428 -41104 17492
rect -41168 17348 -41104 17412
rect -41168 17268 -41104 17332
rect -41168 17188 -41104 17252
rect -41168 17108 -41104 17172
rect -41168 17028 -41104 17092
rect -41168 16948 -41104 17012
rect -41168 16868 -41104 16932
rect -41168 16788 -41104 16852
rect -41168 16708 -41104 16772
rect -41168 16628 -41104 16692
rect -41168 16548 -41104 16612
rect -41168 16468 -41104 16532
rect -41168 16388 -41104 16452
rect -41168 16308 -41104 16372
rect -41168 16228 -41104 16292
rect -41168 16148 -41104 16212
rect -41168 16068 -41104 16132
rect -41168 15988 -41104 16052
rect -41168 15908 -41104 15972
rect -41168 15828 -41104 15892
rect -34849 21908 -34785 21972
rect -34849 21828 -34785 21892
rect -34849 21748 -34785 21812
rect -34849 21668 -34785 21732
rect -34849 21588 -34785 21652
rect -34849 21508 -34785 21572
rect -34849 21428 -34785 21492
rect -34849 21348 -34785 21412
rect -34849 21268 -34785 21332
rect -34849 21188 -34785 21252
rect -34849 21108 -34785 21172
rect -34849 21028 -34785 21092
rect -34849 20948 -34785 21012
rect -34849 20868 -34785 20932
rect -34849 20788 -34785 20852
rect -34849 20708 -34785 20772
rect -34849 20628 -34785 20692
rect -34849 20548 -34785 20612
rect -34849 20468 -34785 20532
rect -34849 20388 -34785 20452
rect -34849 20308 -34785 20372
rect -34849 20228 -34785 20292
rect -34849 20148 -34785 20212
rect -34849 20068 -34785 20132
rect -34849 19988 -34785 20052
rect -34849 19908 -34785 19972
rect -34849 19828 -34785 19892
rect -34849 19748 -34785 19812
rect -34849 19668 -34785 19732
rect -34849 19588 -34785 19652
rect -34849 19508 -34785 19572
rect -34849 19428 -34785 19492
rect -34849 19348 -34785 19412
rect -34849 19268 -34785 19332
rect -34849 19188 -34785 19252
rect -34849 19108 -34785 19172
rect -34849 19028 -34785 19092
rect -34849 18948 -34785 19012
rect -34849 18868 -34785 18932
rect -34849 18788 -34785 18852
rect -34849 18708 -34785 18772
rect -34849 18628 -34785 18692
rect -34849 18548 -34785 18612
rect -34849 18468 -34785 18532
rect -34849 18388 -34785 18452
rect -34849 18308 -34785 18372
rect -34849 18228 -34785 18292
rect -34849 18148 -34785 18212
rect -34849 18068 -34785 18132
rect -34849 17988 -34785 18052
rect -34849 17908 -34785 17972
rect -34849 17828 -34785 17892
rect -34849 17748 -34785 17812
rect -34849 17668 -34785 17732
rect -34849 17588 -34785 17652
rect -34849 17508 -34785 17572
rect -34849 17428 -34785 17492
rect -34849 17348 -34785 17412
rect -34849 17268 -34785 17332
rect -34849 17188 -34785 17252
rect -34849 17108 -34785 17172
rect -34849 17028 -34785 17092
rect -34849 16948 -34785 17012
rect -34849 16868 -34785 16932
rect -34849 16788 -34785 16852
rect -34849 16708 -34785 16772
rect -34849 16628 -34785 16692
rect -34849 16548 -34785 16612
rect -34849 16468 -34785 16532
rect -34849 16388 -34785 16452
rect -34849 16308 -34785 16372
rect -34849 16228 -34785 16292
rect -34849 16148 -34785 16212
rect -34849 16068 -34785 16132
rect -34849 15988 -34785 16052
rect -34849 15908 -34785 15972
rect -34849 15828 -34785 15892
rect -28530 21908 -28466 21972
rect -28530 21828 -28466 21892
rect -28530 21748 -28466 21812
rect -28530 21668 -28466 21732
rect -28530 21588 -28466 21652
rect -28530 21508 -28466 21572
rect -28530 21428 -28466 21492
rect -28530 21348 -28466 21412
rect -28530 21268 -28466 21332
rect -28530 21188 -28466 21252
rect -28530 21108 -28466 21172
rect -28530 21028 -28466 21092
rect -28530 20948 -28466 21012
rect -28530 20868 -28466 20932
rect -28530 20788 -28466 20852
rect -28530 20708 -28466 20772
rect -28530 20628 -28466 20692
rect -28530 20548 -28466 20612
rect -28530 20468 -28466 20532
rect -28530 20388 -28466 20452
rect -28530 20308 -28466 20372
rect -28530 20228 -28466 20292
rect -28530 20148 -28466 20212
rect -28530 20068 -28466 20132
rect -28530 19988 -28466 20052
rect -28530 19908 -28466 19972
rect -28530 19828 -28466 19892
rect -28530 19748 -28466 19812
rect -28530 19668 -28466 19732
rect -28530 19588 -28466 19652
rect -28530 19508 -28466 19572
rect -28530 19428 -28466 19492
rect -28530 19348 -28466 19412
rect -28530 19268 -28466 19332
rect -28530 19188 -28466 19252
rect -28530 19108 -28466 19172
rect -28530 19028 -28466 19092
rect -28530 18948 -28466 19012
rect -28530 18868 -28466 18932
rect -28530 18788 -28466 18852
rect -28530 18708 -28466 18772
rect -28530 18628 -28466 18692
rect -28530 18548 -28466 18612
rect -28530 18468 -28466 18532
rect -28530 18388 -28466 18452
rect -28530 18308 -28466 18372
rect -28530 18228 -28466 18292
rect -28530 18148 -28466 18212
rect -28530 18068 -28466 18132
rect -28530 17988 -28466 18052
rect -28530 17908 -28466 17972
rect -28530 17828 -28466 17892
rect -28530 17748 -28466 17812
rect -28530 17668 -28466 17732
rect -28530 17588 -28466 17652
rect -28530 17508 -28466 17572
rect -28530 17428 -28466 17492
rect -28530 17348 -28466 17412
rect -28530 17268 -28466 17332
rect -28530 17188 -28466 17252
rect -28530 17108 -28466 17172
rect -28530 17028 -28466 17092
rect -28530 16948 -28466 17012
rect -28530 16868 -28466 16932
rect -28530 16788 -28466 16852
rect -28530 16708 -28466 16772
rect -28530 16628 -28466 16692
rect -28530 16548 -28466 16612
rect -28530 16468 -28466 16532
rect -28530 16388 -28466 16452
rect -28530 16308 -28466 16372
rect -28530 16228 -28466 16292
rect -28530 16148 -28466 16212
rect -28530 16068 -28466 16132
rect -28530 15988 -28466 16052
rect -28530 15908 -28466 15972
rect -28530 15828 -28466 15892
rect -22211 21908 -22147 21972
rect -22211 21828 -22147 21892
rect -22211 21748 -22147 21812
rect -22211 21668 -22147 21732
rect -22211 21588 -22147 21652
rect -22211 21508 -22147 21572
rect -22211 21428 -22147 21492
rect -22211 21348 -22147 21412
rect -22211 21268 -22147 21332
rect -22211 21188 -22147 21252
rect -22211 21108 -22147 21172
rect -22211 21028 -22147 21092
rect -22211 20948 -22147 21012
rect -22211 20868 -22147 20932
rect -22211 20788 -22147 20852
rect -22211 20708 -22147 20772
rect -22211 20628 -22147 20692
rect -22211 20548 -22147 20612
rect -22211 20468 -22147 20532
rect -22211 20388 -22147 20452
rect -22211 20308 -22147 20372
rect -22211 20228 -22147 20292
rect -22211 20148 -22147 20212
rect -22211 20068 -22147 20132
rect -22211 19988 -22147 20052
rect -22211 19908 -22147 19972
rect -22211 19828 -22147 19892
rect -22211 19748 -22147 19812
rect -22211 19668 -22147 19732
rect -22211 19588 -22147 19652
rect -22211 19508 -22147 19572
rect -22211 19428 -22147 19492
rect -22211 19348 -22147 19412
rect -22211 19268 -22147 19332
rect -22211 19188 -22147 19252
rect -22211 19108 -22147 19172
rect -22211 19028 -22147 19092
rect -22211 18948 -22147 19012
rect -22211 18868 -22147 18932
rect -22211 18788 -22147 18852
rect -22211 18708 -22147 18772
rect -22211 18628 -22147 18692
rect -22211 18548 -22147 18612
rect -22211 18468 -22147 18532
rect -22211 18388 -22147 18452
rect -22211 18308 -22147 18372
rect -22211 18228 -22147 18292
rect -22211 18148 -22147 18212
rect -22211 18068 -22147 18132
rect -22211 17988 -22147 18052
rect -22211 17908 -22147 17972
rect -22211 17828 -22147 17892
rect -22211 17748 -22147 17812
rect -22211 17668 -22147 17732
rect -22211 17588 -22147 17652
rect -22211 17508 -22147 17572
rect -22211 17428 -22147 17492
rect -22211 17348 -22147 17412
rect -22211 17268 -22147 17332
rect -22211 17188 -22147 17252
rect -22211 17108 -22147 17172
rect -22211 17028 -22147 17092
rect -22211 16948 -22147 17012
rect -22211 16868 -22147 16932
rect -22211 16788 -22147 16852
rect -22211 16708 -22147 16772
rect -22211 16628 -22147 16692
rect -22211 16548 -22147 16612
rect -22211 16468 -22147 16532
rect -22211 16388 -22147 16452
rect -22211 16308 -22147 16372
rect -22211 16228 -22147 16292
rect -22211 16148 -22147 16212
rect -22211 16068 -22147 16132
rect -22211 15988 -22147 16052
rect -22211 15908 -22147 15972
rect -22211 15828 -22147 15892
rect -15892 21908 -15828 21972
rect -15892 21828 -15828 21892
rect -15892 21748 -15828 21812
rect -15892 21668 -15828 21732
rect -15892 21588 -15828 21652
rect -15892 21508 -15828 21572
rect -15892 21428 -15828 21492
rect -15892 21348 -15828 21412
rect -15892 21268 -15828 21332
rect -15892 21188 -15828 21252
rect -15892 21108 -15828 21172
rect -15892 21028 -15828 21092
rect -15892 20948 -15828 21012
rect -15892 20868 -15828 20932
rect -15892 20788 -15828 20852
rect -15892 20708 -15828 20772
rect -15892 20628 -15828 20692
rect -15892 20548 -15828 20612
rect -15892 20468 -15828 20532
rect -15892 20388 -15828 20452
rect -15892 20308 -15828 20372
rect -15892 20228 -15828 20292
rect -15892 20148 -15828 20212
rect -15892 20068 -15828 20132
rect -15892 19988 -15828 20052
rect -15892 19908 -15828 19972
rect -15892 19828 -15828 19892
rect -15892 19748 -15828 19812
rect -15892 19668 -15828 19732
rect -15892 19588 -15828 19652
rect -15892 19508 -15828 19572
rect -15892 19428 -15828 19492
rect -15892 19348 -15828 19412
rect -15892 19268 -15828 19332
rect -15892 19188 -15828 19252
rect -15892 19108 -15828 19172
rect -15892 19028 -15828 19092
rect -15892 18948 -15828 19012
rect -15892 18868 -15828 18932
rect -15892 18788 -15828 18852
rect -15892 18708 -15828 18772
rect -15892 18628 -15828 18692
rect -15892 18548 -15828 18612
rect -15892 18468 -15828 18532
rect -15892 18388 -15828 18452
rect -15892 18308 -15828 18372
rect -15892 18228 -15828 18292
rect -15892 18148 -15828 18212
rect -15892 18068 -15828 18132
rect -15892 17988 -15828 18052
rect -15892 17908 -15828 17972
rect -15892 17828 -15828 17892
rect -15892 17748 -15828 17812
rect -15892 17668 -15828 17732
rect -15892 17588 -15828 17652
rect -15892 17508 -15828 17572
rect -15892 17428 -15828 17492
rect -15892 17348 -15828 17412
rect -15892 17268 -15828 17332
rect -15892 17188 -15828 17252
rect -15892 17108 -15828 17172
rect -15892 17028 -15828 17092
rect -15892 16948 -15828 17012
rect -15892 16868 -15828 16932
rect -15892 16788 -15828 16852
rect -15892 16708 -15828 16772
rect -15892 16628 -15828 16692
rect -15892 16548 -15828 16612
rect -15892 16468 -15828 16532
rect -15892 16388 -15828 16452
rect -15892 16308 -15828 16372
rect -15892 16228 -15828 16292
rect -15892 16148 -15828 16212
rect -15892 16068 -15828 16132
rect -15892 15988 -15828 16052
rect -15892 15908 -15828 15972
rect -15892 15828 -15828 15892
rect -9573 21908 -9509 21972
rect -9573 21828 -9509 21892
rect -9573 21748 -9509 21812
rect -9573 21668 -9509 21732
rect -9573 21588 -9509 21652
rect -9573 21508 -9509 21572
rect -9573 21428 -9509 21492
rect -9573 21348 -9509 21412
rect -9573 21268 -9509 21332
rect -9573 21188 -9509 21252
rect -9573 21108 -9509 21172
rect -9573 21028 -9509 21092
rect -9573 20948 -9509 21012
rect -9573 20868 -9509 20932
rect -9573 20788 -9509 20852
rect -9573 20708 -9509 20772
rect -9573 20628 -9509 20692
rect -9573 20548 -9509 20612
rect -9573 20468 -9509 20532
rect -9573 20388 -9509 20452
rect -9573 20308 -9509 20372
rect -9573 20228 -9509 20292
rect -9573 20148 -9509 20212
rect -9573 20068 -9509 20132
rect -9573 19988 -9509 20052
rect -9573 19908 -9509 19972
rect -9573 19828 -9509 19892
rect -9573 19748 -9509 19812
rect -9573 19668 -9509 19732
rect -9573 19588 -9509 19652
rect -9573 19508 -9509 19572
rect -9573 19428 -9509 19492
rect -9573 19348 -9509 19412
rect -9573 19268 -9509 19332
rect -9573 19188 -9509 19252
rect -9573 19108 -9509 19172
rect -9573 19028 -9509 19092
rect -9573 18948 -9509 19012
rect -9573 18868 -9509 18932
rect -9573 18788 -9509 18852
rect -9573 18708 -9509 18772
rect -9573 18628 -9509 18692
rect -9573 18548 -9509 18612
rect -9573 18468 -9509 18532
rect -9573 18388 -9509 18452
rect -9573 18308 -9509 18372
rect -9573 18228 -9509 18292
rect -9573 18148 -9509 18212
rect -9573 18068 -9509 18132
rect -9573 17988 -9509 18052
rect -9573 17908 -9509 17972
rect -9573 17828 -9509 17892
rect -9573 17748 -9509 17812
rect -9573 17668 -9509 17732
rect -9573 17588 -9509 17652
rect -9573 17508 -9509 17572
rect -9573 17428 -9509 17492
rect -9573 17348 -9509 17412
rect -9573 17268 -9509 17332
rect -9573 17188 -9509 17252
rect -9573 17108 -9509 17172
rect -9573 17028 -9509 17092
rect -9573 16948 -9509 17012
rect -9573 16868 -9509 16932
rect -9573 16788 -9509 16852
rect -9573 16708 -9509 16772
rect -9573 16628 -9509 16692
rect -9573 16548 -9509 16612
rect -9573 16468 -9509 16532
rect -9573 16388 -9509 16452
rect -9573 16308 -9509 16372
rect -9573 16228 -9509 16292
rect -9573 16148 -9509 16212
rect -9573 16068 -9509 16132
rect -9573 15988 -9509 16052
rect -9573 15908 -9509 15972
rect -9573 15828 -9509 15892
rect -3254 21908 -3190 21972
rect -3254 21828 -3190 21892
rect -3254 21748 -3190 21812
rect -3254 21668 -3190 21732
rect -3254 21588 -3190 21652
rect -3254 21508 -3190 21572
rect -3254 21428 -3190 21492
rect -3254 21348 -3190 21412
rect -3254 21268 -3190 21332
rect -3254 21188 -3190 21252
rect -3254 21108 -3190 21172
rect -3254 21028 -3190 21092
rect -3254 20948 -3190 21012
rect -3254 20868 -3190 20932
rect -3254 20788 -3190 20852
rect -3254 20708 -3190 20772
rect -3254 20628 -3190 20692
rect -3254 20548 -3190 20612
rect -3254 20468 -3190 20532
rect -3254 20388 -3190 20452
rect -3254 20308 -3190 20372
rect -3254 20228 -3190 20292
rect -3254 20148 -3190 20212
rect -3254 20068 -3190 20132
rect -3254 19988 -3190 20052
rect -3254 19908 -3190 19972
rect -3254 19828 -3190 19892
rect -3254 19748 -3190 19812
rect -3254 19668 -3190 19732
rect -3254 19588 -3190 19652
rect -3254 19508 -3190 19572
rect -3254 19428 -3190 19492
rect -3254 19348 -3190 19412
rect -3254 19268 -3190 19332
rect -3254 19188 -3190 19252
rect -3254 19108 -3190 19172
rect -3254 19028 -3190 19092
rect -3254 18948 -3190 19012
rect -3254 18868 -3190 18932
rect -3254 18788 -3190 18852
rect -3254 18708 -3190 18772
rect -3254 18628 -3190 18692
rect -3254 18548 -3190 18612
rect -3254 18468 -3190 18532
rect -3254 18388 -3190 18452
rect -3254 18308 -3190 18372
rect -3254 18228 -3190 18292
rect -3254 18148 -3190 18212
rect -3254 18068 -3190 18132
rect -3254 17988 -3190 18052
rect -3254 17908 -3190 17972
rect -3254 17828 -3190 17892
rect -3254 17748 -3190 17812
rect -3254 17668 -3190 17732
rect -3254 17588 -3190 17652
rect -3254 17508 -3190 17572
rect -3254 17428 -3190 17492
rect -3254 17348 -3190 17412
rect -3254 17268 -3190 17332
rect -3254 17188 -3190 17252
rect -3254 17108 -3190 17172
rect -3254 17028 -3190 17092
rect -3254 16948 -3190 17012
rect -3254 16868 -3190 16932
rect -3254 16788 -3190 16852
rect -3254 16708 -3190 16772
rect -3254 16628 -3190 16692
rect -3254 16548 -3190 16612
rect -3254 16468 -3190 16532
rect -3254 16388 -3190 16452
rect -3254 16308 -3190 16372
rect -3254 16228 -3190 16292
rect -3254 16148 -3190 16212
rect -3254 16068 -3190 16132
rect -3254 15988 -3190 16052
rect -3254 15908 -3190 15972
rect -3254 15828 -3190 15892
rect 3065 21908 3129 21972
rect 3065 21828 3129 21892
rect 3065 21748 3129 21812
rect 3065 21668 3129 21732
rect 3065 21588 3129 21652
rect 3065 21508 3129 21572
rect 3065 21428 3129 21492
rect 3065 21348 3129 21412
rect 3065 21268 3129 21332
rect 3065 21188 3129 21252
rect 3065 21108 3129 21172
rect 3065 21028 3129 21092
rect 3065 20948 3129 21012
rect 3065 20868 3129 20932
rect 3065 20788 3129 20852
rect 3065 20708 3129 20772
rect 3065 20628 3129 20692
rect 3065 20548 3129 20612
rect 3065 20468 3129 20532
rect 3065 20388 3129 20452
rect 3065 20308 3129 20372
rect 3065 20228 3129 20292
rect 3065 20148 3129 20212
rect 3065 20068 3129 20132
rect 3065 19988 3129 20052
rect 3065 19908 3129 19972
rect 3065 19828 3129 19892
rect 3065 19748 3129 19812
rect 3065 19668 3129 19732
rect 3065 19588 3129 19652
rect 3065 19508 3129 19572
rect 3065 19428 3129 19492
rect 3065 19348 3129 19412
rect 3065 19268 3129 19332
rect 3065 19188 3129 19252
rect 3065 19108 3129 19172
rect 3065 19028 3129 19092
rect 3065 18948 3129 19012
rect 3065 18868 3129 18932
rect 3065 18788 3129 18852
rect 3065 18708 3129 18772
rect 3065 18628 3129 18692
rect 3065 18548 3129 18612
rect 3065 18468 3129 18532
rect 3065 18388 3129 18452
rect 3065 18308 3129 18372
rect 3065 18228 3129 18292
rect 3065 18148 3129 18212
rect 3065 18068 3129 18132
rect 3065 17988 3129 18052
rect 3065 17908 3129 17972
rect 3065 17828 3129 17892
rect 3065 17748 3129 17812
rect 3065 17668 3129 17732
rect 3065 17588 3129 17652
rect 3065 17508 3129 17572
rect 3065 17428 3129 17492
rect 3065 17348 3129 17412
rect 3065 17268 3129 17332
rect 3065 17188 3129 17252
rect 3065 17108 3129 17172
rect 3065 17028 3129 17092
rect 3065 16948 3129 17012
rect 3065 16868 3129 16932
rect 3065 16788 3129 16852
rect 3065 16708 3129 16772
rect 3065 16628 3129 16692
rect 3065 16548 3129 16612
rect 3065 16468 3129 16532
rect 3065 16388 3129 16452
rect 3065 16308 3129 16372
rect 3065 16228 3129 16292
rect 3065 16148 3129 16212
rect 3065 16068 3129 16132
rect 3065 15988 3129 16052
rect 3065 15908 3129 15972
rect 3065 15828 3129 15892
rect 9384 21908 9448 21972
rect 9384 21828 9448 21892
rect 9384 21748 9448 21812
rect 9384 21668 9448 21732
rect 9384 21588 9448 21652
rect 9384 21508 9448 21572
rect 9384 21428 9448 21492
rect 9384 21348 9448 21412
rect 9384 21268 9448 21332
rect 9384 21188 9448 21252
rect 9384 21108 9448 21172
rect 9384 21028 9448 21092
rect 9384 20948 9448 21012
rect 9384 20868 9448 20932
rect 9384 20788 9448 20852
rect 9384 20708 9448 20772
rect 9384 20628 9448 20692
rect 9384 20548 9448 20612
rect 9384 20468 9448 20532
rect 9384 20388 9448 20452
rect 9384 20308 9448 20372
rect 9384 20228 9448 20292
rect 9384 20148 9448 20212
rect 9384 20068 9448 20132
rect 9384 19988 9448 20052
rect 9384 19908 9448 19972
rect 9384 19828 9448 19892
rect 9384 19748 9448 19812
rect 9384 19668 9448 19732
rect 9384 19588 9448 19652
rect 9384 19508 9448 19572
rect 9384 19428 9448 19492
rect 9384 19348 9448 19412
rect 9384 19268 9448 19332
rect 9384 19188 9448 19252
rect 9384 19108 9448 19172
rect 9384 19028 9448 19092
rect 9384 18948 9448 19012
rect 9384 18868 9448 18932
rect 9384 18788 9448 18852
rect 9384 18708 9448 18772
rect 9384 18628 9448 18692
rect 9384 18548 9448 18612
rect 9384 18468 9448 18532
rect 9384 18388 9448 18452
rect 9384 18308 9448 18372
rect 9384 18228 9448 18292
rect 9384 18148 9448 18212
rect 9384 18068 9448 18132
rect 9384 17988 9448 18052
rect 9384 17908 9448 17972
rect 9384 17828 9448 17892
rect 9384 17748 9448 17812
rect 9384 17668 9448 17732
rect 9384 17588 9448 17652
rect 9384 17508 9448 17572
rect 9384 17428 9448 17492
rect 9384 17348 9448 17412
rect 9384 17268 9448 17332
rect 9384 17188 9448 17252
rect 9384 17108 9448 17172
rect 9384 17028 9448 17092
rect 9384 16948 9448 17012
rect 9384 16868 9448 16932
rect 9384 16788 9448 16852
rect 9384 16708 9448 16772
rect 9384 16628 9448 16692
rect 9384 16548 9448 16612
rect 9384 16468 9448 16532
rect 9384 16388 9448 16452
rect 9384 16308 9448 16372
rect 9384 16228 9448 16292
rect 9384 16148 9448 16212
rect 9384 16068 9448 16132
rect 9384 15988 9448 16052
rect 9384 15908 9448 15972
rect 9384 15828 9448 15892
rect 15703 21908 15767 21972
rect 15703 21828 15767 21892
rect 15703 21748 15767 21812
rect 15703 21668 15767 21732
rect 15703 21588 15767 21652
rect 15703 21508 15767 21572
rect 15703 21428 15767 21492
rect 15703 21348 15767 21412
rect 15703 21268 15767 21332
rect 15703 21188 15767 21252
rect 15703 21108 15767 21172
rect 15703 21028 15767 21092
rect 15703 20948 15767 21012
rect 15703 20868 15767 20932
rect 15703 20788 15767 20852
rect 15703 20708 15767 20772
rect 15703 20628 15767 20692
rect 15703 20548 15767 20612
rect 15703 20468 15767 20532
rect 15703 20388 15767 20452
rect 15703 20308 15767 20372
rect 15703 20228 15767 20292
rect 15703 20148 15767 20212
rect 15703 20068 15767 20132
rect 15703 19988 15767 20052
rect 15703 19908 15767 19972
rect 15703 19828 15767 19892
rect 15703 19748 15767 19812
rect 15703 19668 15767 19732
rect 15703 19588 15767 19652
rect 15703 19508 15767 19572
rect 15703 19428 15767 19492
rect 15703 19348 15767 19412
rect 15703 19268 15767 19332
rect 15703 19188 15767 19252
rect 15703 19108 15767 19172
rect 15703 19028 15767 19092
rect 15703 18948 15767 19012
rect 15703 18868 15767 18932
rect 15703 18788 15767 18852
rect 15703 18708 15767 18772
rect 15703 18628 15767 18692
rect 15703 18548 15767 18612
rect 15703 18468 15767 18532
rect 15703 18388 15767 18452
rect 15703 18308 15767 18372
rect 15703 18228 15767 18292
rect 15703 18148 15767 18212
rect 15703 18068 15767 18132
rect 15703 17988 15767 18052
rect 15703 17908 15767 17972
rect 15703 17828 15767 17892
rect 15703 17748 15767 17812
rect 15703 17668 15767 17732
rect 15703 17588 15767 17652
rect 15703 17508 15767 17572
rect 15703 17428 15767 17492
rect 15703 17348 15767 17412
rect 15703 17268 15767 17332
rect 15703 17188 15767 17252
rect 15703 17108 15767 17172
rect 15703 17028 15767 17092
rect 15703 16948 15767 17012
rect 15703 16868 15767 16932
rect 15703 16788 15767 16852
rect 15703 16708 15767 16772
rect 15703 16628 15767 16692
rect 15703 16548 15767 16612
rect 15703 16468 15767 16532
rect 15703 16388 15767 16452
rect 15703 16308 15767 16372
rect 15703 16228 15767 16292
rect 15703 16148 15767 16212
rect 15703 16068 15767 16132
rect 15703 15988 15767 16052
rect 15703 15908 15767 15972
rect 15703 15828 15767 15892
rect 22022 21908 22086 21972
rect 22022 21828 22086 21892
rect 22022 21748 22086 21812
rect 22022 21668 22086 21732
rect 22022 21588 22086 21652
rect 22022 21508 22086 21572
rect 22022 21428 22086 21492
rect 22022 21348 22086 21412
rect 22022 21268 22086 21332
rect 22022 21188 22086 21252
rect 22022 21108 22086 21172
rect 22022 21028 22086 21092
rect 22022 20948 22086 21012
rect 22022 20868 22086 20932
rect 22022 20788 22086 20852
rect 22022 20708 22086 20772
rect 22022 20628 22086 20692
rect 22022 20548 22086 20612
rect 22022 20468 22086 20532
rect 22022 20388 22086 20452
rect 22022 20308 22086 20372
rect 22022 20228 22086 20292
rect 22022 20148 22086 20212
rect 22022 20068 22086 20132
rect 22022 19988 22086 20052
rect 22022 19908 22086 19972
rect 22022 19828 22086 19892
rect 22022 19748 22086 19812
rect 22022 19668 22086 19732
rect 22022 19588 22086 19652
rect 22022 19508 22086 19572
rect 22022 19428 22086 19492
rect 22022 19348 22086 19412
rect 22022 19268 22086 19332
rect 22022 19188 22086 19252
rect 22022 19108 22086 19172
rect 22022 19028 22086 19092
rect 22022 18948 22086 19012
rect 22022 18868 22086 18932
rect 22022 18788 22086 18852
rect 22022 18708 22086 18772
rect 22022 18628 22086 18692
rect 22022 18548 22086 18612
rect 22022 18468 22086 18532
rect 22022 18388 22086 18452
rect 22022 18308 22086 18372
rect 22022 18228 22086 18292
rect 22022 18148 22086 18212
rect 22022 18068 22086 18132
rect 22022 17988 22086 18052
rect 22022 17908 22086 17972
rect 22022 17828 22086 17892
rect 22022 17748 22086 17812
rect 22022 17668 22086 17732
rect 22022 17588 22086 17652
rect 22022 17508 22086 17572
rect 22022 17428 22086 17492
rect 22022 17348 22086 17412
rect 22022 17268 22086 17332
rect 22022 17188 22086 17252
rect 22022 17108 22086 17172
rect 22022 17028 22086 17092
rect 22022 16948 22086 17012
rect 22022 16868 22086 16932
rect 22022 16788 22086 16852
rect 22022 16708 22086 16772
rect 22022 16628 22086 16692
rect 22022 16548 22086 16612
rect 22022 16468 22086 16532
rect 22022 16388 22086 16452
rect 22022 16308 22086 16372
rect 22022 16228 22086 16292
rect 22022 16148 22086 16212
rect 22022 16068 22086 16132
rect 22022 15988 22086 16052
rect 22022 15908 22086 15972
rect 22022 15828 22086 15892
rect 28341 21908 28405 21972
rect 28341 21828 28405 21892
rect 28341 21748 28405 21812
rect 28341 21668 28405 21732
rect 28341 21588 28405 21652
rect 28341 21508 28405 21572
rect 28341 21428 28405 21492
rect 28341 21348 28405 21412
rect 28341 21268 28405 21332
rect 28341 21188 28405 21252
rect 28341 21108 28405 21172
rect 28341 21028 28405 21092
rect 28341 20948 28405 21012
rect 28341 20868 28405 20932
rect 28341 20788 28405 20852
rect 28341 20708 28405 20772
rect 28341 20628 28405 20692
rect 28341 20548 28405 20612
rect 28341 20468 28405 20532
rect 28341 20388 28405 20452
rect 28341 20308 28405 20372
rect 28341 20228 28405 20292
rect 28341 20148 28405 20212
rect 28341 20068 28405 20132
rect 28341 19988 28405 20052
rect 28341 19908 28405 19972
rect 28341 19828 28405 19892
rect 28341 19748 28405 19812
rect 28341 19668 28405 19732
rect 28341 19588 28405 19652
rect 28341 19508 28405 19572
rect 28341 19428 28405 19492
rect 28341 19348 28405 19412
rect 28341 19268 28405 19332
rect 28341 19188 28405 19252
rect 28341 19108 28405 19172
rect 28341 19028 28405 19092
rect 28341 18948 28405 19012
rect 28341 18868 28405 18932
rect 28341 18788 28405 18852
rect 28341 18708 28405 18772
rect 28341 18628 28405 18692
rect 28341 18548 28405 18612
rect 28341 18468 28405 18532
rect 28341 18388 28405 18452
rect 28341 18308 28405 18372
rect 28341 18228 28405 18292
rect 28341 18148 28405 18212
rect 28341 18068 28405 18132
rect 28341 17988 28405 18052
rect 28341 17908 28405 17972
rect 28341 17828 28405 17892
rect 28341 17748 28405 17812
rect 28341 17668 28405 17732
rect 28341 17588 28405 17652
rect 28341 17508 28405 17572
rect 28341 17428 28405 17492
rect 28341 17348 28405 17412
rect 28341 17268 28405 17332
rect 28341 17188 28405 17252
rect 28341 17108 28405 17172
rect 28341 17028 28405 17092
rect 28341 16948 28405 17012
rect 28341 16868 28405 16932
rect 28341 16788 28405 16852
rect 28341 16708 28405 16772
rect 28341 16628 28405 16692
rect 28341 16548 28405 16612
rect 28341 16468 28405 16532
rect 28341 16388 28405 16452
rect 28341 16308 28405 16372
rect 28341 16228 28405 16292
rect 28341 16148 28405 16212
rect 28341 16068 28405 16132
rect 28341 15988 28405 16052
rect 28341 15908 28405 15972
rect 28341 15828 28405 15892
rect 34660 21908 34724 21972
rect 34660 21828 34724 21892
rect 34660 21748 34724 21812
rect 34660 21668 34724 21732
rect 34660 21588 34724 21652
rect 34660 21508 34724 21572
rect 34660 21428 34724 21492
rect 34660 21348 34724 21412
rect 34660 21268 34724 21332
rect 34660 21188 34724 21252
rect 34660 21108 34724 21172
rect 34660 21028 34724 21092
rect 34660 20948 34724 21012
rect 34660 20868 34724 20932
rect 34660 20788 34724 20852
rect 34660 20708 34724 20772
rect 34660 20628 34724 20692
rect 34660 20548 34724 20612
rect 34660 20468 34724 20532
rect 34660 20388 34724 20452
rect 34660 20308 34724 20372
rect 34660 20228 34724 20292
rect 34660 20148 34724 20212
rect 34660 20068 34724 20132
rect 34660 19988 34724 20052
rect 34660 19908 34724 19972
rect 34660 19828 34724 19892
rect 34660 19748 34724 19812
rect 34660 19668 34724 19732
rect 34660 19588 34724 19652
rect 34660 19508 34724 19572
rect 34660 19428 34724 19492
rect 34660 19348 34724 19412
rect 34660 19268 34724 19332
rect 34660 19188 34724 19252
rect 34660 19108 34724 19172
rect 34660 19028 34724 19092
rect 34660 18948 34724 19012
rect 34660 18868 34724 18932
rect 34660 18788 34724 18852
rect 34660 18708 34724 18772
rect 34660 18628 34724 18692
rect 34660 18548 34724 18612
rect 34660 18468 34724 18532
rect 34660 18388 34724 18452
rect 34660 18308 34724 18372
rect 34660 18228 34724 18292
rect 34660 18148 34724 18212
rect 34660 18068 34724 18132
rect 34660 17988 34724 18052
rect 34660 17908 34724 17972
rect 34660 17828 34724 17892
rect 34660 17748 34724 17812
rect 34660 17668 34724 17732
rect 34660 17588 34724 17652
rect 34660 17508 34724 17572
rect 34660 17428 34724 17492
rect 34660 17348 34724 17412
rect 34660 17268 34724 17332
rect 34660 17188 34724 17252
rect 34660 17108 34724 17172
rect 34660 17028 34724 17092
rect 34660 16948 34724 17012
rect 34660 16868 34724 16932
rect 34660 16788 34724 16852
rect 34660 16708 34724 16772
rect 34660 16628 34724 16692
rect 34660 16548 34724 16612
rect 34660 16468 34724 16532
rect 34660 16388 34724 16452
rect 34660 16308 34724 16372
rect 34660 16228 34724 16292
rect 34660 16148 34724 16212
rect 34660 16068 34724 16132
rect 34660 15988 34724 16052
rect 34660 15908 34724 15972
rect 34660 15828 34724 15892
rect 40979 21908 41043 21972
rect 40979 21828 41043 21892
rect 40979 21748 41043 21812
rect 40979 21668 41043 21732
rect 40979 21588 41043 21652
rect 40979 21508 41043 21572
rect 40979 21428 41043 21492
rect 40979 21348 41043 21412
rect 40979 21268 41043 21332
rect 40979 21188 41043 21252
rect 40979 21108 41043 21172
rect 40979 21028 41043 21092
rect 40979 20948 41043 21012
rect 40979 20868 41043 20932
rect 40979 20788 41043 20852
rect 40979 20708 41043 20772
rect 40979 20628 41043 20692
rect 40979 20548 41043 20612
rect 40979 20468 41043 20532
rect 40979 20388 41043 20452
rect 40979 20308 41043 20372
rect 40979 20228 41043 20292
rect 40979 20148 41043 20212
rect 40979 20068 41043 20132
rect 40979 19988 41043 20052
rect 40979 19908 41043 19972
rect 40979 19828 41043 19892
rect 40979 19748 41043 19812
rect 40979 19668 41043 19732
rect 40979 19588 41043 19652
rect 40979 19508 41043 19572
rect 40979 19428 41043 19492
rect 40979 19348 41043 19412
rect 40979 19268 41043 19332
rect 40979 19188 41043 19252
rect 40979 19108 41043 19172
rect 40979 19028 41043 19092
rect 40979 18948 41043 19012
rect 40979 18868 41043 18932
rect 40979 18788 41043 18852
rect 40979 18708 41043 18772
rect 40979 18628 41043 18692
rect 40979 18548 41043 18612
rect 40979 18468 41043 18532
rect 40979 18388 41043 18452
rect 40979 18308 41043 18372
rect 40979 18228 41043 18292
rect 40979 18148 41043 18212
rect 40979 18068 41043 18132
rect 40979 17988 41043 18052
rect 40979 17908 41043 17972
rect 40979 17828 41043 17892
rect 40979 17748 41043 17812
rect 40979 17668 41043 17732
rect 40979 17588 41043 17652
rect 40979 17508 41043 17572
rect 40979 17428 41043 17492
rect 40979 17348 41043 17412
rect 40979 17268 41043 17332
rect 40979 17188 41043 17252
rect 40979 17108 41043 17172
rect 40979 17028 41043 17092
rect 40979 16948 41043 17012
rect 40979 16868 41043 16932
rect 40979 16788 41043 16852
rect 40979 16708 41043 16772
rect 40979 16628 41043 16692
rect 40979 16548 41043 16612
rect 40979 16468 41043 16532
rect 40979 16388 41043 16452
rect 40979 16308 41043 16372
rect 40979 16228 41043 16292
rect 40979 16148 41043 16212
rect 40979 16068 41043 16132
rect 40979 15988 41043 16052
rect 40979 15908 41043 15972
rect 40979 15828 41043 15892
rect 47298 21908 47362 21972
rect 47298 21828 47362 21892
rect 47298 21748 47362 21812
rect 47298 21668 47362 21732
rect 47298 21588 47362 21652
rect 47298 21508 47362 21572
rect 47298 21428 47362 21492
rect 47298 21348 47362 21412
rect 47298 21268 47362 21332
rect 47298 21188 47362 21252
rect 47298 21108 47362 21172
rect 47298 21028 47362 21092
rect 47298 20948 47362 21012
rect 47298 20868 47362 20932
rect 47298 20788 47362 20852
rect 47298 20708 47362 20772
rect 47298 20628 47362 20692
rect 47298 20548 47362 20612
rect 47298 20468 47362 20532
rect 47298 20388 47362 20452
rect 47298 20308 47362 20372
rect 47298 20228 47362 20292
rect 47298 20148 47362 20212
rect 47298 20068 47362 20132
rect 47298 19988 47362 20052
rect 47298 19908 47362 19972
rect 47298 19828 47362 19892
rect 47298 19748 47362 19812
rect 47298 19668 47362 19732
rect 47298 19588 47362 19652
rect 47298 19508 47362 19572
rect 47298 19428 47362 19492
rect 47298 19348 47362 19412
rect 47298 19268 47362 19332
rect 47298 19188 47362 19252
rect 47298 19108 47362 19172
rect 47298 19028 47362 19092
rect 47298 18948 47362 19012
rect 47298 18868 47362 18932
rect 47298 18788 47362 18852
rect 47298 18708 47362 18772
rect 47298 18628 47362 18692
rect 47298 18548 47362 18612
rect 47298 18468 47362 18532
rect 47298 18388 47362 18452
rect 47298 18308 47362 18372
rect 47298 18228 47362 18292
rect 47298 18148 47362 18212
rect 47298 18068 47362 18132
rect 47298 17988 47362 18052
rect 47298 17908 47362 17972
rect 47298 17828 47362 17892
rect 47298 17748 47362 17812
rect 47298 17668 47362 17732
rect 47298 17588 47362 17652
rect 47298 17508 47362 17572
rect 47298 17428 47362 17492
rect 47298 17348 47362 17412
rect 47298 17268 47362 17332
rect 47298 17188 47362 17252
rect 47298 17108 47362 17172
rect 47298 17028 47362 17092
rect 47298 16948 47362 17012
rect 47298 16868 47362 16932
rect 47298 16788 47362 16852
rect 47298 16708 47362 16772
rect 47298 16628 47362 16692
rect 47298 16548 47362 16612
rect 47298 16468 47362 16532
rect 47298 16388 47362 16452
rect 47298 16308 47362 16372
rect 47298 16228 47362 16292
rect 47298 16148 47362 16212
rect 47298 16068 47362 16132
rect 47298 15988 47362 16052
rect 47298 15908 47362 15972
rect 47298 15828 47362 15892
rect -41168 15608 -41104 15672
rect -41168 15528 -41104 15592
rect -41168 15448 -41104 15512
rect -41168 15368 -41104 15432
rect -41168 15288 -41104 15352
rect -41168 15208 -41104 15272
rect -41168 15128 -41104 15192
rect -41168 15048 -41104 15112
rect -41168 14968 -41104 15032
rect -41168 14888 -41104 14952
rect -41168 14808 -41104 14872
rect -41168 14728 -41104 14792
rect -41168 14648 -41104 14712
rect -41168 14568 -41104 14632
rect -41168 14488 -41104 14552
rect -41168 14408 -41104 14472
rect -41168 14328 -41104 14392
rect -41168 14248 -41104 14312
rect -41168 14168 -41104 14232
rect -41168 14088 -41104 14152
rect -41168 14008 -41104 14072
rect -41168 13928 -41104 13992
rect -41168 13848 -41104 13912
rect -41168 13768 -41104 13832
rect -41168 13688 -41104 13752
rect -41168 13608 -41104 13672
rect -41168 13528 -41104 13592
rect -41168 13448 -41104 13512
rect -41168 13368 -41104 13432
rect -41168 13288 -41104 13352
rect -41168 13208 -41104 13272
rect -41168 13128 -41104 13192
rect -41168 13048 -41104 13112
rect -41168 12968 -41104 13032
rect -41168 12888 -41104 12952
rect -41168 12808 -41104 12872
rect -41168 12728 -41104 12792
rect -41168 12648 -41104 12712
rect -41168 12568 -41104 12632
rect -41168 12488 -41104 12552
rect -41168 12408 -41104 12472
rect -41168 12328 -41104 12392
rect -41168 12248 -41104 12312
rect -41168 12168 -41104 12232
rect -41168 12088 -41104 12152
rect -41168 12008 -41104 12072
rect -41168 11928 -41104 11992
rect -41168 11848 -41104 11912
rect -41168 11768 -41104 11832
rect -41168 11688 -41104 11752
rect -41168 11608 -41104 11672
rect -41168 11528 -41104 11592
rect -41168 11448 -41104 11512
rect -41168 11368 -41104 11432
rect -41168 11288 -41104 11352
rect -41168 11208 -41104 11272
rect -41168 11128 -41104 11192
rect -41168 11048 -41104 11112
rect -41168 10968 -41104 11032
rect -41168 10888 -41104 10952
rect -41168 10808 -41104 10872
rect -41168 10728 -41104 10792
rect -41168 10648 -41104 10712
rect -41168 10568 -41104 10632
rect -41168 10488 -41104 10552
rect -41168 10408 -41104 10472
rect -41168 10328 -41104 10392
rect -41168 10248 -41104 10312
rect -41168 10168 -41104 10232
rect -41168 10088 -41104 10152
rect -41168 10008 -41104 10072
rect -41168 9928 -41104 9992
rect -41168 9848 -41104 9912
rect -41168 9768 -41104 9832
rect -41168 9688 -41104 9752
rect -41168 9608 -41104 9672
rect -41168 9528 -41104 9592
rect -34849 15608 -34785 15672
rect -34849 15528 -34785 15592
rect -34849 15448 -34785 15512
rect -34849 15368 -34785 15432
rect -34849 15288 -34785 15352
rect -34849 15208 -34785 15272
rect -34849 15128 -34785 15192
rect -34849 15048 -34785 15112
rect -34849 14968 -34785 15032
rect -34849 14888 -34785 14952
rect -34849 14808 -34785 14872
rect -34849 14728 -34785 14792
rect -34849 14648 -34785 14712
rect -34849 14568 -34785 14632
rect -34849 14488 -34785 14552
rect -34849 14408 -34785 14472
rect -34849 14328 -34785 14392
rect -34849 14248 -34785 14312
rect -34849 14168 -34785 14232
rect -34849 14088 -34785 14152
rect -34849 14008 -34785 14072
rect -34849 13928 -34785 13992
rect -34849 13848 -34785 13912
rect -34849 13768 -34785 13832
rect -34849 13688 -34785 13752
rect -34849 13608 -34785 13672
rect -34849 13528 -34785 13592
rect -34849 13448 -34785 13512
rect -34849 13368 -34785 13432
rect -34849 13288 -34785 13352
rect -34849 13208 -34785 13272
rect -34849 13128 -34785 13192
rect -34849 13048 -34785 13112
rect -34849 12968 -34785 13032
rect -34849 12888 -34785 12952
rect -34849 12808 -34785 12872
rect -34849 12728 -34785 12792
rect -34849 12648 -34785 12712
rect -34849 12568 -34785 12632
rect -34849 12488 -34785 12552
rect -34849 12408 -34785 12472
rect -34849 12328 -34785 12392
rect -34849 12248 -34785 12312
rect -34849 12168 -34785 12232
rect -34849 12088 -34785 12152
rect -34849 12008 -34785 12072
rect -34849 11928 -34785 11992
rect -34849 11848 -34785 11912
rect -34849 11768 -34785 11832
rect -34849 11688 -34785 11752
rect -34849 11608 -34785 11672
rect -34849 11528 -34785 11592
rect -34849 11448 -34785 11512
rect -34849 11368 -34785 11432
rect -34849 11288 -34785 11352
rect -34849 11208 -34785 11272
rect -34849 11128 -34785 11192
rect -34849 11048 -34785 11112
rect -34849 10968 -34785 11032
rect -34849 10888 -34785 10952
rect -34849 10808 -34785 10872
rect -34849 10728 -34785 10792
rect -34849 10648 -34785 10712
rect -34849 10568 -34785 10632
rect -34849 10488 -34785 10552
rect -34849 10408 -34785 10472
rect -34849 10328 -34785 10392
rect -34849 10248 -34785 10312
rect -34849 10168 -34785 10232
rect -34849 10088 -34785 10152
rect -34849 10008 -34785 10072
rect -34849 9928 -34785 9992
rect -34849 9848 -34785 9912
rect -34849 9768 -34785 9832
rect -34849 9688 -34785 9752
rect -34849 9608 -34785 9672
rect -34849 9528 -34785 9592
rect -28530 15608 -28466 15672
rect -28530 15528 -28466 15592
rect -28530 15448 -28466 15512
rect -28530 15368 -28466 15432
rect -28530 15288 -28466 15352
rect -28530 15208 -28466 15272
rect -28530 15128 -28466 15192
rect -28530 15048 -28466 15112
rect -28530 14968 -28466 15032
rect -28530 14888 -28466 14952
rect -28530 14808 -28466 14872
rect -28530 14728 -28466 14792
rect -28530 14648 -28466 14712
rect -28530 14568 -28466 14632
rect -28530 14488 -28466 14552
rect -28530 14408 -28466 14472
rect -28530 14328 -28466 14392
rect -28530 14248 -28466 14312
rect -28530 14168 -28466 14232
rect -28530 14088 -28466 14152
rect -28530 14008 -28466 14072
rect -28530 13928 -28466 13992
rect -28530 13848 -28466 13912
rect -28530 13768 -28466 13832
rect -28530 13688 -28466 13752
rect -28530 13608 -28466 13672
rect -28530 13528 -28466 13592
rect -28530 13448 -28466 13512
rect -28530 13368 -28466 13432
rect -28530 13288 -28466 13352
rect -28530 13208 -28466 13272
rect -28530 13128 -28466 13192
rect -28530 13048 -28466 13112
rect -28530 12968 -28466 13032
rect -28530 12888 -28466 12952
rect -28530 12808 -28466 12872
rect -28530 12728 -28466 12792
rect -28530 12648 -28466 12712
rect -28530 12568 -28466 12632
rect -28530 12488 -28466 12552
rect -28530 12408 -28466 12472
rect -28530 12328 -28466 12392
rect -28530 12248 -28466 12312
rect -28530 12168 -28466 12232
rect -28530 12088 -28466 12152
rect -28530 12008 -28466 12072
rect -28530 11928 -28466 11992
rect -28530 11848 -28466 11912
rect -28530 11768 -28466 11832
rect -28530 11688 -28466 11752
rect -28530 11608 -28466 11672
rect -28530 11528 -28466 11592
rect -28530 11448 -28466 11512
rect -28530 11368 -28466 11432
rect -28530 11288 -28466 11352
rect -28530 11208 -28466 11272
rect -28530 11128 -28466 11192
rect -28530 11048 -28466 11112
rect -28530 10968 -28466 11032
rect -28530 10888 -28466 10952
rect -28530 10808 -28466 10872
rect -28530 10728 -28466 10792
rect -28530 10648 -28466 10712
rect -28530 10568 -28466 10632
rect -28530 10488 -28466 10552
rect -28530 10408 -28466 10472
rect -28530 10328 -28466 10392
rect -28530 10248 -28466 10312
rect -28530 10168 -28466 10232
rect -28530 10088 -28466 10152
rect -28530 10008 -28466 10072
rect -28530 9928 -28466 9992
rect -28530 9848 -28466 9912
rect -28530 9768 -28466 9832
rect -28530 9688 -28466 9752
rect -28530 9608 -28466 9672
rect -28530 9528 -28466 9592
rect -22211 15608 -22147 15672
rect -22211 15528 -22147 15592
rect -22211 15448 -22147 15512
rect -22211 15368 -22147 15432
rect -22211 15288 -22147 15352
rect -22211 15208 -22147 15272
rect -22211 15128 -22147 15192
rect -22211 15048 -22147 15112
rect -22211 14968 -22147 15032
rect -22211 14888 -22147 14952
rect -22211 14808 -22147 14872
rect -22211 14728 -22147 14792
rect -22211 14648 -22147 14712
rect -22211 14568 -22147 14632
rect -22211 14488 -22147 14552
rect -22211 14408 -22147 14472
rect -22211 14328 -22147 14392
rect -22211 14248 -22147 14312
rect -22211 14168 -22147 14232
rect -22211 14088 -22147 14152
rect -22211 14008 -22147 14072
rect -22211 13928 -22147 13992
rect -22211 13848 -22147 13912
rect -22211 13768 -22147 13832
rect -22211 13688 -22147 13752
rect -22211 13608 -22147 13672
rect -22211 13528 -22147 13592
rect -22211 13448 -22147 13512
rect -22211 13368 -22147 13432
rect -22211 13288 -22147 13352
rect -22211 13208 -22147 13272
rect -22211 13128 -22147 13192
rect -22211 13048 -22147 13112
rect -22211 12968 -22147 13032
rect -22211 12888 -22147 12952
rect -22211 12808 -22147 12872
rect -22211 12728 -22147 12792
rect -22211 12648 -22147 12712
rect -22211 12568 -22147 12632
rect -22211 12488 -22147 12552
rect -22211 12408 -22147 12472
rect -22211 12328 -22147 12392
rect -22211 12248 -22147 12312
rect -22211 12168 -22147 12232
rect -22211 12088 -22147 12152
rect -22211 12008 -22147 12072
rect -22211 11928 -22147 11992
rect -22211 11848 -22147 11912
rect -22211 11768 -22147 11832
rect -22211 11688 -22147 11752
rect -22211 11608 -22147 11672
rect -22211 11528 -22147 11592
rect -22211 11448 -22147 11512
rect -22211 11368 -22147 11432
rect -22211 11288 -22147 11352
rect -22211 11208 -22147 11272
rect -22211 11128 -22147 11192
rect -22211 11048 -22147 11112
rect -22211 10968 -22147 11032
rect -22211 10888 -22147 10952
rect -22211 10808 -22147 10872
rect -22211 10728 -22147 10792
rect -22211 10648 -22147 10712
rect -22211 10568 -22147 10632
rect -22211 10488 -22147 10552
rect -22211 10408 -22147 10472
rect -22211 10328 -22147 10392
rect -22211 10248 -22147 10312
rect -22211 10168 -22147 10232
rect -22211 10088 -22147 10152
rect -22211 10008 -22147 10072
rect -22211 9928 -22147 9992
rect -22211 9848 -22147 9912
rect -22211 9768 -22147 9832
rect -22211 9688 -22147 9752
rect -22211 9608 -22147 9672
rect -22211 9528 -22147 9592
rect -15892 15608 -15828 15672
rect -15892 15528 -15828 15592
rect -15892 15448 -15828 15512
rect -15892 15368 -15828 15432
rect -15892 15288 -15828 15352
rect -15892 15208 -15828 15272
rect -15892 15128 -15828 15192
rect -15892 15048 -15828 15112
rect -15892 14968 -15828 15032
rect -15892 14888 -15828 14952
rect -15892 14808 -15828 14872
rect -15892 14728 -15828 14792
rect -15892 14648 -15828 14712
rect -15892 14568 -15828 14632
rect -15892 14488 -15828 14552
rect -15892 14408 -15828 14472
rect -15892 14328 -15828 14392
rect -15892 14248 -15828 14312
rect -15892 14168 -15828 14232
rect -15892 14088 -15828 14152
rect -15892 14008 -15828 14072
rect -15892 13928 -15828 13992
rect -15892 13848 -15828 13912
rect -15892 13768 -15828 13832
rect -15892 13688 -15828 13752
rect -15892 13608 -15828 13672
rect -15892 13528 -15828 13592
rect -15892 13448 -15828 13512
rect -15892 13368 -15828 13432
rect -15892 13288 -15828 13352
rect -15892 13208 -15828 13272
rect -15892 13128 -15828 13192
rect -15892 13048 -15828 13112
rect -15892 12968 -15828 13032
rect -15892 12888 -15828 12952
rect -15892 12808 -15828 12872
rect -15892 12728 -15828 12792
rect -15892 12648 -15828 12712
rect -15892 12568 -15828 12632
rect -15892 12488 -15828 12552
rect -15892 12408 -15828 12472
rect -15892 12328 -15828 12392
rect -15892 12248 -15828 12312
rect -15892 12168 -15828 12232
rect -15892 12088 -15828 12152
rect -15892 12008 -15828 12072
rect -15892 11928 -15828 11992
rect -15892 11848 -15828 11912
rect -15892 11768 -15828 11832
rect -15892 11688 -15828 11752
rect -15892 11608 -15828 11672
rect -15892 11528 -15828 11592
rect -15892 11448 -15828 11512
rect -15892 11368 -15828 11432
rect -15892 11288 -15828 11352
rect -15892 11208 -15828 11272
rect -15892 11128 -15828 11192
rect -15892 11048 -15828 11112
rect -15892 10968 -15828 11032
rect -15892 10888 -15828 10952
rect -15892 10808 -15828 10872
rect -15892 10728 -15828 10792
rect -15892 10648 -15828 10712
rect -15892 10568 -15828 10632
rect -15892 10488 -15828 10552
rect -15892 10408 -15828 10472
rect -15892 10328 -15828 10392
rect -15892 10248 -15828 10312
rect -15892 10168 -15828 10232
rect -15892 10088 -15828 10152
rect -15892 10008 -15828 10072
rect -15892 9928 -15828 9992
rect -15892 9848 -15828 9912
rect -15892 9768 -15828 9832
rect -15892 9688 -15828 9752
rect -15892 9608 -15828 9672
rect -15892 9528 -15828 9592
rect -9573 15608 -9509 15672
rect -9573 15528 -9509 15592
rect -9573 15448 -9509 15512
rect -9573 15368 -9509 15432
rect -9573 15288 -9509 15352
rect -9573 15208 -9509 15272
rect -9573 15128 -9509 15192
rect -9573 15048 -9509 15112
rect -9573 14968 -9509 15032
rect -9573 14888 -9509 14952
rect -9573 14808 -9509 14872
rect -9573 14728 -9509 14792
rect -9573 14648 -9509 14712
rect -9573 14568 -9509 14632
rect -9573 14488 -9509 14552
rect -9573 14408 -9509 14472
rect -9573 14328 -9509 14392
rect -9573 14248 -9509 14312
rect -9573 14168 -9509 14232
rect -9573 14088 -9509 14152
rect -9573 14008 -9509 14072
rect -9573 13928 -9509 13992
rect -9573 13848 -9509 13912
rect -9573 13768 -9509 13832
rect -9573 13688 -9509 13752
rect -9573 13608 -9509 13672
rect -9573 13528 -9509 13592
rect -9573 13448 -9509 13512
rect -9573 13368 -9509 13432
rect -9573 13288 -9509 13352
rect -9573 13208 -9509 13272
rect -9573 13128 -9509 13192
rect -9573 13048 -9509 13112
rect -9573 12968 -9509 13032
rect -9573 12888 -9509 12952
rect -9573 12808 -9509 12872
rect -9573 12728 -9509 12792
rect -9573 12648 -9509 12712
rect -9573 12568 -9509 12632
rect -9573 12488 -9509 12552
rect -9573 12408 -9509 12472
rect -9573 12328 -9509 12392
rect -9573 12248 -9509 12312
rect -9573 12168 -9509 12232
rect -9573 12088 -9509 12152
rect -9573 12008 -9509 12072
rect -9573 11928 -9509 11992
rect -9573 11848 -9509 11912
rect -9573 11768 -9509 11832
rect -9573 11688 -9509 11752
rect -9573 11608 -9509 11672
rect -9573 11528 -9509 11592
rect -9573 11448 -9509 11512
rect -9573 11368 -9509 11432
rect -9573 11288 -9509 11352
rect -9573 11208 -9509 11272
rect -9573 11128 -9509 11192
rect -9573 11048 -9509 11112
rect -9573 10968 -9509 11032
rect -9573 10888 -9509 10952
rect -9573 10808 -9509 10872
rect -9573 10728 -9509 10792
rect -9573 10648 -9509 10712
rect -9573 10568 -9509 10632
rect -9573 10488 -9509 10552
rect -9573 10408 -9509 10472
rect -9573 10328 -9509 10392
rect -9573 10248 -9509 10312
rect -9573 10168 -9509 10232
rect -9573 10088 -9509 10152
rect -9573 10008 -9509 10072
rect -9573 9928 -9509 9992
rect -9573 9848 -9509 9912
rect -9573 9768 -9509 9832
rect -9573 9688 -9509 9752
rect -9573 9608 -9509 9672
rect -9573 9528 -9509 9592
rect -3254 15608 -3190 15672
rect -3254 15528 -3190 15592
rect -3254 15448 -3190 15512
rect -3254 15368 -3190 15432
rect -3254 15288 -3190 15352
rect -3254 15208 -3190 15272
rect -3254 15128 -3190 15192
rect -3254 15048 -3190 15112
rect -3254 14968 -3190 15032
rect -3254 14888 -3190 14952
rect -3254 14808 -3190 14872
rect -3254 14728 -3190 14792
rect -3254 14648 -3190 14712
rect -3254 14568 -3190 14632
rect -3254 14488 -3190 14552
rect -3254 14408 -3190 14472
rect -3254 14328 -3190 14392
rect -3254 14248 -3190 14312
rect -3254 14168 -3190 14232
rect -3254 14088 -3190 14152
rect -3254 14008 -3190 14072
rect -3254 13928 -3190 13992
rect -3254 13848 -3190 13912
rect -3254 13768 -3190 13832
rect -3254 13688 -3190 13752
rect -3254 13608 -3190 13672
rect -3254 13528 -3190 13592
rect -3254 13448 -3190 13512
rect -3254 13368 -3190 13432
rect -3254 13288 -3190 13352
rect -3254 13208 -3190 13272
rect -3254 13128 -3190 13192
rect -3254 13048 -3190 13112
rect -3254 12968 -3190 13032
rect -3254 12888 -3190 12952
rect -3254 12808 -3190 12872
rect -3254 12728 -3190 12792
rect -3254 12648 -3190 12712
rect -3254 12568 -3190 12632
rect -3254 12488 -3190 12552
rect -3254 12408 -3190 12472
rect -3254 12328 -3190 12392
rect -3254 12248 -3190 12312
rect -3254 12168 -3190 12232
rect -3254 12088 -3190 12152
rect -3254 12008 -3190 12072
rect -3254 11928 -3190 11992
rect -3254 11848 -3190 11912
rect -3254 11768 -3190 11832
rect -3254 11688 -3190 11752
rect -3254 11608 -3190 11672
rect -3254 11528 -3190 11592
rect -3254 11448 -3190 11512
rect -3254 11368 -3190 11432
rect -3254 11288 -3190 11352
rect -3254 11208 -3190 11272
rect -3254 11128 -3190 11192
rect -3254 11048 -3190 11112
rect -3254 10968 -3190 11032
rect -3254 10888 -3190 10952
rect -3254 10808 -3190 10872
rect -3254 10728 -3190 10792
rect -3254 10648 -3190 10712
rect -3254 10568 -3190 10632
rect -3254 10488 -3190 10552
rect -3254 10408 -3190 10472
rect -3254 10328 -3190 10392
rect -3254 10248 -3190 10312
rect -3254 10168 -3190 10232
rect -3254 10088 -3190 10152
rect -3254 10008 -3190 10072
rect -3254 9928 -3190 9992
rect -3254 9848 -3190 9912
rect -3254 9768 -3190 9832
rect -3254 9688 -3190 9752
rect -3254 9608 -3190 9672
rect -3254 9528 -3190 9592
rect 3065 15608 3129 15672
rect 3065 15528 3129 15592
rect 3065 15448 3129 15512
rect 3065 15368 3129 15432
rect 3065 15288 3129 15352
rect 3065 15208 3129 15272
rect 3065 15128 3129 15192
rect 3065 15048 3129 15112
rect 3065 14968 3129 15032
rect 3065 14888 3129 14952
rect 3065 14808 3129 14872
rect 3065 14728 3129 14792
rect 3065 14648 3129 14712
rect 3065 14568 3129 14632
rect 3065 14488 3129 14552
rect 3065 14408 3129 14472
rect 3065 14328 3129 14392
rect 3065 14248 3129 14312
rect 3065 14168 3129 14232
rect 3065 14088 3129 14152
rect 3065 14008 3129 14072
rect 3065 13928 3129 13992
rect 3065 13848 3129 13912
rect 3065 13768 3129 13832
rect 3065 13688 3129 13752
rect 3065 13608 3129 13672
rect 3065 13528 3129 13592
rect 3065 13448 3129 13512
rect 3065 13368 3129 13432
rect 3065 13288 3129 13352
rect 3065 13208 3129 13272
rect 3065 13128 3129 13192
rect 3065 13048 3129 13112
rect 3065 12968 3129 13032
rect 3065 12888 3129 12952
rect 3065 12808 3129 12872
rect 3065 12728 3129 12792
rect 3065 12648 3129 12712
rect 3065 12568 3129 12632
rect 3065 12488 3129 12552
rect 3065 12408 3129 12472
rect 3065 12328 3129 12392
rect 3065 12248 3129 12312
rect 3065 12168 3129 12232
rect 3065 12088 3129 12152
rect 3065 12008 3129 12072
rect 3065 11928 3129 11992
rect 3065 11848 3129 11912
rect 3065 11768 3129 11832
rect 3065 11688 3129 11752
rect 3065 11608 3129 11672
rect 3065 11528 3129 11592
rect 3065 11448 3129 11512
rect 3065 11368 3129 11432
rect 3065 11288 3129 11352
rect 3065 11208 3129 11272
rect 3065 11128 3129 11192
rect 3065 11048 3129 11112
rect 3065 10968 3129 11032
rect 3065 10888 3129 10952
rect 3065 10808 3129 10872
rect 3065 10728 3129 10792
rect 3065 10648 3129 10712
rect 3065 10568 3129 10632
rect 3065 10488 3129 10552
rect 3065 10408 3129 10472
rect 3065 10328 3129 10392
rect 3065 10248 3129 10312
rect 3065 10168 3129 10232
rect 3065 10088 3129 10152
rect 3065 10008 3129 10072
rect 3065 9928 3129 9992
rect 3065 9848 3129 9912
rect 3065 9768 3129 9832
rect 3065 9688 3129 9752
rect 3065 9608 3129 9672
rect 3065 9528 3129 9592
rect 9384 15608 9448 15672
rect 9384 15528 9448 15592
rect 9384 15448 9448 15512
rect 9384 15368 9448 15432
rect 9384 15288 9448 15352
rect 9384 15208 9448 15272
rect 9384 15128 9448 15192
rect 9384 15048 9448 15112
rect 9384 14968 9448 15032
rect 9384 14888 9448 14952
rect 9384 14808 9448 14872
rect 9384 14728 9448 14792
rect 9384 14648 9448 14712
rect 9384 14568 9448 14632
rect 9384 14488 9448 14552
rect 9384 14408 9448 14472
rect 9384 14328 9448 14392
rect 9384 14248 9448 14312
rect 9384 14168 9448 14232
rect 9384 14088 9448 14152
rect 9384 14008 9448 14072
rect 9384 13928 9448 13992
rect 9384 13848 9448 13912
rect 9384 13768 9448 13832
rect 9384 13688 9448 13752
rect 9384 13608 9448 13672
rect 9384 13528 9448 13592
rect 9384 13448 9448 13512
rect 9384 13368 9448 13432
rect 9384 13288 9448 13352
rect 9384 13208 9448 13272
rect 9384 13128 9448 13192
rect 9384 13048 9448 13112
rect 9384 12968 9448 13032
rect 9384 12888 9448 12952
rect 9384 12808 9448 12872
rect 9384 12728 9448 12792
rect 9384 12648 9448 12712
rect 9384 12568 9448 12632
rect 9384 12488 9448 12552
rect 9384 12408 9448 12472
rect 9384 12328 9448 12392
rect 9384 12248 9448 12312
rect 9384 12168 9448 12232
rect 9384 12088 9448 12152
rect 9384 12008 9448 12072
rect 9384 11928 9448 11992
rect 9384 11848 9448 11912
rect 9384 11768 9448 11832
rect 9384 11688 9448 11752
rect 9384 11608 9448 11672
rect 9384 11528 9448 11592
rect 9384 11448 9448 11512
rect 9384 11368 9448 11432
rect 9384 11288 9448 11352
rect 9384 11208 9448 11272
rect 9384 11128 9448 11192
rect 9384 11048 9448 11112
rect 9384 10968 9448 11032
rect 9384 10888 9448 10952
rect 9384 10808 9448 10872
rect 9384 10728 9448 10792
rect 9384 10648 9448 10712
rect 9384 10568 9448 10632
rect 9384 10488 9448 10552
rect 9384 10408 9448 10472
rect 9384 10328 9448 10392
rect 9384 10248 9448 10312
rect 9384 10168 9448 10232
rect 9384 10088 9448 10152
rect 9384 10008 9448 10072
rect 9384 9928 9448 9992
rect 9384 9848 9448 9912
rect 9384 9768 9448 9832
rect 9384 9688 9448 9752
rect 9384 9608 9448 9672
rect 9384 9528 9448 9592
rect 15703 15608 15767 15672
rect 15703 15528 15767 15592
rect 15703 15448 15767 15512
rect 15703 15368 15767 15432
rect 15703 15288 15767 15352
rect 15703 15208 15767 15272
rect 15703 15128 15767 15192
rect 15703 15048 15767 15112
rect 15703 14968 15767 15032
rect 15703 14888 15767 14952
rect 15703 14808 15767 14872
rect 15703 14728 15767 14792
rect 15703 14648 15767 14712
rect 15703 14568 15767 14632
rect 15703 14488 15767 14552
rect 15703 14408 15767 14472
rect 15703 14328 15767 14392
rect 15703 14248 15767 14312
rect 15703 14168 15767 14232
rect 15703 14088 15767 14152
rect 15703 14008 15767 14072
rect 15703 13928 15767 13992
rect 15703 13848 15767 13912
rect 15703 13768 15767 13832
rect 15703 13688 15767 13752
rect 15703 13608 15767 13672
rect 15703 13528 15767 13592
rect 15703 13448 15767 13512
rect 15703 13368 15767 13432
rect 15703 13288 15767 13352
rect 15703 13208 15767 13272
rect 15703 13128 15767 13192
rect 15703 13048 15767 13112
rect 15703 12968 15767 13032
rect 15703 12888 15767 12952
rect 15703 12808 15767 12872
rect 15703 12728 15767 12792
rect 15703 12648 15767 12712
rect 15703 12568 15767 12632
rect 15703 12488 15767 12552
rect 15703 12408 15767 12472
rect 15703 12328 15767 12392
rect 15703 12248 15767 12312
rect 15703 12168 15767 12232
rect 15703 12088 15767 12152
rect 15703 12008 15767 12072
rect 15703 11928 15767 11992
rect 15703 11848 15767 11912
rect 15703 11768 15767 11832
rect 15703 11688 15767 11752
rect 15703 11608 15767 11672
rect 15703 11528 15767 11592
rect 15703 11448 15767 11512
rect 15703 11368 15767 11432
rect 15703 11288 15767 11352
rect 15703 11208 15767 11272
rect 15703 11128 15767 11192
rect 15703 11048 15767 11112
rect 15703 10968 15767 11032
rect 15703 10888 15767 10952
rect 15703 10808 15767 10872
rect 15703 10728 15767 10792
rect 15703 10648 15767 10712
rect 15703 10568 15767 10632
rect 15703 10488 15767 10552
rect 15703 10408 15767 10472
rect 15703 10328 15767 10392
rect 15703 10248 15767 10312
rect 15703 10168 15767 10232
rect 15703 10088 15767 10152
rect 15703 10008 15767 10072
rect 15703 9928 15767 9992
rect 15703 9848 15767 9912
rect 15703 9768 15767 9832
rect 15703 9688 15767 9752
rect 15703 9608 15767 9672
rect 15703 9528 15767 9592
rect 22022 15608 22086 15672
rect 22022 15528 22086 15592
rect 22022 15448 22086 15512
rect 22022 15368 22086 15432
rect 22022 15288 22086 15352
rect 22022 15208 22086 15272
rect 22022 15128 22086 15192
rect 22022 15048 22086 15112
rect 22022 14968 22086 15032
rect 22022 14888 22086 14952
rect 22022 14808 22086 14872
rect 22022 14728 22086 14792
rect 22022 14648 22086 14712
rect 22022 14568 22086 14632
rect 22022 14488 22086 14552
rect 22022 14408 22086 14472
rect 22022 14328 22086 14392
rect 22022 14248 22086 14312
rect 22022 14168 22086 14232
rect 22022 14088 22086 14152
rect 22022 14008 22086 14072
rect 22022 13928 22086 13992
rect 22022 13848 22086 13912
rect 22022 13768 22086 13832
rect 22022 13688 22086 13752
rect 22022 13608 22086 13672
rect 22022 13528 22086 13592
rect 22022 13448 22086 13512
rect 22022 13368 22086 13432
rect 22022 13288 22086 13352
rect 22022 13208 22086 13272
rect 22022 13128 22086 13192
rect 22022 13048 22086 13112
rect 22022 12968 22086 13032
rect 22022 12888 22086 12952
rect 22022 12808 22086 12872
rect 22022 12728 22086 12792
rect 22022 12648 22086 12712
rect 22022 12568 22086 12632
rect 22022 12488 22086 12552
rect 22022 12408 22086 12472
rect 22022 12328 22086 12392
rect 22022 12248 22086 12312
rect 22022 12168 22086 12232
rect 22022 12088 22086 12152
rect 22022 12008 22086 12072
rect 22022 11928 22086 11992
rect 22022 11848 22086 11912
rect 22022 11768 22086 11832
rect 22022 11688 22086 11752
rect 22022 11608 22086 11672
rect 22022 11528 22086 11592
rect 22022 11448 22086 11512
rect 22022 11368 22086 11432
rect 22022 11288 22086 11352
rect 22022 11208 22086 11272
rect 22022 11128 22086 11192
rect 22022 11048 22086 11112
rect 22022 10968 22086 11032
rect 22022 10888 22086 10952
rect 22022 10808 22086 10872
rect 22022 10728 22086 10792
rect 22022 10648 22086 10712
rect 22022 10568 22086 10632
rect 22022 10488 22086 10552
rect 22022 10408 22086 10472
rect 22022 10328 22086 10392
rect 22022 10248 22086 10312
rect 22022 10168 22086 10232
rect 22022 10088 22086 10152
rect 22022 10008 22086 10072
rect 22022 9928 22086 9992
rect 22022 9848 22086 9912
rect 22022 9768 22086 9832
rect 22022 9688 22086 9752
rect 22022 9608 22086 9672
rect 22022 9528 22086 9592
rect 28341 15608 28405 15672
rect 28341 15528 28405 15592
rect 28341 15448 28405 15512
rect 28341 15368 28405 15432
rect 28341 15288 28405 15352
rect 28341 15208 28405 15272
rect 28341 15128 28405 15192
rect 28341 15048 28405 15112
rect 28341 14968 28405 15032
rect 28341 14888 28405 14952
rect 28341 14808 28405 14872
rect 28341 14728 28405 14792
rect 28341 14648 28405 14712
rect 28341 14568 28405 14632
rect 28341 14488 28405 14552
rect 28341 14408 28405 14472
rect 28341 14328 28405 14392
rect 28341 14248 28405 14312
rect 28341 14168 28405 14232
rect 28341 14088 28405 14152
rect 28341 14008 28405 14072
rect 28341 13928 28405 13992
rect 28341 13848 28405 13912
rect 28341 13768 28405 13832
rect 28341 13688 28405 13752
rect 28341 13608 28405 13672
rect 28341 13528 28405 13592
rect 28341 13448 28405 13512
rect 28341 13368 28405 13432
rect 28341 13288 28405 13352
rect 28341 13208 28405 13272
rect 28341 13128 28405 13192
rect 28341 13048 28405 13112
rect 28341 12968 28405 13032
rect 28341 12888 28405 12952
rect 28341 12808 28405 12872
rect 28341 12728 28405 12792
rect 28341 12648 28405 12712
rect 28341 12568 28405 12632
rect 28341 12488 28405 12552
rect 28341 12408 28405 12472
rect 28341 12328 28405 12392
rect 28341 12248 28405 12312
rect 28341 12168 28405 12232
rect 28341 12088 28405 12152
rect 28341 12008 28405 12072
rect 28341 11928 28405 11992
rect 28341 11848 28405 11912
rect 28341 11768 28405 11832
rect 28341 11688 28405 11752
rect 28341 11608 28405 11672
rect 28341 11528 28405 11592
rect 28341 11448 28405 11512
rect 28341 11368 28405 11432
rect 28341 11288 28405 11352
rect 28341 11208 28405 11272
rect 28341 11128 28405 11192
rect 28341 11048 28405 11112
rect 28341 10968 28405 11032
rect 28341 10888 28405 10952
rect 28341 10808 28405 10872
rect 28341 10728 28405 10792
rect 28341 10648 28405 10712
rect 28341 10568 28405 10632
rect 28341 10488 28405 10552
rect 28341 10408 28405 10472
rect 28341 10328 28405 10392
rect 28341 10248 28405 10312
rect 28341 10168 28405 10232
rect 28341 10088 28405 10152
rect 28341 10008 28405 10072
rect 28341 9928 28405 9992
rect 28341 9848 28405 9912
rect 28341 9768 28405 9832
rect 28341 9688 28405 9752
rect 28341 9608 28405 9672
rect 28341 9528 28405 9592
rect 34660 15608 34724 15672
rect 34660 15528 34724 15592
rect 34660 15448 34724 15512
rect 34660 15368 34724 15432
rect 34660 15288 34724 15352
rect 34660 15208 34724 15272
rect 34660 15128 34724 15192
rect 34660 15048 34724 15112
rect 34660 14968 34724 15032
rect 34660 14888 34724 14952
rect 34660 14808 34724 14872
rect 34660 14728 34724 14792
rect 34660 14648 34724 14712
rect 34660 14568 34724 14632
rect 34660 14488 34724 14552
rect 34660 14408 34724 14472
rect 34660 14328 34724 14392
rect 34660 14248 34724 14312
rect 34660 14168 34724 14232
rect 34660 14088 34724 14152
rect 34660 14008 34724 14072
rect 34660 13928 34724 13992
rect 34660 13848 34724 13912
rect 34660 13768 34724 13832
rect 34660 13688 34724 13752
rect 34660 13608 34724 13672
rect 34660 13528 34724 13592
rect 34660 13448 34724 13512
rect 34660 13368 34724 13432
rect 34660 13288 34724 13352
rect 34660 13208 34724 13272
rect 34660 13128 34724 13192
rect 34660 13048 34724 13112
rect 34660 12968 34724 13032
rect 34660 12888 34724 12952
rect 34660 12808 34724 12872
rect 34660 12728 34724 12792
rect 34660 12648 34724 12712
rect 34660 12568 34724 12632
rect 34660 12488 34724 12552
rect 34660 12408 34724 12472
rect 34660 12328 34724 12392
rect 34660 12248 34724 12312
rect 34660 12168 34724 12232
rect 34660 12088 34724 12152
rect 34660 12008 34724 12072
rect 34660 11928 34724 11992
rect 34660 11848 34724 11912
rect 34660 11768 34724 11832
rect 34660 11688 34724 11752
rect 34660 11608 34724 11672
rect 34660 11528 34724 11592
rect 34660 11448 34724 11512
rect 34660 11368 34724 11432
rect 34660 11288 34724 11352
rect 34660 11208 34724 11272
rect 34660 11128 34724 11192
rect 34660 11048 34724 11112
rect 34660 10968 34724 11032
rect 34660 10888 34724 10952
rect 34660 10808 34724 10872
rect 34660 10728 34724 10792
rect 34660 10648 34724 10712
rect 34660 10568 34724 10632
rect 34660 10488 34724 10552
rect 34660 10408 34724 10472
rect 34660 10328 34724 10392
rect 34660 10248 34724 10312
rect 34660 10168 34724 10232
rect 34660 10088 34724 10152
rect 34660 10008 34724 10072
rect 34660 9928 34724 9992
rect 34660 9848 34724 9912
rect 34660 9768 34724 9832
rect 34660 9688 34724 9752
rect 34660 9608 34724 9672
rect 34660 9528 34724 9592
rect 40979 15608 41043 15672
rect 40979 15528 41043 15592
rect 40979 15448 41043 15512
rect 40979 15368 41043 15432
rect 40979 15288 41043 15352
rect 40979 15208 41043 15272
rect 40979 15128 41043 15192
rect 40979 15048 41043 15112
rect 40979 14968 41043 15032
rect 40979 14888 41043 14952
rect 40979 14808 41043 14872
rect 40979 14728 41043 14792
rect 40979 14648 41043 14712
rect 40979 14568 41043 14632
rect 40979 14488 41043 14552
rect 40979 14408 41043 14472
rect 40979 14328 41043 14392
rect 40979 14248 41043 14312
rect 40979 14168 41043 14232
rect 40979 14088 41043 14152
rect 40979 14008 41043 14072
rect 40979 13928 41043 13992
rect 40979 13848 41043 13912
rect 40979 13768 41043 13832
rect 40979 13688 41043 13752
rect 40979 13608 41043 13672
rect 40979 13528 41043 13592
rect 40979 13448 41043 13512
rect 40979 13368 41043 13432
rect 40979 13288 41043 13352
rect 40979 13208 41043 13272
rect 40979 13128 41043 13192
rect 40979 13048 41043 13112
rect 40979 12968 41043 13032
rect 40979 12888 41043 12952
rect 40979 12808 41043 12872
rect 40979 12728 41043 12792
rect 40979 12648 41043 12712
rect 40979 12568 41043 12632
rect 40979 12488 41043 12552
rect 40979 12408 41043 12472
rect 40979 12328 41043 12392
rect 40979 12248 41043 12312
rect 40979 12168 41043 12232
rect 40979 12088 41043 12152
rect 40979 12008 41043 12072
rect 40979 11928 41043 11992
rect 40979 11848 41043 11912
rect 40979 11768 41043 11832
rect 40979 11688 41043 11752
rect 40979 11608 41043 11672
rect 40979 11528 41043 11592
rect 40979 11448 41043 11512
rect 40979 11368 41043 11432
rect 40979 11288 41043 11352
rect 40979 11208 41043 11272
rect 40979 11128 41043 11192
rect 40979 11048 41043 11112
rect 40979 10968 41043 11032
rect 40979 10888 41043 10952
rect 40979 10808 41043 10872
rect 40979 10728 41043 10792
rect 40979 10648 41043 10712
rect 40979 10568 41043 10632
rect 40979 10488 41043 10552
rect 40979 10408 41043 10472
rect 40979 10328 41043 10392
rect 40979 10248 41043 10312
rect 40979 10168 41043 10232
rect 40979 10088 41043 10152
rect 40979 10008 41043 10072
rect 40979 9928 41043 9992
rect 40979 9848 41043 9912
rect 40979 9768 41043 9832
rect 40979 9688 41043 9752
rect 40979 9608 41043 9672
rect 40979 9528 41043 9592
rect 47298 15608 47362 15672
rect 47298 15528 47362 15592
rect 47298 15448 47362 15512
rect 47298 15368 47362 15432
rect 47298 15288 47362 15352
rect 47298 15208 47362 15272
rect 47298 15128 47362 15192
rect 47298 15048 47362 15112
rect 47298 14968 47362 15032
rect 47298 14888 47362 14952
rect 47298 14808 47362 14872
rect 47298 14728 47362 14792
rect 47298 14648 47362 14712
rect 47298 14568 47362 14632
rect 47298 14488 47362 14552
rect 47298 14408 47362 14472
rect 47298 14328 47362 14392
rect 47298 14248 47362 14312
rect 47298 14168 47362 14232
rect 47298 14088 47362 14152
rect 47298 14008 47362 14072
rect 47298 13928 47362 13992
rect 47298 13848 47362 13912
rect 47298 13768 47362 13832
rect 47298 13688 47362 13752
rect 47298 13608 47362 13672
rect 47298 13528 47362 13592
rect 47298 13448 47362 13512
rect 47298 13368 47362 13432
rect 47298 13288 47362 13352
rect 47298 13208 47362 13272
rect 47298 13128 47362 13192
rect 47298 13048 47362 13112
rect 47298 12968 47362 13032
rect 47298 12888 47362 12952
rect 47298 12808 47362 12872
rect 47298 12728 47362 12792
rect 47298 12648 47362 12712
rect 47298 12568 47362 12632
rect 47298 12488 47362 12552
rect 47298 12408 47362 12472
rect 47298 12328 47362 12392
rect 47298 12248 47362 12312
rect 47298 12168 47362 12232
rect 47298 12088 47362 12152
rect 47298 12008 47362 12072
rect 47298 11928 47362 11992
rect 47298 11848 47362 11912
rect 47298 11768 47362 11832
rect 47298 11688 47362 11752
rect 47298 11608 47362 11672
rect 47298 11528 47362 11592
rect 47298 11448 47362 11512
rect 47298 11368 47362 11432
rect 47298 11288 47362 11352
rect 47298 11208 47362 11272
rect 47298 11128 47362 11192
rect 47298 11048 47362 11112
rect 47298 10968 47362 11032
rect 47298 10888 47362 10952
rect 47298 10808 47362 10872
rect 47298 10728 47362 10792
rect 47298 10648 47362 10712
rect 47298 10568 47362 10632
rect 47298 10488 47362 10552
rect 47298 10408 47362 10472
rect 47298 10328 47362 10392
rect 47298 10248 47362 10312
rect 47298 10168 47362 10232
rect 47298 10088 47362 10152
rect 47298 10008 47362 10072
rect 47298 9928 47362 9992
rect 47298 9848 47362 9912
rect 47298 9768 47362 9832
rect 47298 9688 47362 9752
rect 47298 9608 47362 9672
rect 47298 9528 47362 9592
rect -41168 9308 -41104 9372
rect -41168 9228 -41104 9292
rect -41168 9148 -41104 9212
rect -41168 9068 -41104 9132
rect -41168 8988 -41104 9052
rect -41168 8908 -41104 8972
rect -41168 8828 -41104 8892
rect -41168 8748 -41104 8812
rect -41168 8668 -41104 8732
rect -41168 8588 -41104 8652
rect -41168 8508 -41104 8572
rect -41168 8428 -41104 8492
rect -41168 8348 -41104 8412
rect -41168 8268 -41104 8332
rect -41168 8188 -41104 8252
rect -41168 8108 -41104 8172
rect -41168 8028 -41104 8092
rect -41168 7948 -41104 8012
rect -41168 7868 -41104 7932
rect -41168 7788 -41104 7852
rect -41168 7708 -41104 7772
rect -41168 7628 -41104 7692
rect -41168 7548 -41104 7612
rect -41168 7468 -41104 7532
rect -41168 7388 -41104 7452
rect -41168 7308 -41104 7372
rect -41168 7228 -41104 7292
rect -41168 7148 -41104 7212
rect -41168 7068 -41104 7132
rect -41168 6988 -41104 7052
rect -41168 6908 -41104 6972
rect -41168 6828 -41104 6892
rect -41168 6748 -41104 6812
rect -41168 6668 -41104 6732
rect -41168 6588 -41104 6652
rect -41168 6508 -41104 6572
rect -41168 6428 -41104 6492
rect -41168 6348 -41104 6412
rect -41168 6268 -41104 6332
rect -41168 6188 -41104 6252
rect -41168 6108 -41104 6172
rect -41168 6028 -41104 6092
rect -41168 5948 -41104 6012
rect -41168 5868 -41104 5932
rect -41168 5788 -41104 5852
rect -41168 5708 -41104 5772
rect -41168 5628 -41104 5692
rect -41168 5548 -41104 5612
rect -41168 5468 -41104 5532
rect -41168 5388 -41104 5452
rect -41168 5308 -41104 5372
rect -41168 5228 -41104 5292
rect -41168 5148 -41104 5212
rect -41168 5068 -41104 5132
rect -41168 4988 -41104 5052
rect -41168 4908 -41104 4972
rect -41168 4828 -41104 4892
rect -41168 4748 -41104 4812
rect -41168 4668 -41104 4732
rect -41168 4588 -41104 4652
rect -41168 4508 -41104 4572
rect -41168 4428 -41104 4492
rect -41168 4348 -41104 4412
rect -41168 4268 -41104 4332
rect -41168 4188 -41104 4252
rect -41168 4108 -41104 4172
rect -41168 4028 -41104 4092
rect -41168 3948 -41104 4012
rect -41168 3868 -41104 3932
rect -41168 3788 -41104 3852
rect -41168 3708 -41104 3772
rect -41168 3628 -41104 3692
rect -41168 3548 -41104 3612
rect -41168 3468 -41104 3532
rect -41168 3388 -41104 3452
rect -41168 3308 -41104 3372
rect -41168 3228 -41104 3292
rect -34849 9308 -34785 9372
rect -34849 9228 -34785 9292
rect -34849 9148 -34785 9212
rect -34849 9068 -34785 9132
rect -34849 8988 -34785 9052
rect -34849 8908 -34785 8972
rect -34849 8828 -34785 8892
rect -34849 8748 -34785 8812
rect -34849 8668 -34785 8732
rect -34849 8588 -34785 8652
rect -34849 8508 -34785 8572
rect -34849 8428 -34785 8492
rect -34849 8348 -34785 8412
rect -34849 8268 -34785 8332
rect -34849 8188 -34785 8252
rect -34849 8108 -34785 8172
rect -34849 8028 -34785 8092
rect -34849 7948 -34785 8012
rect -34849 7868 -34785 7932
rect -34849 7788 -34785 7852
rect -34849 7708 -34785 7772
rect -34849 7628 -34785 7692
rect -34849 7548 -34785 7612
rect -34849 7468 -34785 7532
rect -34849 7388 -34785 7452
rect -34849 7308 -34785 7372
rect -34849 7228 -34785 7292
rect -34849 7148 -34785 7212
rect -34849 7068 -34785 7132
rect -34849 6988 -34785 7052
rect -34849 6908 -34785 6972
rect -34849 6828 -34785 6892
rect -34849 6748 -34785 6812
rect -34849 6668 -34785 6732
rect -34849 6588 -34785 6652
rect -34849 6508 -34785 6572
rect -34849 6428 -34785 6492
rect -34849 6348 -34785 6412
rect -34849 6268 -34785 6332
rect -34849 6188 -34785 6252
rect -34849 6108 -34785 6172
rect -34849 6028 -34785 6092
rect -34849 5948 -34785 6012
rect -34849 5868 -34785 5932
rect -34849 5788 -34785 5852
rect -34849 5708 -34785 5772
rect -34849 5628 -34785 5692
rect -34849 5548 -34785 5612
rect -34849 5468 -34785 5532
rect -34849 5388 -34785 5452
rect -34849 5308 -34785 5372
rect -34849 5228 -34785 5292
rect -34849 5148 -34785 5212
rect -34849 5068 -34785 5132
rect -34849 4988 -34785 5052
rect -34849 4908 -34785 4972
rect -34849 4828 -34785 4892
rect -34849 4748 -34785 4812
rect -34849 4668 -34785 4732
rect -34849 4588 -34785 4652
rect -34849 4508 -34785 4572
rect -34849 4428 -34785 4492
rect -34849 4348 -34785 4412
rect -34849 4268 -34785 4332
rect -34849 4188 -34785 4252
rect -34849 4108 -34785 4172
rect -34849 4028 -34785 4092
rect -34849 3948 -34785 4012
rect -34849 3868 -34785 3932
rect -34849 3788 -34785 3852
rect -34849 3708 -34785 3772
rect -34849 3628 -34785 3692
rect -34849 3548 -34785 3612
rect -34849 3468 -34785 3532
rect -34849 3388 -34785 3452
rect -34849 3308 -34785 3372
rect -34849 3228 -34785 3292
rect -28530 9308 -28466 9372
rect -28530 9228 -28466 9292
rect -28530 9148 -28466 9212
rect -28530 9068 -28466 9132
rect -28530 8988 -28466 9052
rect -28530 8908 -28466 8972
rect -28530 8828 -28466 8892
rect -28530 8748 -28466 8812
rect -28530 8668 -28466 8732
rect -28530 8588 -28466 8652
rect -28530 8508 -28466 8572
rect -28530 8428 -28466 8492
rect -28530 8348 -28466 8412
rect -28530 8268 -28466 8332
rect -28530 8188 -28466 8252
rect -28530 8108 -28466 8172
rect -28530 8028 -28466 8092
rect -28530 7948 -28466 8012
rect -28530 7868 -28466 7932
rect -28530 7788 -28466 7852
rect -28530 7708 -28466 7772
rect -28530 7628 -28466 7692
rect -28530 7548 -28466 7612
rect -28530 7468 -28466 7532
rect -28530 7388 -28466 7452
rect -28530 7308 -28466 7372
rect -28530 7228 -28466 7292
rect -28530 7148 -28466 7212
rect -28530 7068 -28466 7132
rect -28530 6988 -28466 7052
rect -28530 6908 -28466 6972
rect -28530 6828 -28466 6892
rect -28530 6748 -28466 6812
rect -28530 6668 -28466 6732
rect -28530 6588 -28466 6652
rect -28530 6508 -28466 6572
rect -28530 6428 -28466 6492
rect -28530 6348 -28466 6412
rect -28530 6268 -28466 6332
rect -28530 6188 -28466 6252
rect -28530 6108 -28466 6172
rect -28530 6028 -28466 6092
rect -28530 5948 -28466 6012
rect -28530 5868 -28466 5932
rect -28530 5788 -28466 5852
rect -28530 5708 -28466 5772
rect -28530 5628 -28466 5692
rect -28530 5548 -28466 5612
rect -28530 5468 -28466 5532
rect -28530 5388 -28466 5452
rect -28530 5308 -28466 5372
rect -28530 5228 -28466 5292
rect -28530 5148 -28466 5212
rect -28530 5068 -28466 5132
rect -28530 4988 -28466 5052
rect -28530 4908 -28466 4972
rect -28530 4828 -28466 4892
rect -28530 4748 -28466 4812
rect -28530 4668 -28466 4732
rect -28530 4588 -28466 4652
rect -28530 4508 -28466 4572
rect -28530 4428 -28466 4492
rect -28530 4348 -28466 4412
rect -28530 4268 -28466 4332
rect -28530 4188 -28466 4252
rect -28530 4108 -28466 4172
rect -28530 4028 -28466 4092
rect -28530 3948 -28466 4012
rect -28530 3868 -28466 3932
rect -28530 3788 -28466 3852
rect -28530 3708 -28466 3772
rect -28530 3628 -28466 3692
rect -28530 3548 -28466 3612
rect -28530 3468 -28466 3532
rect -28530 3388 -28466 3452
rect -28530 3308 -28466 3372
rect -28530 3228 -28466 3292
rect -22211 9308 -22147 9372
rect -22211 9228 -22147 9292
rect -22211 9148 -22147 9212
rect -22211 9068 -22147 9132
rect -22211 8988 -22147 9052
rect -22211 8908 -22147 8972
rect -22211 8828 -22147 8892
rect -22211 8748 -22147 8812
rect -22211 8668 -22147 8732
rect -22211 8588 -22147 8652
rect -22211 8508 -22147 8572
rect -22211 8428 -22147 8492
rect -22211 8348 -22147 8412
rect -22211 8268 -22147 8332
rect -22211 8188 -22147 8252
rect -22211 8108 -22147 8172
rect -22211 8028 -22147 8092
rect -22211 7948 -22147 8012
rect -22211 7868 -22147 7932
rect -22211 7788 -22147 7852
rect -22211 7708 -22147 7772
rect -22211 7628 -22147 7692
rect -22211 7548 -22147 7612
rect -22211 7468 -22147 7532
rect -22211 7388 -22147 7452
rect -22211 7308 -22147 7372
rect -22211 7228 -22147 7292
rect -22211 7148 -22147 7212
rect -22211 7068 -22147 7132
rect -22211 6988 -22147 7052
rect -22211 6908 -22147 6972
rect -22211 6828 -22147 6892
rect -22211 6748 -22147 6812
rect -22211 6668 -22147 6732
rect -22211 6588 -22147 6652
rect -22211 6508 -22147 6572
rect -22211 6428 -22147 6492
rect -22211 6348 -22147 6412
rect -22211 6268 -22147 6332
rect -22211 6188 -22147 6252
rect -22211 6108 -22147 6172
rect -22211 6028 -22147 6092
rect -22211 5948 -22147 6012
rect -22211 5868 -22147 5932
rect -22211 5788 -22147 5852
rect -22211 5708 -22147 5772
rect -22211 5628 -22147 5692
rect -22211 5548 -22147 5612
rect -22211 5468 -22147 5532
rect -22211 5388 -22147 5452
rect -22211 5308 -22147 5372
rect -22211 5228 -22147 5292
rect -22211 5148 -22147 5212
rect -22211 5068 -22147 5132
rect -22211 4988 -22147 5052
rect -22211 4908 -22147 4972
rect -22211 4828 -22147 4892
rect -22211 4748 -22147 4812
rect -22211 4668 -22147 4732
rect -22211 4588 -22147 4652
rect -22211 4508 -22147 4572
rect -22211 4428 -22147 4492
rect -22211 4348 -22147 4412
rect -22211 4268 -22147 4332
rect -22211 4188 -22147 4252
rect -22211 4108 -22147 4172
rect -22211 4028 -22147 4092
rect -22211 3948 -22147 4012
rect -22211 3868 -22147 3932
rect -22211 3788 -22147 3852
rect -22211 3708 -22147 3772
rect -22211 3628 -22147 3692
rect -22211 3548 -22147 3612
rect -22211 3468 -22147 3532
rect -22211 3388 -22147 3452
rect -22211 3308 -22147 3372
rect -22211 3228 -22147 3292
rect -15892 9308 -15828 9372
rect -15892 9228 -15828 9292
rect -15892 9148 -15828 9212
rect -15892 9068 -15828 9132
rect -15892 8988 -15828 9052
rect -15892 8908 -15828 8972
rect -15892 8828 -15828 8892
rect -15892 8748 -15828 8812
rect -15892 8668 -15828 8732
rect -15892 8588 -15828 8652
rect -15892 8508 -15828 8572
rect -15892 8428 -15828 8492
rect -15892 8348 -15828 8412
rect -15892 8268 -15828 8332
rect -15892 8188 -15828 8252
rect -15892 8108 -15828 8172
rect -15892 8028 -15828 8092
rect -15892 7948 -15828 8012
rect -15892 7868 -15828 7932
rect -15892 7788 -15828 7852
rect -15892 7708 -15828 7772
rect -15892 7628 -15828 7692
rect -15892 7548 -15828 7612
rect -15892 7468 -15828 7532
rect -15892 7388 -15828 7452
rect -15892 7308 -15828 7372
rect -15892 7228 -15828 7292
rect -15892 7148 -15828 7212
rect -15892 7068 -15828 7132
rect -15892 6988 -15828 7052
rect -15892 6908 -15828 6972
rect -15892 6828 -15828 6892
rect -15892 6748 -15828 6812
rect -15892 6668 -15828 6732
rect -15892 6588 -15828 6652
rect -15892 6508 -15828 6572
rect -15892 6428 -15828 6492
rect -15892 6348 -15828 6412
rect -15892 6268 -15828 6332
rect -15892 6188 -15828 6252
rect -15892 6108 -15828 6172
rect -15892 6028 -15828 6092
rect -15892 5948 -15828 6012
rect -15892 5868 -15828 5932
rect -15892 5788 -15828 5852
rect -15892 5708 -15828 5772
rect -15892 5628 -15828 5692
rect -15892 5548 -15828 5612
rect -15892 5468 -15828 5532
rect -15892 5388 -15828 5452
rect -15892 5308 -15828 5372
rect -15892 5228 -15828 5292
rect -15892 5148 -15828 5212
rect -15892 5068 -15828 5132
rect -15892 4988 -15828 5052
rect -15892 4908 -15828 4972
rect -15892 4828 -15828 4892
rect -15892 4748 -15828 4812
rect -15892 4668 -15828 4732
rect -15892 4588 -15828 4652
rect -15892 4508 -15828 4572
rect -15892 4428 -15828 4492
rect -15892 4348 -15828 4412
rect -15892 4268 -15828 4332
rect -15892 4188 -15828 4252
rect -15892 4108 -15828 4172
rect -15892 4028 -15828 4092
rect -15892 3948 -15828 4012
rect -15892 3868 -15828 3932
rect -15892 3788 -15828 3852
rect -15892 3708 -15828 3772
rect -15892 3628 -15828 3692
rect -15892 3548 -15828 3612
rect -15892 3468 -15828 3532
rect -15892 3388 -15828 3452
rect -15892 3308 -15828 3372
rect -15892 3228 -15828 3292
rect -9573 9308 -9509 9372
rect -9573 9228 -9509 9292
rect -9573 9148 -9509 9212
rect -9573 9068 -9509 9132
rect -9573 8988 -9509 9052
rect -9573 8908 -9509 8972
rect -9573 8828 -9509 8892
rect -9573 8748 -9509 8812
rect -9573 8668 -9509 8732
rect -9573 8588 -9509 8652
rect -9573 8508 -9509 8572
rect -9573 8428 -9509 8492
rect -9573 8348 -9509 8412
rect -9573 8268 -9509 8332
rect -9573 8188 -9509 8252
rect -9573 8108 -9509 8172
rect -9573 8028 -9509 8092
rect -9573 7948 -9509 8012
rect -9573 7868 -9509 7932
rect -9573 7788 -9509 7852
rect -9573 7708 -9509 7772
rect -9573 7628 -9509 7692
rect -9573 7548 -9509 7612
rect -9573 7468 -9509 7532
rect -9573 7388 -9509 7452
rect -9573 7308 -9509 7372
rect -9573 7228 -9509 7292
rect -9573 7148 -9509 7212
rect -9573 7068 -9509 7132
rect -9573 6988 -9509 7052
rect -9573 6908 -9509 6972
rect -9573 6828 -9509 6892
rect -9573 6748 -9509 6812
rect -9573 6668 -9509 6732
rect -9573 6588 -9509 6652
rect -9573 6508 -9509 6572
rect -9573 6428 -9509 6492
rect -9573 6348 -9509 6412
rect -9573 6268 -9509 6332
rect -9573 6188 -9509 6252
rect -9573 6108 -9509 6172
rect -9573 6028 -9509 6092
rect -9573 5948 -9509 6012
rect -9573 5868 -9509 5932
rect -9573 5788 -9509 5852
rect -9573 5708 -9509 5772
rect -9573 5628 -9509 5692
rect -9573 5548 -9509 5612
rect -9573 5468 -9509 5532
rect -9573 5388 -9509 5452
rect -9573 5308 -9509 5372
rect -9573 5228 -9509 5292
rect -9573 5148 -9509 5212
rect -9573 5068 -9509 5132
rect -9573 4988 -9509 5052
rect -9573 4908 -9509 4972
rect -9573 4828 -9509 4892
rect -9573 4748 -9509 4812
rect -9573 4668 -9509 4732
rect -9573 4588 -9509 4652
rect -9573 4508 -9509 4572
rect -9573 4428 -9509 4492
rect -9573 4348 -9509 4412
rect -9573 4268 -9509 4332
rect -9573 4188 -9509 4252
rect -9573 4108 -9509 4172
rect -9573 4028 -9509 4092
rect -9573 3948 -9509 4012
rect -9573 3868 -9509 3932
rect -9573 3788 -9509 3852
rect -9573 3708 -9509 3772
rect -9573 3628 -9509 3692
rect -9573 3548 -9509 3612
rect -9573 3468 -9509 3532
rect -9573 3388 -9509 3452
rect -9573 3308 -9509 3372
rect -9573 3228 -9509 3292
rect -3254 9308 -3190 9372
rect -3254 9228 -3190 9292
rect -3254 9148 -3190 9212
rect -3254 9068 -3190 9132
rect -3254 8988 -3190 9052
rect -3254 8908 -3190 8972
rect -3254 8828 -3190 8892
rect -3254 8748 -3190 8812
rect -3254 8668 -3190 8732
rect -3254 8588 -3190 8652
rect -3254 8508 -3190 8572
rect -3254 8428 -3190 8492
rect -3254 8348 -3190 8412
rect -3254 8268 -3190 8332
rect -3254 8188 -3190 8252
rect -3254 8108 -3190 8172
rect -3254 8028 -3190 8092
rect -3254 7948 -3190 8012
rect -3254 7868 -3190 7932
rect -3254 7788 -3190 7852
rect -3254 7708 -3190 7772
rect -3254 7628 -3190 7692
rect -3254 7548 -3190 7612
rect -3254 7468 -3190 7532
rect -3254 7388 -3190 7452
rect -3254 7308 -3190 7372
rect -3254 7228 -3190 7292
rect -3254 7148 -3190 7212
rect -3254 7068 -3190 7132
rect -3254 6988 -3190 7052
rect -3254 6908 -3190 6972
rect -3254 6828 -3190 6892
rect -3254 6748 -3190 6812
rect -3254 6668 -3190 6732
rect -3254 6588 -3190 6652
rect -3254 6508 -3190 6572
rect -3254 6428 -3190 6492
rect -3254 6348 -3190 6412
rect -3254 6268 -3190 6332
rect -3254 6188 -3190 6252
rect -3254 6108 -3190 6172
rect -3254 6028 -3190 6092
rect -3254 5948 -3190 6012
rect -3254 5868 -3190 5932
rect -3254 5788 -3190 5852
rect -3254 5708 -3190 5772
rect -3254 5628 -3190 5692
rect -3254 5548 -3190 5612
rect -3254 5468 -3190 5532
rect -3254 5388 -3190 5452
rect -3254 5308 -3190 5372
rect -3254 5228 -3190 5292
rect -3254 5148 -3190 5212
rect -3254 5068 -3190 5132
rect -3254 4988 -3190 5052
rect -3254 4908 -3190 4972
rect -3254 4828 -3190 4892
rect -3254 4748 -3190 4812
rect -3254 4668 -3190 4732
rect -3254 4588 -3190 4652
rect -3254 4508 -3190 4572
rect -3254 4428 -3190 4492
rect -3254 4348 -3190 4412
rect -3254 4268 -3190 4332
rect -3254 4188 -3190 4252
rect -3254 4108 -3190 4172
rect -3254 4028 -3190 4092
rect -3254 3948 -3190 4012
rect -3254 3868 -3190 3932
rect -3254 3788 -3190 3852
rect -3254 3708 -3190 3772
rect -3254 3628 -3190 3692
rect -3254 3548 -3190 3612
rect -3254 3468 -3190 3532
rect -3254 3388 -3190 3452
rect -3254 3308 -3190 3372
rect -3254 3228 -3190 3292
rect 3065 9308 3129 9372
rect 3065 9228 3129 9292
rect 3065 9148 3129 9212
rect 3065 9068 3129 9132
rect 3065 8988 3129 9052
rect 3065 8908 3129 8972
rect 3065 8828 3129 8892
rect 3065 8748 3129 8812
rect 3065 8668 3129 8732
rect 3065 8588 3129 8652
rect 3065 8508 3129 8572
rect 3065 8428 3129 8492
rect 3065 8348 3129 8412
rect 3065 8268 3129 8332
rect 3065 8188 3129 8252
rect 3065 8108 3129 8172
rect 3065 8028 3129 8092
rect 3065 7948 3129 8012
rect 3065 7868 3129 7932
rect 3065 7788 3129 7852
rect 3065 7708 3129 7772
rect 3065 7628 3129 7692
rect 3065 7548 3129 7612
rect 3065 7468 3129 7532
rect 3065 7388 3129 7452
rect 3065 7308 3129 7372
rect 3065 7228 3129 7292
rect 3065 7148 3129 7212
rect 3065 7068 3129 7132
rect 3065 6988 3129 7052
rect 3065 6908 3129 6972
rect 3065 6828 3129 6892
rect 3065 6748 3129 6812
rect 3065 6668 3129 6732
rect 3065 6588 3129 6652
rect 3065 6508 3129 6572
rect 3065 6428 3129 6492
rect 3065 6348 3129 6412
rect 3065 6268 3129 6332
rect 3065 6188 3129 6252
rect 3065 6108 3129 6172
rect 3065 6028 3129 6092
rect 3065 5948 3129 6012
rect 3065 5868 3129 5932
rect 3065 5788 3129 5852
rect 3065 5708 3129 5772
rect 3065 5628 3129 5692
rect 3065 5548 3129 5612
rect 3065 5468 3129 5532
rect 3065 5388 3129 5452
rect 3065 5308 3129 5372
rect 3065 5228 3129 5292
rect 3065 5148 3129 5212
rect 3065 5068 3129 5132
rect 3065 4988 3129 5052
rect 3065 4908 3129 4972
rect 3065 4828 3129 4892
rect 3065 4748 3129 4812
rect 3065 4668 3129 4732
rect 3065 4588 3129 4652
rect 3065 4508 3129 4572
rect 3065 4428 3129 4492
rect 3065 4348 3129 4412
rect 3065 4268 3129 4332
rect 3065 4188 3129 4252
rect 3065 4108 3129 4172
rect 3065 4028 3129 4092
rect 3065 3948 3129 4012
rect 3065 3868 3129 3932
rect 3065 3788 3129 3852
rect 3065 3708 3129 3772
rect 3065 3628 3129 3692
rect 3065 3548 3129 3612
rect 3065 3468 3129 3532
rect 3065 3388 3129 3452
rect 3065 3308 3129 3372
rect 3065 3228 3129 3292
rect 9384 9308 9448 9372
rect 9384 9228 9448 9292
rect 9384 9148 9448 9212
rect 9384 9068 9448 9132
rect 9384 8988 9448 9052
rect 9384 8908 9448 8972
rect 9384 8828 9448 8892
rect 9384 8748 9448 8812
rect 9384 8668 9448 8732
rect 9384 8588 9448 8652
rect 9384 8508 9448 8572
rect 9384 8428 9448 8492
rect 9384 8348 9448 8412
rect 9384 8268 9448 8332
rect 9384 8188 9448 8252
rect 9384 8108 9448 8172
rect 9384 8028 9448 8092
rect 9384 7948 9448 8012
rect 9384 7868 9448 7932
rect 9384 7788 9448 7852
rect 9384 7708 9448 7772
rect 9384 7628 9448 7692
rect 9384 7548 9448 7612
rect 9384 7468 9448 7532
rect 9384 7388 9448 7452
rect 9384 7308 9448 7372
rect 9384 7228 9448 7292
rect 9384 7148 9448 7212
rect 9384 7068 9448 7132
rect 9384 6988 9448 7052
rect 9384 6908 9448 6972
rect 9384 6828 9448 6892
rect 9384 6748 9448 6812
rect 9384 6668 9448 6732
rect 9384 6588 9448 6652
rect 9384 6508 9448 6572
rect 9384 6428 9448 6492
rect 9384 6348 9448 6412
rect 9384 6268 9448 6332
rect 9384 6188 9448 6252
rect 9384 6108 9448 6172
rect 9384 6028 9448 6092
rect 9384 5948 9448 6012
rect 9384 5868 9448 5932
rect 9384 5788 9448 5852
rect 9384 5708 9448 5772
rect 9384 5628 9448 5692
rect 9384 5548 9448 5612
rect 9384 5468 9448 5532
rect 9384 5388 9448 5452
rect 9384 5308 9448 5372
rect 9384 5228 9448 5292
rect 9384 5148 9448 5212
rect 9384 5068 9448 5132
rect 9384 4988 9448 5052
rect 9384 4908 9448 4972
rect 9384 4828 9448 4892
rect 9384 4748 9448 4812
rect 9384 4668 9448 4732
rect 9384 4588 9448 4652
rect 9384 4508 9448 4572
rect 9384 4428 9448 4492
rect 9384 4348 9448 4412
rect 9384 4268 9448 4332
rect 9384 4188 9448 4252
rect 9384 4108 9448 4172
rect 9384 4028 9448 4092
rect 9384 3948 9448 4012
rect 9384 3868 9448 3932
rect 9384 3788 9448 3852
rect 9384 3708 9448 3772
rect 9384 3628 9448 3692
rect 9384 3548 9448 3612
rect 9384 3468 9448 3532
rect 9384 3388 9448 3452
rect 9384 3308 9448 3372
rect 9384 3228 9448 3292
rect 15703 9308 15767 9372
rect 15703 9228 15767 9292
rect 15703 9148 15767 9212
rect 15703 9068 15767 9132
rect 15703 8988 15767 9052
rect 15703 8908 15767 8972
rect 15703 8828 15767 8892
rect 15703 8748 15767 8812
rect 15703 8668 15767 8732
rect 15703 8588 15767 8652
rect 15703 8508 15767 8572
rect 15703 8428 15767 8492
rect 15703 8348 15767 8412
rect 15703 8268 15767 8332
rect 15703 8188 15767 8252
rect 15703 8108 15767 8172
rect 15703 8028 15767 8092
rect 15703 7948 15767 8012
rect 15703 7868 15767 7932
rect 15703 7788 15767 7852
rect 15703 7708 15767 7772
rect 15703 7628 15767 7692
rect 15703 7548 15767 7612
rect 15703 7468 15767 7532
rect 15703 7388 15767 7452
rect 15703 7308 15767 7372
rect 15703 7228 15767 7292
rect 15703 7148 15767 7212
rect 15703 7068 15767 7132
rect 15703 6988 15767 7052
rect 15703 6908 15767 6972
rect 15703 6828 15767 6892
rect 15703 6748 15767 6812
rect 15703 6668 15767 6732
rect 15703 6588 15767 6652
rect 15703 6508 15767 6572
rect 15703 6428 15767 6492
rect 15703 6348 15767 6412
rect 15703 6268 15767 6332
rect 15703 6188 15767 6252
rect 15703 6108 15767 6172
rect 15703 6028 15767 6092
rect 15703 5948 15767 6012
rect 15703 5868 15767 5932
rect 15703 5788 15767 5852
rect 15703 5708 15767 5772
rect 15703 5628 15767 5692
rect 15703 5548 15767 5612
rect 15703 5468 15767 5532
rect 15703 5388 15767 5452
rect 15703 5308 15767 5372
rect 15703 5228 15767 5292
rect 15703 5148 15767 5212
rect 15703 5068 15767 5132
rect 15703 4988 15767 5052
rect 15703 4908 15767 4972
rect 15703 4828 15767 4892
rect 15703 4748 15767 4812
rect 15703 4668 15767 4732
rect 15703 4588 15767 4652
rect 15703 4508 15767 4572
rect 15703 4428 15767 4492
rect 15703 4348 15767 4412
rect 15703 4268 15767 4332
rect 15703 4188 15767 4252
rect 15703 4108 15767 4172
rect 15703 4028 15767 4092
rect 15703 3948 15767 4012
rect 15703 3868 15767 3932
rect 15703 3788 15767 3852
rect 15703 3708 15767 3772
rect 15703 3628 15767 3692
rect 15703 3548 15767 3612
rect 15703 3468 15767 3532
rect 15703 3388 15767 3452
rect 15703 3308 15767 3372
rect 15703 3228 15767 3292
rect 22022 9308 22086 9372
rect 22022 9228 22086 9292
rect 22022 9148 22086 9212
rect 22022 9068 22086 9132
rect 22022 8988 22086 9052
rect 22022 8908 22086 8972
rect 22022 8828 22086 8892
rect 22022 8748 22086 8812
rect 22022 8668 22086 8732
rect 22022 8588 22086 8652
rect 22022 8508 22086 8572
rect 22022 8428 22086 8492
rect 22022 8348 22086 8412
rect 22022 8268 22086 8332
rect 22022 8188 22086 8252
rect 22022 8108 22086 8172
rect 22022 8028 22086 8092
rect 22022 7948 22086 8012
rect 22022 7868 22086 7932
rect 22022 7788 22086 7852
rect 22022 7708 22086 7772
rect 22022 7628 22086 7692
rect 22022 7548 22086 7612
rect 22022 7468 22086 7532
rect 22022 7388 22086 7452
rect 22022 7308 22086 7372
rect 22022 7228 22086 7292
rect 22022 7148 22086 7212
rect 22022 7068 22086 7132
rect 22022 6988 22086 7052
rect 22022 6908 22086 6972
rect 22022 6828 22086 6892
rect 22022 6748 22086 6812
rect 22022 6668 22086 6732
rect 22022 6588 22086 6652
rect 22022 6508 22086 6572
rect 22022 6428 22086 6492
rect 22022 6348 22086 6412
rect 22022 6268 22086 6332
rect 22022 6188 22086 6252
rect 22022 6108 22086 6172
rect 22022 6028 22086 6092
rect 22022 5948 22086 6012
rect 22022 5868 22086 5932
rect 22022 5788 22086 5852
rect 22022 5708 22086 5772
rect 22022 5628 22086 5692
rect 22022 5548 22086 5612
rect 22022 5468 22086 5532
rect 22022 5388 22086 5452
rect 22022 5308 22086 5372
rect 22022 5228 22086 5292
rect 22022 5148 22086 5212
rect 22022 5068 22086 5132
rect 22022 4988 22086 5052
rect 22022 4908 22086 4972
rect 22022 4828 22086 4892
rect 22022 4748 22086 4812
rect 22022 4668 22086 4732
rect 22022 4588 22086 4652
rect 22022 4508 22086 4572
rect 22022 4428 22086 4492
rect 22022 4348 22086 4412
rect 22022 4268 22086 4332
rect 22022 4188 22086 4252
rect 22022 4108 22086 4172
rect 22022 4028 22086 4092
rect 22022 3948 22086 4012
rect 22022 3868 22086 3932
rect 22022 3788 22086 3852
rect 22022 3708 22086 3772
rect 22022 3628 22086 3692
rect 22022 3548 22086 3612
rect 22022 3468 22086 3532
rect 22022 3388 22086 3452
rect 22022 3308 22086 3372
rect 22022 3228 22086 3292
rect 28341 9308 28405 9372
rect 28341 9228 28405 9292
rect 28341 9148 28405 9212
rect 28341 9068 28405 9132
rect 28341 8988 28405 9052
rect 28341 8908 28405 8972
rect 28341 8828 28405 8892
rect 28341 8748 28405 8812
rect 28341 8668 28405 8732
rect 28341 8588 28405 8652
rect 28341 8508 28405 8572
rect 28341 8428 28405 8492
rect 28341 8348 28405 8412
rect 28341 8268 28405 8332
rect 28341 8188 28405 8252
rect 28341 8108 28405 8172
rect 28341 8028 28405 8092
rect 28341 7948 28405 8012
rect 28341 7868 28405 7932
rect 28341 7788 28405 7852
rect 28341 7708 28405 7772
rect 28341 7628 28405 7692
rect 28341 7548 28405 7612
rect 28341 7468 28405 7532
rect 28341 7388 28405 7452
rect 28341 7308 28405 7372
rect 28341 7228 28405 7292
rect 28341 7148 28405 7212
rect 28341 7068 28405 7132
rect 28341 6988 28405 7052
rect 28341 6908 28405 6972
rect 28341 6828 28405 6892
rect 28341 6748 28405 6812
rect 28341 6668 28405 6732
rect 28341 6588 28405 6652
rect 28341 6508 28405 6572
rect 28341 6428 28405 6492
rect 28341 6348 28405 6412
rect 28341 6268 28405 6332
rect 28341 6188 28405 6252
rect 28341 6108 28405 6172
rect 28341 6028 28405 6092
rect 28341 5948 28405 6012
rect 28341 5868 28405 5932
rect 28341 5788 28405 5852
rect 28341 5708 28405 5772
rect 28341 5628 28405 5692
rect 28341 5548 28405 5612
rect 28341 5468 28405 5532
rect 28341 5388 28405 5452
rect 28341 5308 28405 5372
rect 28341 5228 28405 5292
rect 28341 5148 28405 5212
rect 28341 5068 28405 5132
rect 28341 4988 28405 5052
rect 28341 4908 28405 4972
rect 28341 4828 28405 4892
rect 28341 4748 28405 4812
rect 28341 4668 28405 4732
rect 28341 4588 28405 4652
rect 28341 4508 28405 4572
rect 28341 4428 28405 4492
rect 28341 4348 28405 4412
rect 28341 4268 28405 4332
rect 28341 4188 28405 4252
rect 28341 4108 28405 4172
rect 28341 4028 28405 4092
rect 28341 3948 28405 4012
rect 28341 3868 28405 3932
rect 28341 3788 28405 3852
rect 28341 3708 28405 3772
rect 28341 3628 28405 3692
rect 28341 3548 28405 3612
rect 28341 3468 28405 3532
rect 28341 3388 28405 3452
rect 28341 3308 28405 3372
rect 28341 3228 28405 3292
rect 34660 9308 34724 9372
rect 34660 9228 34724 9292
rect 34660 9148 34724 9212
rect 34660 9068 34724 9132
rect 34660 8988 34724 9052
rect 34660 8908 34724 8972
rect 34660 8828 34724 8892
rect 34660 8748 34724 8812
rect 34660 8668 34724 8732
rect 34660 8588 34724 8652
rect 34660 8508 34724 8572
rect 34660 8428 34724 8492
rect 34660 8348 34724 8412
rect 34660 8268 34724 8332
rect 34660 8188 34724 8252
rect 34660 8108 34724 8172
rect 34660 8028 34724 8092
rect 34660 7948 34724 8012
rect 34660 7868 34724 7932
rect 34660 7788 34724 7852
rect 34660 7708 34724 7772
rect 34660 7628 34724 7692
rect 34660 7548 34724 7612
rect 34660 7468 34724 7532
rect 34660 7388 34724 7452
rect 34660 7308 34724 7372
rect 34660 7228 34724 7292
rect 34660 7148 34724 7212
rect 34660 7068 34724 7132
rect 34660 6988 34724 7052
rect 34660 6908 34724 6972
rect 34660 6828 34724 6892
rect 34660 6748 34724 6812
rect 34660 6668 34724 6732
rect 34660 6588 34724 6652
rect 34660 6508 34724 6572
rect 34660 6428 34724 6492
rect 34660 6348 34724 6412
rect 34660 6268 34724 6332
rect 34660 6188 34724 6252
rect 34660 6108 34724 6172
rect 34660 6028 34724 6092
rect 34660 5948 34724 6012
rect 34660 5868 34724 5932
rect 34660 5788 34724 5852
rect 34660 5708 34724 5772
rect 34660 5628 34724 5692
rect 34660 5548 34724 5612
rect 34660 5468 34724 5532
rect 34660 5388 34724 5452
rect 34660 5308 34724 5372
rect 34660 5228 34724 5292
rect 34660 5148 34724 5212
rect 34660 5068 34724 5132
rect 34660 4988 34724 5052
rect 34660 4908 34724 4972
rect 34660 4828 34724 4892
rect 34660 4748 34724 4812
rect 34660 4668 34724 4732
rect 34660 4588 34724 4652
rect 34660 4508 34724 4572
rect 34660 4428 34724 4492
rect 34660 4348 34724 4412
rect 34660 4268 34724 4332
rect 34660 4188 34724 4252
rect 34660 4108 34724 4172
rect 34660 4028 34724 4092
rect 34660 3948 34724 4012
rect 34660 3868 34724 3932
rect 34660 3788 34724 3852
rect 34660 3708 34724 3772
rect 34660 3628 34724 3692
rect 34660 3548 34724 3612
rect 34660 3468 34724 3532
rect 34660 3388 34724 3452
rect 34660 3308 34724 3372
rect 34660 3228 34724 3292
rect 40979 9308 41043 9372
rect 40979 9228 41043 9292
rect 40979 9148 41043 9212
rect 40979 9068 41043 9132
rect 40979 8988 41043 9052
rect 40979 8908 41043 8972
rect 40979 8828 41043 8892
rect 40979 8748 41043 8812
rect 40979 8668 41043 8732
rect 40979 8588 41043 8652
rect 40979 8508 41043 8572
rect 40979 8428 41043 8492
rect 40979 8348 41043 8412
rect 40979 8268 41043 8332
rect 40979 8188 41043 8252
rect 40979 8108 41043 8172
rect 40979 8028 41043 8092
rect 40979 7948 41043 8012
rect 40979 7868 41043 7932
rect 40979 7788 41043 7852
rect 40979 7708 41043 7772
rect 40979 7628 41043 7692
rect 40979 7548 41043 7612
rect 40979 7468 41043 7532
rect 40979 7388 41043 7452
rect 40979 7308 41043 7372
rect 40979 7228 41043 7292
rect 40979 7148 41043 7212
rect 40979 7068 41043 7132
rect 40979 6988 41043 7052
rect 40979 6908 41043 6972
rect 40979 6828 41043 6892
rect 40979 6748 41043 6812
rect 40979 6668 41043 6732
rect 40979 6588 41043 6652
rect 40979 6508 41043 6572
rect 40979 6428 41043 6492
rect 40979 6348 41043 6412
rect 40979 6268 41043 6332
rect 40979 6188 41043 6252
rect 40979 6108 41043 6172
rect 40979 6028 41043 6092
rect 40979 5948 41043 6012
rect 40979 5868 41043 5932
rect 40979 5788 41043 5852
rect 40979 5708 41043 5772
rect 40979 5628 41043 5692
rect 40979 5548 41043 5612
rect 40979 5468 41043 5532
rect 40979 5388 41043 5452
rect 40979 5308 41043 5372
rect 40979 5228 41043 5292
rect 40979 5148 41043 5212
rect 40979 5068 41043 5132
rect 40979 4988 41043 5052
rect 40979 4908 41043 4972
rect 40979 4828 41043 4892
rect 40979 4748 41043 4812
rect 40979 4668 41043 4732
rect 40979 4588 41043 4652
rect 40979 4508 41043 4572
rect 40979 4428 41043 4492
rect 40979 4348 41043 4412
rect 40979 4268 41043 4332
rect 40979 4188 41043 4252
rect 40979 4108 41043 4172
rect 40979 4028 41043 4092
rect 40979 3948 41043 4012
rect 40979 3868 41043 3932
rect 40979 3788 41043 3852
rect 40979 3708 41043 3772
rect 40979 3628 41043 3692
rect 40979 3548 41043 3612
rect 40979 3468 41043 3532
rect 40979 3388 41043 3452
rect 40979 3308 41043 3372
rect 40979 3228 41043 3292
rect 47298 9308 47362 9372
rect 47298 9228 47362 9292
rect 47298 9148 47362 9212
rect 47298 9068 47362 9132
rect 47298 8988 47362 9052
rect 47298 8908 47362 8972
rect 47298 8828 47362 8892
rect 47298 8748 47362 8812
rect 47298 8668 47362 8732
rect 47298 8588 47362 8652
rect 47298 8508 47362 8572
rect 47298 8428 47362 8492
rect 47298 8348 47362 8412
rect 47298 8268 47362 8332
rect 47298 8188 47362 8252
rect 47298 8108 47362 8172
rect 47298 8028 47362 8092
rect 47298 7948 47362 8012
rect 47298 7868 47362 7932
rect 47298 7788 47362 7852
rect 47298 7708 47362 7772
rect 47298 7628 47362 7692
rect 47298 7548 47362 7612
rect 47298 7468 47362 7532
rect 47298 7388 47362 7452
rect 47298 7308 47362 7372
rect 47298 7228 47362 7292
rect 47298 7148 47362 7212
rect 47298 7068 47362 7132
rect 47298 6988 47362 7052
rect 47298 6908 47362 6972
rect 47298 6828 47362 6892
rect 47298 6748 47362 6812
rect 47298 6668 47362 6732
rect 47298 6588 47362 6652
rect 47298 6508 47362 6572
rect 47298 6428 47362 6492
rect 47298 6348 47362 6412
rect 47298 6268 47362 6332
rect 47298 6188 47362 6252
rect 47298 6108 47362 6172
rect 47298 6028 47362 6092
rect 47298 5948 47362 6012
rect 47298 5868 47362 5932
rect 47298 5788 47362 5852
rect 47298 5708 47362 5772
rect 47298 5628 47362 5692
rect 47298 5548 47362 5612
rect 47298 5468 47362 5532
rect 47298 5388 47362 5452
rect 47298 5308 47362 5372
rect 47298 5228 47362 5292
rect 47298 5148 47362 5212
rect 47298 5068 47362 5132
rect 47298 4988 47362 5052
rect 47298 4908 47362 4972
rect 47298 4828 47362 4892
rect 47298 4748 47362 4812
rect 47298 4668 47362 4732
rect 47298 4588 47362 4652
rect 47298 4508 47362 4572
rect 47298 4428 47362 4492
rect 47298 4348 47362 4412
rect 47298 4268 47362 4332
rect 47298 4188 47362 4252
rect 47298 4108 47362 4172
rect 47298 4028 47362 4092
rect 47298 3948 47362 4012
rect 47298 3868 47362 3932
rect 47298 3788 47362 3852
rect 47298 3708 47362 3772
rect 47298 3628 47362 3692
rect 47298 3548 47362 3612
rect 47298 3468 47362 3532
rect 47298 3388 47362 3452
rect 47298 3308 47362 3372
rect 47298 3228 47362 3292
rect -41168 3008 -41104 3072
rect -41168 2928 -41104 2992
rect -41168 2848 -41104 2912
rect -41168 2768 -41104 2832
rect -41168 2688 -41104 2752
rect -41168 2608 -41104 2672
rect -41168 2528 -41104 2592
rect -41168 2448 -41104 2512
rect -41168 2368 -41104 2432
rect -41168 2288 -41104 2352
rect -41168 2208 -41104 2272
rect -41168 2128 -41104 2192
rect -41168 2048 -41104 2112
rect -41168 1968 -41104 2032
rect -41168 1888 -41104 1952
rect -41168 1808 -41104 1872
rect -41168 1728 -41104 1792
rect -41168 1648 -41104 1712
rect -41168 1568 -41104 1632
rect -41168 1488 -41104 1552
rect -41168 1408 -41104 1472
rect -41168 1328 -41104 1392
rect -41168 1248 -41104 1312
rect -41168 1168 -41104 1232
rect -41168 1088 -41104 1152
rect -41168 1008 -41104 1072
rect -41168 928 -41104 992
rect -41168 848 -41104 912
rect -41168 768 -41104 832
rect -41168 688 -41104 752
rect -41168 608 -41104 672
rect -41168 528 -41104 592
rect -41168 448 -41104 512
rect -41168 368 -41104 432
rect -41168 288 -41104 352
rect -41168 208 -41104 272
rect -41168 128 -41104 192
rect -41168 48 -41104 112
rect -41168 -32 -41104 32
rect -41168 -112 -41104 -48
rect -41168 -192 -41104 -128
rect -41168 -272 -41104 -208
rect -41168 -352 -41104 -288
rect -41168 -432 -41104 -368
rect -41168 -512 -41104 -448
rect -41168 -592 -41104 -528
rect -41168 -672 -41104 -608
rect -41168 -752 -41104 -688
rect -41168 -832 -41104 -768
rect -41168 -912 -41104 -848
rect -41168 -992 -41104 -928
rect -41168 -1072 -41104 -1008
rect -41168 -1152 -41104 -1088
rect -41168 -1232 -41104 -1168
rect -41168 -1312 -41104 -1248
rect -41168 -1392 -41104 -1328
rect -41168 -1472 -41104 -1408
rect -41168 -1552 -41104 -1488
rect -41168 -1632 -41104 -1568
rect -41168 -1712 -41104 -1648
rect -41168 -1792 -41104 -1728
rect -41168 -1872 -41104 -1808
rect -41168 -1952 -41104 -1888
rect -41168 -2032 -41104 -1968
rect -41168 -2112 -41104 -2048
rect -41168 -2192 -41104 -2128
rect -41168 -2272 -41104 -2208
rect -41168 -2352 -41104 -2288
rect -41168 -2432 -41104 -2368
rect -41168 -2512 -41104 -2448
rect -41168 -2592 -41104 -2528
rect -41168 -2672 -41104 -2608
rect -41168 -2752 -41104 -2688
rect -41168 -2832 -41104 -2768
rect -41168 -2912 -41104 -2848
rect -41168 -2992 -41104 -2928
rect -41168 -3072 -41104 -3008
rect -34849 3008 -34785 3072
rect -34849 2928 -34785 2992
rect -34849 2848 -34785 2912
rect -34849 2768 -34785 2832
rect -34849 2688 -34785 2752
rect -34849 2608 -34785 2672
rect -34849 2528 -34785 2592
rect -34849 2448 -34785 2512
rect -34849 2368 -34785 2432
rect -34849 2288 -34785 2352
rect -34849 2208 -34785 2272
rect -34849 2128 -34785 2192
rect -34849 2048 -34785 2112
rect -34849 1968 -34785 2032
rect -34849 1888 -34785 1952
rect -34849 1808 -34785 1872
rect -34849 1728 -34785 1792
rect -34849 1648 -34785 1712
rect -34849 1568 -34785 1632
rect -34849 1488 -34785 1552
rect -34849 1408 -34785 1472
rect -34849 1328 -34785 1392
rect -34849 1248 -34785 1312
rect -34849 1168 -34785 1232
rect -34849 1088 -34785 1152
rect -34849 1008 -34785 1072
rect -34849 928 -34785 992
rect -34849 848 -34785 912
rect -34849 768 -34785 832
rect -34849 688 -34785 752
rect -34849 608 -34785 672
rect -34849 528 -34785 592
rect -34849 448 -34785 512
rect -34849 368 -34785 432
rect -34849 288 -34785 352
rect -34849 208 -34785 272
rect -34849 128 -34785 192
rect -34849 48 -34785 112
rect -34849 -32 -34785 32
rect -34849 -112 -34785 -48
rect -34849 -192 -34785 -128
rect -34849 -272 -34785 -208
rect -34849 -352 -34785 -288
rect -34849 -432 -34785 -368
rect -34849 -512 -34785 -448
rect -34849 -592 -34785 -528
rect -34849 -672 -34785 -608
rect -34849 -752 -34785 -688
rect -34849 -832 -34785 -768
rect -34849 -912 -34785 -848
rect -34849 -992 -34785 -928
rect -34849 -1072 -34785 -1008
rect -34849 -1152 -34785 -1088
rect -34849 -1232 -34785 -1168
rect -34849 -1312 -34785 -1248
rect -34849 -1392 -34785 -1328
rect -34849 -1472 -34785 -1408
rect -34849 -1552 -34785 -1488
rect -34849 -1632 -34785 -1568
rect -34849 -1712 -34785 -1648
rect -34849 -1792 -34785 -1728
rect -34849 -1872 -34785 -1808
rect -34849 -1952 -34785 -1888
rect -34849 -2032 -34785 -1968
rect -34849 -2112 -34785 -2048
rect -34849 -2192 -34785 -2128
rect -34849 -2272 -34785 -2208
rect -34849 -2352 -34785 -2288
rect -34849 -2432 -34785 -2368
rect -34849 -2512 -34785 -2448
rect -34849 -2592 -34785 -2528
rect -34849 -2672 -34785 -2608
rect -34849 -2752 -34785 -2688
rect -34849 -2832 -34785 -2768
rect -34849 -2912 -34785 -2848
rect -34849 -2992 -34785 -2928
rect -34849 -3072 -34785 -3008
rect -28530 3008 -28466 3072
rect -28530 2928 -28466 2992
rect -28530 2848 -28466 2912
rect -28530 2768 -28466 2832
rect -28530 2688 -28466 2752
rect -28530 2608 -28466 2672
rect -28530 2528 -28466 2592
rect -28530 2448 -28466 2512
rect -28530 2368 -28466 2432
rect -28530 2288 -28466 2352
rect -28530 2208 -28466 2272
rect -28530 2128 -28466 2192
rect -28530 2048 -28466 2112
rect -28530 1968 -28466 2032
rect -28530 1888 -28466 1952
rect -28530 1808 -28466 1872
rect -28530 1728 -28466 1792
rect -28530 1648 -28466 1712
rect -28530 1568 -28466 1632
rect -28530 1488 -28466 1552
rect -28530 1408 -28466 1472
rect -28530 1328 -28466 1392
rect -28530 1248 -28466 1312
rect -28530 1168 -28466 1232
rect -28530 1088 -28466 1152
rect -28530 1008 -28466 1072
rect -28530 928 -28466 992
rect -28530 848 -28466 912
rect -28530 768 -28466 832
rect -28530 688 -28466 752
rect -28530 608 -28466 672
rect -28530 528 -28466 592
rect -28530 448 -28466 512
rect -28530 368 -28466 432
rect -28530 288 -28466 352
rect -28530 208 -28466 272
rect -28530 128 -28466 192
rect -28530 48 -28466 112
rect -28530 -32 -28466 32
rect -28530 -112 -28466 -48
rect -28530 -192 -28466 -128
rect -28530 -272 -28466 -208
rect -28530 -352 -28466 -288
rect -28530 -432 -28466 -368
rect -28530 -512 -28466 -448
rect -28530 -592 -28466 -528
rect -28530 -672 -28466 -608
rect -28530 -752 -28466 -688
rect -28530 -832 -28466 -768
rect -28530 -912 -28466 -848
rect -28530 -992 -28466 -928
rect -28530 -1072 -28466 -1008
rect -28530 -1152 -28466 -1088
rect -28530 -1232 -28466 -1168
rect -28530 -1312 -28466 -1248
rect -28530 -1392 -28466 -1328
rect -28530 -1472 -28466 -1408
rect -28530 -1552 -28466 -1488
rect -28530 -1632 -28466 -1568
rect -28530 -1712 -28466 -1648
rect -28530 -1792 -28466 -1728
rect -28530 -1872 -28466 -1808
rect -28530 -1952 -28466 -1888
rect -28530 -2032 -28466 -1968
rect -28530 -2112 -28466 -2048
rect -28530 -2192 -28466 -2128
rect -28530 -2272 -28466 -2208
rect -28530 -2352 -28466 -2288
rect -28530 -2432 -28466 -2368
rect -28530 -2512 -28466 -2448
rect -28530 -2592 -28466 -2528
rect -28530 -2672 -28466 -2608
rect -28530 -2752 -28466 -2688
rect -28530 -2832 -28466 -2768
rect -28530 -2912 -28466 -2848
rect -28530 -2992 -28466 -2928
rect -28530 -3072 -28466 -3008
rect -22211 3008 -22147 3072
rect -22211 2928 -22147 2992
rect -22211 2848 -22147 2912
rect -22211 2768 -22147 2832
rect -22211 2688 -22147 2752
rect -22211 2608 -22147 2672
rect -22211 2528 -22147 2592
rect -22211 2448 -22147 2512
rect -22211 2368 -22147 2432
rect -22211 2288 -22147 2352
rect -22211 2208 -22147 2272
rect -22211 2128 -22147 2192
rect -22211 2048 -22147 2112
rect -22211 1968 -22147 2032
rect -22211 1888 -22147 1952
rect -22211 1808 -22147 1872
rect -22211 1728 -22147 1792
rect -22211 1648 -22147 1712
rect -22211 1568 -22147 1632
rect -22211 1488 -22147 1552
rect -22211 1408 -22147 1472
rect -22211 1328 -22147 1392
rect -22211 1248 -22147 1312
rect -22211 1168 -22147 1232
rect -22211 1088 -22147 1152
rect -22211 1008 -22147 1072
rect -22211 928 -22147 992
rect -22211 848 -22147 912
rect -22211 768 -22147 832
rect -22211 688 -22147 752
rect -22211 608 -22147 672
rect -22211 528 -22147 592
rect -22211 448 -22147 512
rect -22211 368 -22147 432
rect -22211 288 -22147 352
rect -22211 208 -22147 272
rect -22211 128 -22147 192
rect -22211 48 -22147 112
rect -22211 -32 -22147 32
rect -22211 -112 -22147 -48
rect -22211 -192 -22147 -128
rect -22211 -272 -22147 -208
rect -22211 -352 -22147 -288
rect -22211 -432 -22147 -368
rect -22211 -512 -22147 -448
rect -22211 -592 -22147 -528
rect -22211 -672 -22147 -608
rect -22211 -752 -22147 -688
rect -22211 -832 -22147 -768
rect -22211 -912 -22147 -848
rect -22211 -992 -22147 -928
rect -22211 -1072 -22147 -1008
rect -22211 -1152 -22147 -1088
rect -22211 -1232 -22147 -1168
rect -22211 -1312 -22147 -1248
rect -22211 -1392 -22147 -1328
rect -22211 -1472 -22147 -1408
rect -22211 -1552 -22147 -1488
rect -22211 -1632 -22147 -1568
rect -22211 -1712 -22147 -1648
rect -22211 -1792 -22147 -1728
rect -22211 -1872 -22147 -1808
rect -22211 -1952 -22147 -1888
rect -22211 -2032 -22147 -1968
rect -22211 -2112 -22147 -2048
rect -22211 -2192 -22147 -2128
rect -22211 -2272 -22147 -2208
rect -22211 -2352 -22147 -2288
rect -22211 -2432 -22147 -2368
rect -22211 -2512 -22147 -2448
rect -22211 -2592 -22147 -2528
rect -22211 -2672 -22147 -2608
rect -22211 -2752 -22147 -2688
rect -22211 -2832 -22147 -2768
rect -22211 -2912 -22147 -2848
rect -22211 -2992 -22147 -2928
rect -22211 -3072 -22147 -3008
rect -15892 3008 -15828 3072
rect -15892 2928 -15828 2992
rect -15892 2848 -15828 2912
rect -15892 2768 -15828 2832
rect -15892 2688 -15828 2752
rect -15892 2608 -15828 2672
rect -15892 2528 -15828 2592
rect -15892 2448 -15828 2512
rect -15892 2368 -15828 2432
rect -15892 2288 -15828 2352
rect -15892 2208 -15828 2272
rect -15892 2128 -15828 2192
rect -15892 2048 -15828 2112
rect -15892 1968 -15828 2032
rect -15892 1888 -15828 1952
rect -15892 1808 -15828 1872
rect -15892 1728 -15828 1792
rect -15892 1648 -15828 1712
rect -15892 1568 -15828 1632
rect -15892 1488 -15828 1552
rect -15892 1408 -15828 1472
rect -15892 1328 -15828 1392
rect -15892 1248 -15828 1312
rect -15892 1168 -15828 1232
rect -15892 1088 -15828 1152
rect -15892 1008 -15828 1072
rect -15892 928 -15828 992
rect -15892 848 -15828 912
rect -15892 768 -15828 832
rect -15892 688 -15828 752
rect -15892 608 -15828 672
rect -15892 528 -15828 592
rect -15892 448 -15828 512
rect -15892 368 -15828 432
rect -15892 288 -15828 352
rect -15892 208 -15828 272
rect -15892 128 -15828 192
rect -15892 48 -15828 112
rect -15892 -32 -15828 32
rect -15892 -112 -15828 -48
rect -15892 -192 -15828 -128
rect -15892 -272 -15828 -208
rect -15892 -352 -15828 -288
rect -15892 -432 -15828 -368
rect -15892 -512 -15828 -448
rect -15892 -592 -15828 -528
rect -15892 -672 -15828 -608
rect -15892 -752 -15828 -688
rect -15892 -832 -15828 -768
rect -15892 -912 -15828 -848
rect -15892 -992 -15828 -928
rect -15892 -1072 -15828 -1008
rect -15892 -1152 -15828 -1088
rect -15892 -1232 -15828 -1168
rect -15892 -1312 -15828 -1248
rect -15892 -1392 -15828 -1328
rect -15892 -1472 -15828 -1408
rect -15892 -1552 -15828 -1488
rect -15892 -1632 -15828 -1568
rect -15892 -1712 -15828 -1648
rect -15892 -1792 -15828 -1728
rect -15892 -1872 -15828 -1808
rect -15892 -1952 -15828 -1888
rect -15892 -2032 -15828 -1968
rect -15892 -2112 -15828 -2048
rect -15892 -2192 -15828 -2128
rect -15892 -2272 -15828 -2208
rect -15892 -2352 -15828 -2288
rect -15892 -2432 -15828 -2368
rect -15892 -2512 -15828 -2448
rect -15892 -2592 -15828 -2528
rect -15892 -2672 -15828 -2608
rect -15892 -2752 -15828 -2688
rect -15892 -2832 -15828 -2768
rect -15892 -2912 -15828 -2848
rect -15892 -2992 -15828 -2928
rect -15892 -3072 -15828 -3008
rect -9573 3008 -9509 3072
rect -9573 2928 -9509 2992
rect -9573 2848 -9509 2912
rect -9573 2768 -9509 2832
rect -9573 2688 -9509 2752
rect -9573 2608 -9509 2672
rect -9573 2528 -9509 2592
rect -9573 2448 -9509 2512
rect -9573 2368 -9509 2432
rect -9573 2288 -9509 2352
rect -9573 2208 -9509 2272
rect -9573 2128 -9509 2192
rect -9573 2048 -9509 2112
rect -9573 1968 -9509 2032
rect -9573 1888 -9509 1952
rect -9573 1808 -9509 1872
rect -9573 1728 -9509 1792
rect -9573 1648 -9509 1712
rect -9573 1568 -9509 1632
rect -9573 1488 -9509 1552
rect -9573 1408 -9509 1472
rect -9573 1328 -9509 1392
rect -9573 1248 -9509 1312
rect -9573 1168 -9509 1232
rect -9573 1088 -9509 1152
rect -9573 1008 -9509 1072
rect -9573 928 -9509 992
rect -9573 848 -9509 912
rect -9573 768 -9509 832
rect -9573 688 -9509 752
rect -9573 608 -9509 672
rect -9573 528 -9509 592
rect -9573 448 -9509 512
rect -9573 368 -9509 432
rect -9573 288 -9509 352
rect -9573 208 -9509 272
rect -9573 128 -9509 192
rect -9573 48 -9509 112
rect -9573 -32 -9509 32
rect -9573 -112 -9509 -48
rect -9573 -192 -9509 -128
rect -9573 -272 -9509 -208
rect -9573 -352 -9509 -288
rect -9573 -432 -9509 -368
rect -9573 -512 -9509 -448
rect -9573 -592 -9509 -528
rect -9573 -672 -9509 -608
rect -9573 -752 -9509 -688
rect -9573 -832 -9509 -768
rect -9573 -912 -9509 -848
rect -9573 -992 -9509 -928
rect -9573 -1072 -9509 -1008
rect -9573 -1152 -9509 -1088
rect -9573 -1232 -9509 -1168
rect -9573 -1312 -9509 -1248
rect -9573 -1392 -9509 -1328
rect -9573 -1472 -9509 -1408
rect -9573 -1552 -9509 -1488
rect -9573 -1632 -9509 -1568
rect -9573 -1712 -9509 -1648
rect -9573 -1792 -9509 -1728
rect -9573 -1872 -9509 -1808
rect -9573 -1952 -9509 -1888
rect -9573 -2032 -9509 -1968
rect -9573 -2112 -9509 -2048
rect -9573 -2192 -9509 -2128
rect -9573 -2272 -9509 -2208
rect -9573 -2352 -9509 -2288
rect -9573 -2432 -9509 -2368
rect -9573 -2512 -9509 -2448
rect -9573 -2592 -9509 -2528
rect -9573 -2672 -9509 -2608
rect -9573 -2752 -9509 -2688
rect -9573 -2832 -9509 -2768
rect -9573 -2912 -9509 -2848
rect -9573 -2992 -9509 -2928
rect -9573 -3072 -9509 -3008
rect -3254 3008 -3190 3072
rect -3254 2928 -3190 2992
rect -3254 2848 -3190 2912
rect -3254 2768 -3190 2832
rect -3254 2688 -3190 2752
rect -3254 2608 -3190 2672
rect -3254 2528 -3190 2592
rect -3254 2448 -3190 2512
rect -3254 2368 -3190 2432
rect -3254 2288 -3190 2352
rect -3254 2208 -3190 2272
rect -3254 2128 -3190 2192
rect -3254 2048 -3190 2112
rect -3254 1968 -3190 2032
rect -3254 1888 -3190 1952
rect -3254 1808 -3190 1872
rect -3254 1728 -3190 1792
rect -3254 1648 -3190 1712
rect -3254 1568 -3190 1632
rect -3254 1488 -3190 1552
rect -3254 1408 -3190 1472
rect -3254 1328 -3190 1392
rect -3254 1248 -3190 1312
rect -3254 1168 -3190 1232
rect -3254 1088 -3190 1152
rect -3254 1008 -3190 1072
rect -3254 928 -3190 992
rect -3254 848 -3190 912
rect -3254 768 -3190 832
rect -3254 688 -3190 752
rect -3254 608 -3190 672
rect -3254 528 -3190 592
rect -3254 448 -3190 512
rect -3254 368 -3190 432
rect -3254 288 -3190 352
rect -3254 208 -3190 272
rect -3254 128 -3190 192
rect -3254 48 -3190 112
rect -3254 -32 -3190 32
rect -3254 -112 -3190 -48
rect -3254 -192 -3190 -128
rect -3254 -272 -3190 -208
rect -3254 -352 -3190 -288
rect -3254 -432 -3190 -368
rect -3254 -512 -3190 -448
rect -3254 -592 -3190 -528
rect -3254 -672 -3190 -608
rect -3254 -752 -3190 -688
rect -3254 -832 -3190 -768
rect -3254 -912 -3190 -848
rect -3254 -992 -3190 -928
rect -3254 -1072 -3190 -1008
rect -3254 -1152 -3190 -1088
rect -3254 -1232 -3190 -1168
rect -3254 -1312 -3190 -1248
rect -3254 -1392 -3190 -1328
rect -3254 -1472 -3190 -1408
rect -3254 -1552 -3190 -1488
rect -3254 -1632 -3190 -1568
rect -3254 -1712 -3190 -1648
rect -3254 -1792 -3190 -1728
rect -3254 -1872 -3190 -1808
rect -3254 -1952 -3190 -1888
rect -3254 -2032 -3190 -1968
rect -3254 -2112 -3190 -2048
rect -3254 -2192 -3190 -2128
rect -3254 -2272 -3190 -2208
rect -3254 -2352 -3190 -2288
rect -3254 -2432 -3190 -2368
rect -3254 -2512 -3190 -2448
rect -3254 -2592 -3190 -2528
rect -3254 -2672 -3190 -2608
rect -3254 -2752 -3190 -2688
rect -3254 -2832 -3190 -2768
rect -3254 -2912 -3190 -2848
rect -3254 -2992 -3190 -2928
rect -3254 -3072 -3190 -3008
rect 3065 3008 3129 3072
rect 3065 2928 3129 2992
rect 3065 2848 3129 2912
rect 3065 2768 3129 2832
rect 3065 2688 3129 2752
rect 3065 2608 3129 2672
rect 3065 2528 3129 2592
rect 3065 2448 3129 2512
rect 3065 2368 3129 2432
rect 3065 2288 3129 2352
rect 3065 2208 3129 2272
rect 3065 2128 3129 2192
rect 3065 2048 3129 2112
rect 3065 1968 3129 2032
rect 3065 1888 3129 1952
rect 3065 1808 3129 1872
rect 3065 1728 3129 1792
rect 3065 1648 3129 1712
rect 3065 1568 3129 1632
rect 3065 1488 3129 1552
rect 3065 1408 3129 1472
rect 3065 1328 3129 1392
rect 3065 1248 3129 1312
rect 3065 1168 3129 1232
rect 3065 1088 3129 1152
rect 3065 1008 3129 1072
rect 3065 928 3129 992
rect 3065 848 3129 912
rect 3065 768 3129 832
rect 3065 688 3129 752
rect 3065 608 3129 672
rect 3065 528 3129 592
rect 3065 448 3129 512
rect 3065 368 3129 432
rect 3065 288 3129 352
rect 3065 208 3129 272
rect 3065 128 3129 192
rect 3065 48 3129 112
rect 3065 -32 3129 32
rect 3065 -112 3129 -48
rect 3065 -192 3129 -128
rect 3065 -272 3129 -208
rect 3065 -352 3129 -288
rect 3065 -432 3129 -368
rect 3065 -512 3129 -448
rect 3065 -592 3129 -528
rect 3065 -672 3129 -608
rect 3065 -752 3129 -688
rect 3065 -832 3129 -768
rect 3065 -912 3129 -848
rect 3065 -992 3129 -928
rect 3065 -1072 3129 -1008
rect 3065 -1152 3129 -1088
rect 3065 -1232 3129 -1168
rect 3065 -1312 3129 -1248
rect 3065 -1392 3129 -1328
rect 3065 -1472 3129 -1408
rect 3065 -1552 3129 -1488
rect 3065 -1632 3129 -1568
rect 3065 -1712 3129 -1648
rect 3065 -1792 3129 -1728
rect 3065 -1872 3129 -1808
rect 3065 -1952 3129 -1888
rect 3065 -2032 3129 -1968
rect 3065 -2112 3129 -2048
rect 3065 -2192 3129 -2128
rect 3065 -2272 3129 -2208
rect 3065 -2352 3129 -2288
rect 3065 -2432 3129 -2368
rect 3065 -2512 3129 -2448
rect 3065 -2592 3129 -2528
rect 3065 -2672 3129 -2608
rect 3065 -2752 3129 -2688
rect 3065 -2832 3129 -2768
rect 3065 -2912 3129 -2848
rect 3065 -2992 3129 -2928
rect 3065 -3072 3129 -3008
rect 9384 3008 9448 3072
rect 9384 2928 9448 2992
rect 9384 2848 9448 2912
rect 9384 2768 9448 2832
rect 9384 2688 9448 2752
rect 9384 2608 9448 2672
rect 9384 2528 9448 2592
rect 9384 2448 9448 2512
rect 9384 2368 9448 2432
rect 9384 2288 9448 2352
rect 9384 2208 9448 2272
rect 9384 2128 9448 2192
rect 9384 2048 9448 2112
rect 9384 1968 9448 2032
rect 9384 1888 9448 1952
rect 9384 1808 9448 1872
rect 9384 1728 9448 1792
rect 9384 1648 9448 1712
rect 9384 1568 9448 1632
rect 9384 1488 9448 1552
rect 9384 1408 9448 1472
rect 9384 1328 9448 1392
rect 9384 1248 9448 1312
rect 9384 1168 9448 1232
rect 9384 1088 9448 1152
rect 9384 1008 9448 1072
rect 9384 928 9448 992
rect 9384 848 9448 912
rect 9384 768 9448 832
rect 9384 688 9448 752
rect 9384 608 9448 672
rect 9384 528 9448 592
rect 9384 448 9448 512
rect 9384 368 9448 432
rect 9384 288 9448 352
rect 9384 208 9448 272
rect 9384 128 9448 192
rect 9384 48 9448 112
rect 9384 -32 9448 32
rect 9384 -112 9448 -48
rect 9384 -192 9448 -128
rect 9384 -272 9448 -208
rect 9384 -352 9448 -288
rect 9384 -432 9448 -368
rect 9384 -512 9448 -448
rect 9384 -592 9448 -528
rect 9384 -672 9448 -608
rect 9384 -752 9448 -688
rect 9384 -832 9448 -768
rect 9384 -912 9448 -848
rect 9384 -992 9448 -928
rect 9384 -1072 9448 -1008
rect 9384 -1152 9448 -1088
rect 9384 -1232 9448 -1168
rect 9384 -1312 9448 -1248
rect 9384 -1392 9448 -1328
rect 9384 -1472 9448 -1408
rect 9384 -1552 9448 -1488
rect 9384 -1632 9448 -1568
rect 9384 -1712 9448 -1648
rect 9384 -1792 9448 -1728
rect 9384 -1872 9448 -1808
rect 9384 -1952 9448 -1888
rect 9384 -2032 9448 -1968
rect 9384 -2112 9448 -2048
rect 9384 -2192 9448 -2128
rect 9384 -2272 9448 -2208
rect 9384 -2352 9448 -2288
rect 9384 -2432 9448 -2368
rect 9384 -2512 9448 -2448
rect 9384 -2592 9448 -2528
rect 9384 -2672 9448 -2608
rect 9384 -2752 9448 -2688
rect 9384 -2832 9448 -2768
rect 9384 -2912 9448 -2848
rect 9384 -2992 9448 -2928
rect 9384 -3072 9448 -3008
rect 15703 3008 15767 3072
rect 15703 2928 15767 2992
rect 15703 2848 15767 2912
rect 15703 2768 15767 2832
rect 15703 2688 15767 2752
rect 15703 2608 15767 2672
rect 15703 2528 15767 2592
rect 15703 2448 15767 2512
rect 15703 2368 15767 2432
rect 15703 2288 15767 2352
rect 15703 2208 15767 2272
rect 15703 2128 15767 2192
rect 15703 2048 15767 2112
rect 15703 1968 15767 2032
rect 15703 1888 15767 1952
rect 15703 1808 15767 1872
rect 15703 1728 15767 1792
rect 15703 1648 15767 1712
rect 15703 1568 15767 1632
rect 15703 1488 15767 1552
rect 15703 1408 15767 1472
rect 15703 1328 15767 1392
rect 15703 1248 15767 1312
rect 15703 1168 15767 1232
rect 15703 1088 15767 1152
rect 15703 1008 15767 1072
rect 15703 928 15767 992
rect 15703 848 15767 912
rect 15703 768 15767 832
rect 15703 688 15767 752
rect 15703 608 15767 672
rect 15703 528 15767 592
rect 15703 448 15767 512
rect 15703 368 15767 432
rect 15703 288 15767 352
rect 15703 208 15767 272
rect 15703 128 15767 192
rect 15703 48 15767 112
rect 15703 -32 15767 32
rect 15703 -112 15767 -48
rect 15703 -192 15767 -128
rect 15703 -272 15767 -208
rect 15703 -352 15767 -288
rect 15703 -432 15767 -368
rect 15703 -512 15767 -448
rect 15703 -592 15767 -528
rect 15703 -672 15767 -608
rect 15703 -752 15767 -688
rect 15703 -832 15767 -768
rect 15703 -912 15767 -848
rect 15703 -992 15767 -928
rect 15703 -1072 15767 -1008
rect 15703 -1152 15767 -1088
rect 15703 -1232 15767 -1168
rect 15703 -1312 15767 -1248
rect 15703 -1392 15767 -1328
rect 15703 -1472 15767 -1408
rect 15703 -1552 15767 -1488
rect 15703 -1632 15767 -1568
rect 15703 -1712 15767 -1648
rect 15703 -1792 15767 -1728
rect 15703 -1872 15767 -1808
rect 15703 -1952 15767 -1888
rect 15703 -2032 15767 -1968
rect 15703 -2112 15767 -2048
rect 15703 -2192 15767 -2128
rect 15703 -2272 15767 -2208
rect 15703 -2352 15767 -2288
rect 15703 -2432 15767 -2368
rect 15703 -2512 15767 -2448
rect 15703 -2592 15767 -2528
rect 15703 -2672 15767 -2608
rect 15703 -2752 15767 -2688
rect 15703 -2832 15767 -2768
rect 15703 -2912 15767 -2848
rect 15703 -2992 15767 -2928
rect 15703 -3072 15767 -3008
rect 22022 3008 22086 3072
rect 22022 2928 22086 2992
rect 22022 2848 22086 2912
rect 22022 2768 22086 2832
rect 22022 2688 22086 2752
rect 22022 2608 22086 2672
rect 22022 2528 22086 2592
rect 22022 2448 22086 2512
rect 22022 2368 22086 2432
rect 22022 2288 22086 2352
rect 22022 2208 22086 2272
rect 22022 2128 22086 2192
rect 22022 2048 22086 2112
rect 22022 1968 22086 2032
rect 22022 1888 22086 1952
rect 22022 1808 22086 1872
rect 22022 1728 22086 1792
rect 22022 1648 22086 1712
rect 22022 1568 22086 1632
rect 22022 1488 22086 1552
rect 22022 1408 22086 1472
rect 22022 1328 22086 1392
rect 22022 1248 22086 1312
rect 22022 1168 22086 1232
rect 22022 1088 22086 1152
rect 22022 1008 22086 1072
rect 22022 928 22086 992
rect 22022 848 22086 912
rect 22022 768 22086 832
rect 22022 688 22086 752
rect 22022 608 22086 672
rect 22022 528 22086 592
rect 22022 448 22086 512
rect 22022 368 22086 432
rect 22022 288 22086 352
rect 22022 208 22086 272
rect 22022 128 22086 192
rect 22022 48 22086 112
rect 22022 -32 22086 32
rect 22022 -112 22086 -48
rect 22022 -192 22086 -128
rect 22022 -272 22086 -208
rect 22022 -352 22086 -288
rect 22022 -432 22086 -368
rect 22022 -512 22086 -448
rect 22022 -592 22086 -528
rect 22022 -672 22086 -608
rect 22022 -752 22086 -688
rect 22022 -832 22086 -768
rect 22022 -912 22086 -848
rect 22022 -992 22086 -928
rect 22022 -1072 22086 -1008
rect 22022 -1152 22086 -1088
rect 22022 -1232 22086 -1168
rect 22022 -1312 22086 -1248
rect 22022 -1392 22086 -1328
rect 22022 -1472 22086 -1408
rect 22022 -1552 22086 -1488
rect 22022 -1632 22086 -1568
rect 22022 -1712 22086 -1648
rect 22022 -1792 22086 -1728
rect 22022 -1872 22086 -1808
rect 22022 -1952 22086 -1888
rect 22022 -2032 22086 -1968
rect 22022 -2112 22086 -2048
rect 22022 -2192 22086 -2128
rect 22022 -2272 22086 -2208
rect 22022 -2352 22086 -2288
rect 22022 -2432 22086 -2368
rect 22022 -2512 22086 -2448
rect 22022 -2592 22086 -2528
rect 22022 -2672 22086 -2608
rect 22022 -2752 22086 -2688
rect 22022 -2832 22086 -2768
rect 22022 -2912 22086 -2848
rect 22022 -2992 22086 -2928
rect 22022 -3072 22086 -3008
rect 28341 3008 28405 3072
rect 28341 2928 28405 2992
rect 28341 2848 28405 2912
rect 28341 2768 28405 2832
rect 28341 2688 28405 2752
rect 28341 2608 28405 2672
rect 28341 2528 28405 2592
rect 28341 2448 28405 2512
rect 28341 2368 28405 2432
rect 28341 2288 28405 2352
rect 28341 2208 28405 2272
rect 28341 2128 28405 2192
rect 28341 2048 28405 2112
rect 28341 1968 28405 2032
rect 28341 1888 28405 1952
rect 28341 1808 28405 1872
rect 28341 1728 28405 1792
rect 28341 1648 28405 1712
rect 28341 1568 28405 1632
rect 28341 1488 28405 1552
rect 28341 1408 28405 1472
rect 28341 1328 28405 1392
rect 28341 1248 28405 1312
rect 28341 1168 28405 1232
rect 28341 1088 28405 1152
rect 28341 1008 28405 1072
rect 28341 928 28405 992
rect 28341 848 28405 912
rect 28341 768 28405 832
rect 28341 688 28405 752
rect 28341 608 28405 672
rect 28341 528 28405 592
rect 28341 448 28405 512
rect 28341 368 28405 432
rect 28341 288 28405 352
rect 28341 208 28405 272
rect 28341 128 28405 192
rect 28341 48 28405 112
rect 28341 -32 28405 32
rect 28341 -112 28405 -48
rect 28341 -192 28405 -128
rect 28341 -272 28405 -208
rect 28341 -352 28405 -288
rect 28341 -432 28405 -368
rect 28341 -512 28405 -448
rect 28341 -592 28405 -528
rect 28341 -672 28405 -608
rect 28341 -752 28405 -688
rect 28341 -832 28405 -768
rect 28341 -912 28405 -848
rect 28341 -992 28405 -928
rect 28341 -1072 28405 -1008
rect 28341 -1152 28405 -1088
rect 28341 -1232 28405 -1168
rect 28341 -1312 28405 -1248
rect 28341 -1392 28405 -1328
rect 28341 -1472 28405 -1408
rect 28341 -1552 28405 -1488
rect 28341 -1632 28405 -1568
rect 28341 -1712 28405 -1648
rect 28341 -1792 28405 -1728
rect 28341 -1872 28405 -1808
rect 28341 -1952 28405 -1888
rect 28341 -2032 28405 -1968
rect 28341 -2112 28405 -2048
rect 28341 -2192 28405 -2128
rect 28341 -2272 28405 -2208
rect 28341 -2352 28405 -2288
rect 28341 -2432 28405 -2368
rect 28341 -2512 28405 -2448
rect 28341 -2592 28405 -2528
rect 28341 -2672 28405 -2608
rect 28341 -2752 28405 -2688
rect 28341 -2832 28405 -2768
rect 28341 -2912 28405 -2848
rect 28341 -2992 28405 -2928
rect 28341 -3072 28405 -3008
rect 34660 3008 34724 3072
rect 34660 2928 34724 2992
rect 34660 2848 34724 2912
rect 34660 2768 34724 2832
rect 34660 2688 34724 2752
rect 34660 2608 34724 2672
rect 34660 2528 34724 2592
rect 34660 2448 34724 2512
rect 34660 2368 34724 2432
rect 34660 2288 34724 2352
rect 34660 2208 34724 2272
rect 34660 2128 34724 2192
rect 34660 2048 34724 2112
rect 34660 1968 34724 2032
rect 34660 1888 34724 1952
rect 34660 1808 34724 1872
rect 34660 1728 34724 1792
rect 34660 1648 34724 1712
rect 34660 1568 34724 1632
rect 34660 1488 34724 1552
rect 34660 1408 34724 1472
rect 34660 1328 34724 1392
rect 34660 1248 34724 1312
rect 34660 1168 34724 1232
rect 34660 1088 34724 1152
rect 34660 1008 34724 1072
rect 34660 928 34724 992
rect 34660 848 34724 912
rect 34660 768 34724 832
rect 34660 688 34724 752
rect 34660 608 34724 672
rect 34660 528 34724 592
rect 34660 448 34724 512
rect 34660 368 34724 432
rect 34660 288 34724 352
rect 34660 208 34724 272
rect 34660 128 34724 192
rect 34660 48 34724 112
rect 34660 -32 34724 32
rect 34660 -112 34724 -48
rect 34660 -192 34724 -128
rect 34660 -272 34724 -208
rect 34660 -352 34724 -288
rect 34660 -432 34724 -368
rect 34660 -512 34724 -448
rect 34660 -592 34724 -528
rect 34660 -672 34724 -608
rect 34660 -752 34724 -688
rect 34660 -832 34724 -768
rect 34660 -912 34724 -848
rect 34660 -992 34724 -928
rect 34660 -1072 34724 -1008
rect 34660 -1152 34724 -1088
rect 34660 -1232 34724 -1168
rect 34660 -1312 34724 -1248
rect 34660 -1392 34724 -1328
rect 34660 -1472 34724 -1408
rect 34660 -1552 34724 -1488
rect 34660 -1632 34724 -1568
rect 34660 -1712 34724 -1648
rect 34660 -1792 34724 -1728
rect 34660 -1872 34724 -1808
rect 34660 -1952 34724 -1888
rect 34660 -2032 34724 -1968
rect 34660 -2112 34724 -2048
rect 34660 -2192 34724 -2128
rect 34660 -2272 34724 -2208
rect 34660 -2352 34724 -2288
rect 34660 -2432 34724 -2368
rect 34660 -2512 34724 -2448
rect 34660 -2592 34724 -2528
rect 34660 -2672 34724 -2608
rect 34660 -2752 34724 -2688
rect 34660 -2832 34724 -2768
rect 34660 -2912 34724 -2848
rect 34660 -2992 34724 -2928
rect 34660 -3072 34724 -3008
rect 40979 3008 41043 3072
rect 40979 2928 41043 2992
rect 40979 2848 41043 2912
rect 40979 2768 41043 2832
rect 40979 2688 41043 2752
rect 40979 2608 41043 2672
rect 40979 2528 41043 2592
rect 40979 2448 41043 2512
rect 40979 2368 41043 2432
rect 40979 2288 41043 2352
rect 40979 2208 41043 2272
rect 40979 2128 41043 2192
rect 40979 2048 41043 2112
rect 40979 1968 41043 2032
rect 40979 1888 41043 1952
rect 40979 1808 41043 1872
rect 40979 1728 41043 1792
rect 40979 1648 41043 1712
rect 40979 1568 41043 1632
rect 40979 1488 41043 1552
rect 40979 1408 41043 1472
rect 40979 1328 41043 1392
rect 40979 1248 41043 1312
rect 40979 1168 41043 1232
rect 40979 1088 41043 1152
rect 40979 1008 41043 1072
rect 40979 928 41043 992
rect 40979 848 41043 912
rect 40979 768 41043 832
rect 40979 688 41043 752
rect 40979 608 41043 672
rect 40979 528 41043 592
rect 40979 448 41043 512
rect 40979 368 41043 432
rect 40979 288 41043 352
rect 40979 208 41043 272
rect 40979 128 41043 192
rect 40979 48 41043 112
rect 40979 -32 41043 32
rect 40979 -112 41043 -48
rect 40979 -192 41043 -128
rect 40979 -272 41043 -208
rect 40979 -352 41043 -288
rect 40979 -432 41043 -368
rect 40979 -512 41043 -448
rect 40979 -592 41043 -528
rect 40979 -672 41043 -608
rect 40979 -752 41043 -688
rect 40979 -832 41043 -768
rect 40979 -912 41043 -848
rect 40979 -992 41043 -928
rect 40979 -1072 41043 -1008
rect 40979 -1152 41043 -1088
rect 40979 -1232 41043 -1168
rect 40979 -1312 41043 -1248
rect 40979 -1392 41043 -1328
rect 40979 -1472 41043 -1408
rect 40979 -1552 41043 -1488
rect 40979 -1632 41043 -1568
rect 40979 -1712 41043 -1648
rect 40979 -1792 41043 -1728
rect 40979 -1872 41043 -1808
rect 40979 -1952 41043 -1888
rect 40979 -2032 41043 -1968
rect 40979 -2112 41043 -2048
rect 40979 -2192 41043 -2128
rect 40979 -2272 41043 -2208
rect 40979 -2352 41043 -2288
rect 40979 -2432 41043 -2368
rect 40979 -2512 41043 -2448
rect 40979 -2592 41043 -2528
rect 40979 -2672 41043 -2608
rect 40979 -2752 41043 -2688
rect 40979 -2832 41043 -2768
rect 40979 -2912 41043 -2848
rect 40979 -2992 41043 -2928
rect 40979 -3072 41043 -3008
rect 47298 3008 47362 3072
rect 47298 2928 47362 2992
rect 47298 2848 47362 2912
rect 47298 2768 47362 2832
rect 47298 2688 47362 2752
rect 47298 2608 47362 2672
rect 47298 2528 47362 2592
rect 47298 2448 47362 2512
rect 47298 2368 47362 2432
rect 47298 2288 47362 2352
rect 47298 2208 47362 2272
rect 47298 2128 47362 2192
rect 47298 2048 47362 2112
rect 47298 1968 47362 2032
rect 47298 1888 47362 1952
rect 47298 1808 47362 1872
rect 47298 1728 47362 1792
rect 47298 1648 47362 1712
rect 47298 1568 47362 1632
rect 47298 1488 47362 1552
rect 47298 1408 47362 1472
rect 47298 1328 47362 1392
rect 47298 1248 47362 1312
rect 47298 1168 47362 1232
rect 47298 1088 47362 1152
rect 47298 1008 47362 1072
rect 47298 928 47362 992
rect 47298 848 47362 912
rect 47298 768 47362 832
rect 47298 688 47362 752
rect 47298 608 47362 672
rect 47298 528 47362 592
rect 47298 448 47362 512
rect 47298 368 47362 432
rect 47298 288 47362 352
rect 47298 208 47362 272
rect 47298 128 47362 192
rect 47298 48 47362 112
rect 47298 -32 47362 32
rect 47298 -112 47362 -48
rect 47298 -192 47362 -128
rect 47298 -272 47362 -208
rect 47298 -352 47362 -288
rect 47298 -432 47362 -368
rect 47298 -512 47362 -448
rect 47298 -592 47362 -528
rect 47298 -672 47362 -608
rect 47298 -752 47362 -688
rect 47298 -832 47362 -768
rect 47298 -912 47362 -848
rect 47298 -992 47362 -928
rect 47298 -1072 47362 -1008
rect 47298 -1152 47362 -1088
rect 47298 -1232 47362 -1168
rect 47298 -1312 47362 -1248
rect 47298 -1392 47362 -1328
rect 47298 -1472 47362 -1408
rect 47298 -1552 47362 -1488
rect 47298 -1632 47362 -1568
rect 47298 -1712 47362 -1648
rect 47298 -1792 47362 -1728
rect 47298 -1872 47362 -1808
rect 47298 -1952 47362 -1888
rect 47298 -2032 47362 -1968
rect 47298 -2112 47362 -2048
rect 47298 -2192 47362 -2128
rect 47298 -2272 47362 -2208
rect 47298 -2352 47362 -2288
rect 47298 -2432 47362 -2368
rect 47298 -2512 47362 -2448
rect 47298 -2592 47362 -2528
rect 47298 -2672 47362 -2608
rect 47298 -2752 47362 -2688
rect 47298 -2832 47362 -2768
rect 47298 -2912 47362 -2848
rect 47298 -2992 47362 -2928
rect 47298 -3072 47362 -3008
rect -41168 -3292 -41104 -3228
rect -41168 -3372 -41104 -3308
rect -41168 -3452 -41104 -3388
rect -41168 -3532 -41104 -3468
rect -41168 -3612 -41104 -3548
rect -41168 -3692 -41104 -3628
rect -41168 -3772 -41104 -3708
rect -41168 -3852 -41104 -3788
rect -41168 -3932 -41104 -3868
rect -41168 -4012 -41104 -3948
rect -41168 -4092 -41104 -4028
rect -41168 -4172 -41104 -4108
rect -41168 -4252 -41104 -4188
rect -41168 -4332 -41104 -4268
rect -41168 -4412 -41104 -4348
rect -41168 -4492 -41104 -4428
rect -41168 -4572 -41104 -4508
rect -41168 -4652 -41104 -4588
rect -41168 -4732 -41104 -4668
rect -41168 -4812 -41104 -4748
rect -41168 -4892 -41104 -4828
rect -41168 -4972 -41104 -4908
rect -41168 -5052 -41104 -4988
rect -41168 -5132 -41104 -5068
rect -41168 -5212 -41104 -5148
rect -41168 -5292 -41104 -5228
rect -41168 -5372 -41104 -5308
rect -41168 -5452 -41104 -5388
rect -41168 -5532 -41104 -5468
rect -41168 -5612 -41104 -5548
rect -41168 -5692 -41104 -5628
rect -41168 -5772 -41104 -5708
rect -41168 -5852 -41104 -5788
rect -41168 -5932 -41104 -5868
rect -41168 -6012 -41104 -5948
rect -41168 -6092 -41104 -6028
rect -41168 -6172 -41104 -6108
rect -41168 -6252 -41104 -6188
rect -41168 -6332 -41104 -6268
rect -41168 -6412 -41104 -6348
rect -41168 -6492 -41104 -6428
rect -41168 -6572 -41104 -6508
rect -41168 -6652 -41104 -6588
rect -41168 -6732 -41104 -6668
rect -41168 -6812 -41104 -6748
rect -41168 -6892 -41104 -6828
rect -41168 -6972 -41104 -6908
rect -41168 -7052 -41104 -6988
rect -41168 -7132 -41104 -7068
rect -41168 -7212 -41104 -7148
rect -41168 -7292 -41104 -7228
rect -41168 -7372 -41104 -7308
rect -41168 -7452 -41104 -7388
rect -41168 -7532 -41104 -7468
rect -41168 -7612 -41104 -7548
rect -41168 -7692 -41104 -7628
rect -41168 -7772 -41104 -7708
rect -41168 -7852 -41104 -7788
rect -41168 -7932 -41104 -7868
rect -41168 -8012 -41104 -7948
rect -41168 -8092 -41104 -8028
rect -41168 -8172 -41104 -8108
rect -41168 -8252 -41104 -8188
rect -41168 -8332 -41104 -8268
rect -41168 -8412 -41104 -8348
rect -41168 -8492 -41104 -8428
rect -41168 -8572 -41104 -8508
rect -41168 -8652 -41104 -8588
rect -41168 -8732 -41104 -8668
rect -41168 -8812 -41104 -8748
rect -41168 -8892 -41104 -8828
rect -41168 -8972 -41104 -8908
rect -41168 -9052 -41104 -8988
rect -41168 -9132 -41104 -9068
rect -41168 -9212 -41104 -9148
rect -41168 -9292 -41104 -9228
rect -41168 -9372 -41104 -9308
rect -34849 -3292 -34785 -3228
rect -34849 -3372 -34785 -3308
rect -34849 -3452 -34785 -3388
rect -34849 -3532 -34785 -3468
rect -34849 -3612 -34785 -3548
rect -34849 -3692 -34785 -3628
rect -34849 -3772 -34785 -3708
rect -34849 -3852 -34785 -3788
rect -34849 -3932 -34785 -3868
rect -34849 -4012 -34785 -3948
rect -34849 -4092 -34785 -4028
rect -34849 -4172 -34785 -4108
rect -34849 -4252 -34785 -4188
rect -34849 -4332 -34785 -4268
rect -34849 -4412 -34785 -4348
rect -34849 -4492 -34785 -4428
rect -34849 -4572 -34785 -4508
rect -34849 -4652 -34785 -4588
rect -34849 -4732 -34785 -4668
rect -34849 -4812 -34785 -4748
rect -34849 -4892 -34785 -4828
rect -34849 -4972 -34785 -4908
rect -34849 -5052 -34785 -4988
rect -34849 -5132 -34785 -5068
rect -34849 -5212 -34785 -5148
rect -34849 -5292 -34785 -5228
rect -34849 -5372 -34785 -5308
rect -34849 -5452 -34785 -5388
rect -34849 -5532 -34785 -5468
rect -34849 -5612 -34785 -5548
rect -34849 -5692 -34785 -5628
rect -34849 -5772 -34785 -5708
rect -34849 -5852 -34785 -5788
rect -34849 -5932 -34785 -5868
rect -34849 -6012 -34785 -5948
rect -34849 -6092 -34785 -6028
rect -34849 -6172 -34785 -6108
rect -34849 -6252 -34785 -6188
rect -34849 -6332 -34785 -6268
rect -34849 -6412 -34785 -6348
rect -34849 -6492 -34785 -6428
rect -34849 -6572 -34785 -6508
rect -34849 -6652 -34785 -6588
rect -34849 -6732 -34785 -6668
rect -34849 -6812 -34785 -6748
rect -34849 -6892 -34785 -6828
rect -34849 -6972 -34785 -6908
rect -34849 -7052 -34785 -6988
rect -34849 -7132 -34785 -7068
rect -34849 -7212 -34785 -7148
rect -34849 -7292 -34785 -7228
rect -34849 -7372 -34785 -7308
rect -34849 -7452 -34785 -7388
rect -34849 -7532 -34785 -7468
rect -34849 -7612 -34785 -7548
rect -34849 -7692 -34785 -7628
rect -34849 -7772 -34785 -7708
rect -34849 -7852 -34785 -7788
rect -34849 -7932 -34785 -7868
rect -34849 -8012 -34785 -7948
rect -34849 -8092 -34785 -8028
rect -34849 -8172 -34785 -8108
rect -34849 -8252 -34785 -8188
rect -34849 -8332 -34785 -8268
rect -34849 -8412 -34785 -8348
rect -34849 -8492 -34785 -8428
rect -34849 -8572 -34785 -8508
rect -34849 -8652 -34785 -8588
rect -34849 -8732 -34785 -8668
rect -34849 -8812 -34785 -8748
rect -34849 -8892 -34785 -8828
rect -34849 -8972 -34785 -8908
rect -34849 -9052 -34785 -8988
rect -34849 -9132 -34785 -9068
rect -34849 -9212 -34785 -9148
rect -34849 -9292 -34785 -9228
rect -34849 -9372 -34785 -9308
rect -28530 -3292 -28466 -3228
rect -28530 -3372 -28466 -3308
rect -28530 -3452 -28466 -3388
rect -28530 -3532 -28466 -3468
rect -28530 -3612 -28466 -3548
rect -28530 -3692 -28466 -3628
rect -28530 -3772 -28466 -3708
rect -28530 -3852 -28466 -3788
rect -28530 -3932 -28466 -3868
rect -28530 -4012 -28466 -3948
rect -28530 -4092 -28466 -4028
rect -28530 -4172 -28466 -4108
rect -28530 -4252 -28466 -4188
rect -28530 -4332 -28466 -4268
rect -28530 -4412 -28466 -4348
rect -28530 -4492 -28466 -4428
rect -28530 -4572 -28466 -4508
rect -28530 -4652 -28466 -4588
rect -28530 -4732 -28466 -4668
rect -28530 -4812 -28466 -4748
rect -28530 -4892 -28466 -4828
rect -28530 -4972 -28466 -4908
rect -28530 -5052 -28466 -4988
rect -28530 -5132 -28466 -5068
rect -28530 -5212 -28466 -5148
rect -28530 -5292 -28466 -5228
rect -28530 -5372 -28466 -5308
rect -28530 -5452 -28466 -5388
rect -28530 -5532 -28466 -5468
rect -28530 -5612 -28466 -5548
rect -28530 -5692 -28466 -5628
rect -28530 -5772 -28466 -5708
rect -28530 -5852 -28466 -5788
rect -28530 -5932 -28466 -5868
rect -28530 -6012 -28466 -5948
rect -28530 -6092 -28466 -6028
rect -28530 -6172 -28466 -6108
rect -28530 -6252 -28466 -6188
rect -28530 -6332 -28466 -6268
rect -28530 -6412 -28466 -6348
rect -28530 -6492 -28466 -6428
rect -28530 -6572 -28466 -6508
rect -28530 -6652 -28466 -6588
rect -28530 -6732 -28466 -6668
rect -28530 -6812 -28466 -6748
rect -28530 -6892 -28466 -6828
rect -28530 -6972 -28466 -6908
rect -28530 -7052 -28466 -6988
rect -28530 -7132 -28466 -7068
rect -28530 -7212 -28466 -7148
rect -28530 -7292 -28466 -7228
rect -28530 -7372 -28466 -7308
rect -28530 -7452 -28466 -7388
rect -28530 -7532 -28466 -7468
rect -28530 -7612 -28466 -7548
rect -28530 -7692 -28466 -7628
rect -28530 -7772 -28466 -7708
rect -28530 -7852 -28466 -7788
rect -28530 -7932 -28466 -7868
rect -28530 -8012 -28466 -7948
rect -28530 -8092 -28466 -8028
rect -28530 -8172 -28466 -8108
rect -28530 -8252 -28466 -8188
rect -28530 -8332 -28466 -8268
rect -28530 -8412 -28466 -8348
rect -28530 -8492 -28466 -8428
rect -28530 -8572 -28466 -8508
rect -28530 -8652 -28466 -8588
rect -28530 -8732 -28466 -8668
rect -28530 -8812 -28466 -8748
rect -28530 -8892 -28466 -8828
rect -28530 -8972 -28466 -8908
rect -28530 -9052 -28466 -8988
rect -28530 -9132 -28466 -9068
rect -28530 -9212 -28466 -9148
rect -28530 -9292 -28466 -9228
rect -28530 -9372 -28466 -9308
rect -22211 -3292 -22147 -3228
rect -22211 -3372 -22147 -3308
rect -22211 -3452 -22147 -3388
rect -22211 -3532 -22147 -3468
rect -22211 -3612 -22147 -3548
rect -22211 -3692 -22147 -3628
rect -22211 -3772 -22147 -3708
rect -22211 -3852 -22147 -3788
rect -22211 -3932 -22147 -3868
rect -22211 -4012 -22147 -3948
rect -22211 -4092 -22147 -4028
rect -22211 -4172 -22147 -4108
rect -22211 -4252 -22147 -4188
rect -22211 -4332 -22147 -4268
rect -22211 -4412 -22147 -4348
rect -22211 -4492 -22147 -4428
rect -22211 -4572 -22147 -4508
rect -22211 -4652 -22147 -4588
rect -22211 -4732 -22147 -4668
rect -22211 -4812 -22147 -4748
rect -22211 -4892 -22147 -4828
rect -22211 -4972 -22147 -4908
rect -22211 -5052 -22147 -4988
rect -22211 -5132 -22147 -5068
rect -22211 -5212 -22147 -5148
rect -22211 -5292 -22147 -5228
rect -22211 -5372 -22147 -5308
rect -22211 -5452 -22147 -5388
rect -22211 -5532 -22147 -5468
rect -22211 -5612 -22147 -5548
rect -22211 -5692 -22147 -5628
rect -22211 -5772 -22147 -5708
rect -22211 -5852 -22147 -5788
rect -22211 -5932 -22147 -5868
rect -22211 -6012 -22147 -5948
rect -22211 -6092 -22147 -6028
rect -22211 -6172 -22147 -6108
rect -22211 -6252 -22147 -6188
rect -22211 -6332 -22147 -6268
rect -22211 -6412 -22147 -6348
rect -22211 -6492 -22147 -6428
rect -22211 -6572 -22147 -6508
rect -22211 -6652 -22147 -6588
rect -22211 -6732 -22147 -6668
rect -22211 -6812 -22147 -6748
rect -22211 -6892 -22147 -6828
rect -22211 -6972 -22147 -6908
rect -22211 -7052 -22147 -6988
rect -22211 -7132 -22147 -7068
rect -22211 -7212 -22147 -7148
rect -22211 -7292 -22147 -7228
rect -22211 -7372 -22147 -7308
rect -22211 -7452 -22147 -7388
rect -22211 -7532 -22147 -7468
rect -22211 -7612 -22147 -7548
rect -22211 -7692 -22147 -7628
rect -22211 -7772 -22147 -7708
rect -22211 -7852 -22147 -7788
rect -22211 -7932 -22147 -7868
rect -22211 -8012 -22147 -7948
rect -22211 -8092 -22147 -8028
rect -22211 -8172 -22147 -8108
rect -22211 -8252 -22147 -8188
rect -22211 -8332 -22147 -8268
rect -22211 -8412 -22147 -8348
rect -22211 -8492 -22147 -8428
rect -22211 -8572 -22147 -8508
rect -22211 -8652 -22147 -8588
rect -22211 -8732 -22147 -8668
rect -22211 -8812 -22147 -8748
rect -22211 -8892 -22147 -8828
rect -22211 -8972 -22147 -8908
rect -22211 -9052 -22147 -8988
rect -22211 -9132 -22147 -9068
rect -22211 -9212 -22147 -9148
rect -22211 -9292 -22147 -9228
rect -22211 -9372 -22147 -9308
rect -15892 -3292 -15828 -3228
rect -15892 -3372 -15828 -3308
rect -15892 -3452 -15828 -3388
rect -15892 -3532 -15828 -3468
rect -15892 -3612 -15828 -3548
rect -15892 -3692 -15828 -3628
rect -15892 -3772 -15828 -3708
rect -15892 -3852 -15828 -3788
rect -15892 -3932 -15828 -3868
rect -15892 -4012 -15828 -3948
rect -15892 -4092 -15828 -4028
rect -15892 -4172 -15828 -4108
rect -15892 -4252 -15828 -4188
rect -15892 -4332 -15828 -4268
rect -15892 -4412 -15828 -4348
rect -15892 -4492 -15828 -4428
rect -15892 -4572 -15828 -4508
rect -15892 -4652 -15828 -4588
rect -15892 -4732 -15828 -4668
rect -15892 -4812 -15828 -4748
rect -15892 -4892 -15828 -4828
rect -15892 -4972 -15828 -4908
rect -15892 -5052 -15828 -4988
rect -15892 -5132 -15828 -5068
rect -15892 -5212 -15828 -5148
rect -15892 -5292 -15828 -5228
rect -15892 -5372 -15828 -5308
rect -15892 -5452 -15828 -5388
rect -15892 -5532 -15828 -5468
rect -15892 -5612 -15828 -5548
rect -15892 -5692 -15828 -5628
rect -15892 -5772 -15828 -5708
rect -15892 -5852 -15828 -5788
rect -15892 -5932 -15828 -5868
rect -15892 -6012 -15828 -5948
rect -15892 -6092 -15828 -6028
rect -15892 -6172 -15828 -6108
rect -15892 -6252 -15828 -6188
rect -15892 -6332 -15828 -6268
rect -15892 -6412 -15828 -6348
rect -15892 -6492 -15828 -6428
rect -15892 -6572 -15828 -6508
rect -15892 -6652 -15828 -6588
rect -15892 -6732 -15828 -6668
rect -15892 -6812 -15828 -6748
rect -15892 -6892 -15828 -6828
rect -15892 -6972 -15828 -6908
rect -15892 -7052 -15828 -6988
rect -15892 -7132 -15828 -7068
rect -15892 -7212 -15828 -7148
rect -15892 -7292 -15828 -7228
rect -15892 -7372 -15828 -7308
rect -15892 -7452 -15828 -7388
rect -15892 -7532 -15828 -7468
rect -15892 -7612 -15828 -7548
rect -15892 -7692 -15828 -7628
rect -15892 -7772 -15828 -7708
rect -15892 -7852 -15828 -7788
rect -15892 -7932 -15828 -7868
rect -15892 -8012 -15828 -7948
rect -15892 -8092 -15828 -8028
rect -15892 -8172 -15828 -8108
rect -15892 -8252 -15828 -8188
rect -15892 -8332 -15828 -8268
rect -15892 -8412 -15828 -8348
rect -15892 -8492 -15828 -8428
rect -15892 -8572 -15828 -8508
rect -15892 -8652 -15828 -8588
rect -15892 -8732 -15828 -8668
rect -15892 -8812 -15828 -8748
rect -15892 -8892 -15828 -8828
rect -15892 -8972 -15828 -8908
rect -15892 -9052 -15828 -8988
rect -15892 -9132 -15828 -9068
rect -15892 -9212 -15828 -9148
rect -15892 -9292 -15828 -9228
rect -15892 -9372 -15828 -9308
rect -9573 -3292 -9509 -3228
rect -9573 -3372 -9509 -3308
rect -9573 -3452 -9509 -3388
rect -9573 -3532 -9509 -3468
rect -9573 -3612 -9509 -3548
rect -9573 -3692 -9509 -3628
rect -9573 -3772 -9509 -3708
rect -9573 -3852 -9509 -3788
rect -9573 -3932 -9509 -3868
rect -9573 -4012 -9509 -3948
rect -9573 -4092 -9509 -4028
rect -9573 -4172 -9509 -4108
rect -9573 -4252 -9509 -4188
rect -9573 -4332 -9509 -4268
rect -9573 -4412 -9509 -4348
rect -9573 -4492 -9509 -4428
rect -9573 -4572 -9509 -4508
rect -9573 -4652 -9509 -4588
rect -9573 -4732 -9509 -4668
rect -9573 -4812 -9509 -4748
rect -9573 -4892 -9509 -4828
rect -9573 -4972 -9509 -4908
rect -9573 -5052 -9509 -4988
rect -9573 -5132 -9509 -5068
rect -9573 -5212 -9509 -5148
rect -9573 -5292 -9509 -5228
rect -9573 -5372 -9509 -5308
rect -9573 -5452 -9509 -5388
rect -9573 -5532 -9509 -5468
rect -9573 -5612 -9509 -5548
rect -9573 -5692 -9509 -5628
rect -9573 -5772 -9509 -5708
rect -9573 -5852 -9509 -5788
rect -9573 -5932 -9509 -5868
rect -9573 -6012 -9509 -5948
rect -9573 -6092 -9509 -6028
rect -9573 -6172 -9509 -6108
rect -9573 -6252 -9509 -6188
rect -9573 -6332 -9509 -6268
rect -9573 -6412 -9509 -6348
rect -9573 -6492 -9509 -6428
rect -9573 -6572 -9509 -6508
rect -9573 -6652 -9509 -6588
rect -9573 -6732 -9509 -6668
rect -9573 -6812 -9509 -6748
rect -9573 -6892 -9509 -6828
rect -9573 -6972 -9509 -6908
rect -9573 -7052 -9509 -6988
rect -9573 -7132 -9509 -7068
rect -9573 -7212 -9509 -7148
rect -9573 -7292 -9509 -7228
rect -9573 -7372 -9509 -7308
rect -9573 -7452 -9509 -7388
rect -9573 -7532 -9509 -7468
rect -9573 -7612 -9509 -7548
rect -9573 -7692 -9509 -7628
rect -9573 -7772 -9509 -7708
rect -9573 -7852 -9509 -7788
rect -9573 -7932 -9509 -7868
rect -9573 -8012 -9509 -7948
rect -9573 -8092 -9509 -8028
rect -9573 -8172 -9509 -8108
rect -9573 -8252 -9509 -8188
rect -9573 -8332 -9509 -8268
rect -9573 -8412 -9509 -8348
rect -9573 -8492 -9509 -8428
rect -9573 -8572 -9509 -8508
rect -9573 -8652 -9509 -8588
rect -9573 -8732 -9509 -8668
rect -9573 -8812 -9509 -8748
rect -9573 -8892 -9509 -8828
rect -9573 -8972 -9509 -8908
rect -9573 -9052 -9509 -8988
rect -9573 -9132 -9509 -9068
rect -9573 -9212 -9509 -9148
rect -9573 -9292 -9509 -9228
rect -9573 -9372 -9509 -9308
rect -3254 -3292 -3190 -3228
rect -3254 -3372 -3190 -3308
rect -3254 -3452 -3190 -3388
rect -3254 -3532 -3190 -3468
rect -3254 -3612 -3190 -3548
rect -3254 -3692 -3190 -3628
rect -3254 -3772 -3190 -3708
rect -3254 -3852 -3190 -3788
rect -3254 -3932 -3190 -3868
rect -3254 -4012 -3190 -3948
rect -3254 -4092 -3190 -4028
rect -3254 -4172 -3190 -4108
rect -3254 -4252 -3190 -4188
rect -3254 -4332 -3190 -4268
rect -3254 -4412 -3190 -4348
rect -3254 -4492 -3190 -4428
rect -3254 -4572 -3190 -4508
rect -3254 -4652 -3190 -4588
rect -3254 -4732 -3190 -4668
rect -3254 -4812 -3190 -4748
rect -3254 -4892 -3190 -4828
rect -3254 -4972 -3190 -4908
rect -3254 -5052 -3190 -4988
rect -3254 -5132 -3190 -5068
rect -3254 -5212 -3190 -5148
rect -3254 -5292 -3190 -5228
rect -3254 -5372 -3190 -5308
rect -3254 -5452 -3190 -5388
rect -3254 -5532 -3190 -5468
rect -3254 -5612 -3190 -5548
rect -3254 -5692 -3190 -5628
rect -3254 -5772 -3190 -5708
rect -3254 -5852 -3190 -5788
rect -3254 -5932 -3190 -5868
rect -3254 -6012 -3190 -5948
rect -3254 -6092 -3190 -6028
rect -3254 -6172 -3190 -6108
rect -3254 -6252 -3190 -6188
rect -3254 -6332 -3190 -6268
rect -3254 -6412 -3190 -6348
rect -3254 -6492 -3190 -6428
rect -3254 -6572 -3190 -6508
rect -3254 -6652 -3190 -6588
rect -3254 -6732 -3190 -6668
rect -3254 -6812 -3190 -6748
rect -3254 -6892 -3190 -6828
rect -3254 -6972 -3190 -6908
rect -3254 -7052 -3190 -6988
rect -3254 -7132 -3190 -7068
rect -3254 -7212 -3190 -7148
rect -3254 -7292 -3190 -7228
rect -3254 -7372 -3190 -7308
rect -3254 -7452 -3190 -7388
rect -3254 -7532 -3190 -7468
rect -3254 -7612 -3190 -7548
rect -3254 -7692 -3190 -7628
rect -3254 -7772 -3190 -7708
rect -3254 -7852 -3190 -7788
rect -3254 -7932 -3190 -7868
rect -3254 -8012 -3190 -7948
rect -3254 -8092 -3190 -8028
rect -3254 -8172 -3190 -8108
rect -3254 -8252 -3190 -8188
rect -3254 -8332 -3190 -8268
rect -3254 -8412 -3190 -8348
rect -3254 -8492 -3190 -8428
rect -3254 -8572 -3190 -8508
rect -3254 -8652 -3190 -8588
rect -3254 -8732 -3190 -8668
rect -3254 -8812 -3190 -8748
rect -3254 -8892 -3190 -8828
rect -3254 -8972 -3190 -8908
rect -3254 -9052 -3190 -8988
rect -3254 -9132 -3190 -9068
rect -3254 -9212 -3190 -9148
rect -3254 -9292 -3190 -9228
rect -3254 -9372 -3190 -9308
rect 3065 -3292 3129 -3228
rect 3065 -3372 3129 -3308
rect 3065 -3452 3129 -3388
rect 3065 -3532 3129 -3468
rect 3065 -3612 3129 -3548
rect 3065 -3692 3129 -3628
rect 3065 -3772 3129 -3708
rect 3065 -3852 3129 -3788
rect 3065 -3932 3129 -3868
rect 3065 -4012 3129 -3948
rect 3065 -4092 3129 -4028
rect 3065 -4172 3129 -4108
rect 3065 -4252 3129 -4188
rect 3065 -4332 3129 -4268
rect 3065 -4412 3129 -4348
rect 3065 -4492 3129 -4428
rect 3065 -4572 3129 -4508
rect 3065 -4652 3129 -4588
rect 3065 -4732 3129 -4668
rect 3065 -4812 3129 -4748
rect 3065 -4892 3129 -4828
rect 3065 -4972 3129 -4908
rect 3065 -5052 3129 -4988
rect 3065 -5132 3129 -5068
rect 3065 -5212 3129 -5148
rect 3065 -5292 3129 -5228
rect 3065 -5372 3129 -5308
rect 3065 -5452 3129 -5388
rect 3065 -5532 3129 -5468
rect 3065 -5612 3129 -5548
rect 3065 -5692 3129 -5628
rect 3065 -5772 3129 -5708
rect 3065 -5852 3129 -5788
rect 3065 -5932 3129 -5868
rect 3065 -6012 3129 -5948
rect 3065 -6092 3129 -6028
rect 3065 -6172 3129 -6108
rect 3065 -6252 3129 -6188
rect 3065 -6332 3129 -6268
rect 3065 -6412 3129 -6348
rect 3065 -6492 3129 -6428
rect 3065 -6572 3129 -6508
rect 3065 -6652 3129 -6588
rect 3065 -6732 3129 -6668
rect 3065 -6812 3129 -6748
rect 3065 -6892 3129 -6828
rect 3065 -6972 3129 -6908
rect 3065 -7052 3129 -6988
rect 3065 -7132 3129 -7068
rect 3065 -7212 3129 -7148
rect 3065 -7292 3129 -7228
rect 3065 -7372 3129 -7308
rect 3065 -7452 3129 -7388
rect 3065 -7532 3129 -7468
rect 3065 -7612 3129 -7548
rect 3065 -7692 3129 -7628
rect 3065 -7772 3129 -7708
rect 3065 -7852 3129 -7788
rect 3065 -7932 3129 -7868
rect 3065 -8012 3129 -7948
rect 3065 -8092 3129 -8028
rect 3065 -8172 3129 -8108
rect 3065 -8252 3129 -8188
rect 3065 -8332 3129 -8268
rect 3065 -8412 3129 -8348
rect 3065 -8492 3129 -8428
rect 3065 -8572 3129 -8508
rect 3065 -8652 3129 -8588
rect 3065 -8732 3129 -8668
rect 3065 -8812 3129 -8748
rect 3065 -8892 3129 -8828
rect 3065 -8972 3129 -8908
rect 3065 -9052 3129 -8988
rect 3065 -9132 3129 -9068
rect 3065 -9212 3129 -9148
rect 3065 -9292 3129 -9228
rect 3065 -9372 3129 -9308
rect 9384 -3292 9448 -3228
rect 9384 -3372 9448 -3308
rect 9384 -3452 9448 -3388
rect 9384 -3532 9448 -3468
rect 9384 -3612 9448 -3548
rect 9384 -3692 9448 -3628
rect 9384 -3772 9448 -3708
rect 9384 -3852 9448 -3788
rect 9384 -3932 9448 -3868
rect 9384 -4012 9448 -3948
rect 9384 -4092 9448 -4028
rect 9384 -4172 9448 -4108
rect 9384 -4252 9448 -4188
rect 9384 -4332 9448 -4268
rect 9384 -4412 9448 -4348
rect 9384 -4492 9448 -4428
rect 9384 -4572 9448 -4508
rect 9384 -4652 9448 -4588
rect 9384 -4732 9448 -4668
rect 9384 -4812 9448 -4748
rect 9384 -4892 9448 -4828
rect 9384 -4972 9448 -4908
rect 9384 -5052 9448 -4988
rect 9384 -5132 9448 -5068
rect 9384 -5212 9448 -5148
rect 9384 -5292 9448 -5228
rect 9384 -5372 9448 -5308
rect 9384 -5452 9448 -5388
rect 9384 -5532 9448 -5468
rect 9384 -5612 9448 -5548
rect 9384 -5692 9448 -5628
rect 9384 -5772 9448 -5708
rect 9384 -5852 9448 -5788
rect 9384 -5932 9448 -5868
rect 9384 -6012 9448 -5948
rect 9384 -6092 9448 -6028
rect 9384 -6172 9448 -6108
rect 9384 -6252 9448 -6188
rect 9384 -6332 9448 -6268
rect 9384 -6412 9448 -6348
rect 9384 -6492 9448 -6428
rect 9384 -6572 9448 -6508
rect 9384 -6652 9448 -6588
rect 9384 -6732 9448 -6668
rect 9384 -6812 9448 -6748
rect 9384 -6892 9448 -6828
rect 9384 -6972 9448 -6908
rect 9384 -7052 9448 -6988
rect 9384 -7132 9448 -7068
rect 9384 -7212 9448 -7148
rect 9384 -7292 9448 -7228
rect 9384 -7372 9448 -7308
rect 9384 -7452 9448 -7388
rect 9384 -7532 9448 -7468
rect 9384 -7612 9448 -7548
rect 9384 -7692 9448 -7628
rect 9384 -7772 9448 -7708
rect 9384 -7852 9448 -7788
rect 9384 -7932 9448 -7868
rect 9384 -8012 9448 -7948
rect 9384 -8092 9448 -8028
rect 9384 -8172 9448 -8108
rect 9384 -8252 9448 -8188
rect 9384 -8332 9448 -8268
rect 9384 -8412 9448 -8348
rect 9384 -8492 9448 -8428
rect 9384 -8572 9448 -8508
rect 9384 -8652 9448 -8588
rect 9384 -8732 9448 -8668
rect 9384 -8812 9448 -8748
rect 9384 -8892 9448 -8828
rect 9384 -8972 9448 -8908
rect 9384 -9052 9448 -8988
rect 9384 -9132 9448 -9068
rect 9384 -9212 9448 -9148
rect 9384 -9292 9448 -9228
rect 9384 -9372 9448 -9308
rect 15703 -3292 15767 -3228
rect 15703 -3372 15767 -3308
rect 15703 -3452 15767 -3388
rect 15703 -3532 15767 -3468
rect 15703 -3612 15767 -3548
rect 15703 -3692 15767 -3628
rect 15703 -3772 15767 -3708
rect 15703 -3852 15767 -3788
rect 15703 -3932 15767 -3868
rect 15703 -4012 15767 -3948
rect 15703 -4092 15767 -4028
rect 15703 -4172 15767 -4108
rect 15703 -4252 15767 -4188
rect 15703 -4332 15767 -4268
rect 15703 -4412 15767 -4348
rect 15703 -4492 15767 -4428
rect 15703 -4572 15767 -4508
rect 15703 -4652 15767 -4588
rect 15703 -4732 15767 -4668
rect 15703 -4812 15767 -4748
rect 15703 -4892 15767 -4828
rect 15703 -4972 15767 -4908
rect 15703 -5052 15767 -4988
rect 15703 -5132 15767 -5068
rect 15703 -5212 15767 -5148
rect 15703 -5292 15767 -5228
rect 15703 -5372 15767 -5308
rect 15703 -5452 15767 -5388
rect 15703 -5532 15767 -5468
rect 15703 -5612 15767 -5548
rect 15703 -5692 15767 -5628
rect 15703 -5772 15767 -5708
rect 15703 -5852 15767 -5788
rect 15703 -5932 15767 -5868
rect 15703 -6012 15767 -5948
rect 15703 -6092 15767 -6028
rect 15703 -6172 15767 -6108
rect 15703 -6252 15767 -6188
rect 15703 -6332 15767 -6268
rect 15703 -6412 15767 -6348
rect 15703 -6492 15767 -6428
rect 15703 -6572 15767 -6508
rect 15703 -6652 15767 -6588
rect 15703 -6732 15767 -6668
rect 15703 -6812 15767 -6748
rect 15703 -6892 15767 -6828
rect 15703 -6972 15767 -6908
rect 15703 -7052 15767 -6988
rect 15703 -7132 15767 -7068
rect 15703 -7212 15767 -7148
rect 15703 -7292 15767 -7228
rect 15703 -7372 15767 -7308
rect 15703 -7452 15767 -7388
rect 15703 -7532 15767 -7468
rect 15703 -7612 15767 -7548
rect 15703 -7692 15767 -7628
rect 15703 -7772 15767 -7708
rect 15703 -7852 15767 -7788
rect 15703 -7932 15767 -7868
rect 15703 -8012 15767 -7948
rect 15703 -8092 15767 -8028
rect 15703 -8172 15767 -8108
rect 15703 -8252 15767 -8188
rect 15703 -8332 15767 -8268
rect 15703 -8412 15767 -8348
rect 15703 -8492 15767 -8428
rect 15703 -8572 15767 -8508
rect 15703 -8652 15767 -8588
rect 15703 -8732 15767 -8668
rect 15703 -8812 15767 -8748
rect 15703 -8892 15767 -8828
rect 15703 -8972 15767 -8908
rect 15703 -9052 15767 -8988
rect 15703 -9132 15767 -9068
rect 15703 -9212 15767 -9148
rect 15703 -9292 15767 -9228
rect 15703 -9372 15767 -9308
rect 22022 -3292 22086 -3228
rect 22022 -3372 22086 -3308
rect 22022 -3452 22086 -3388
rect 22022 -3532 22086 -3468
rect 22022 -3612 22086 -3548
rect 22022 -3692 22086 -3628
rect 22022 -3772 22086 -3708
rect 22022 -3852 22086 -3788
rect 22022 -3932 22086 -3868
rect 22022 -4012 22086 -3948
rect 22022 -4092 22086 -4028
rect 22022 -4172 22086 -4108
rect 22022 -4252 22086 -4188
rect 22022 -4332 22086 -4268
rect 22022 -4412 22086 -4348
rect 22022 -4492 22086 -4428
rect 22022 -4572 22086 -4508
rect 22022 -4652 22086 -4588
rect 22022 -4732 22086 -4668
rect 22022 -4812 22086 -4748
rect 22022 -4892 22086 -4828
rect 22022 -4972 22086 -4908
rect 22022 -5052 22086 -4988
rect 22022 -5132 22086 -5068
rect 22022 -5212 22086 -5148
rect 22022 -5292 22086 -5228
rect 22022 -5372 22086 -5308
rect 22022 -5452 22086 -5388
rect 22022 -5532 22086 -5468
rect 22022 -5612 22086 -5548
rect 22022 -5692 22086 -5628
rect 22022 -5772 22086 -5708
rect 22022 -5852 22086 -5788
rect 22022 -5932 22086 -5868
rect 22022 -6012 22086 -5948
rect 22022 -6092 22086 -6028
rect 22022 -6172 22086 -6108
rect 22022 -6252 22086 -6188
rect 22022 -6332 22086 -6268
rect 22022 -6412 22086 -6348
rect 22022 -6492 22086 -6428
rect 22022 -6572 22086 -6508
rect 22022 -6652 22086 -6588
rect 22022 -6732 22086 -6668
rect 22022 -6812 22086 -6748
rect 22022 -6892 22086 -6828
rect 22022 -6972 22086 -6908
rect 22022 -7052 22086 -6988
rect 22022 -7132 22086 -7068
rect 22022 -7212 22086 -7148
rect 22022 -7292 22086 -7228
rect 22022 -7372 22086 -7308
rect 22022 -7452 22086 -7388
rect 22022 -7532 22086 -7468
rect 22022 -7612 22086 -7548
rect 22022 -7692 22086 -7628
rect 22022 -7772 22086 -7708
rect 22022 -7852 22086 -7788
rect 22022 -7932 22086 -7868
rect 22022 -8012 22086 -7948
rect 22022 -8092 22086 -8028
rect 22022 -8172 22086 -8108
rect 22022 -8252 22086 -8188
rect 22022 -8332 22086 -8268
rect 22022 -8412 22086 -8348
rect 22022 -8492 22086 -8428
rect 22022 -8572 22086 -8508
rect 22022 -8652 22086 -8588
rect 22022 -8732 22086 -8668
rect 22022 -8812 22086 -8748
rect 22022 -8892 22086 -8828
rect 22022 -8972 22086 -8908
rect 22022 -9052 22086 -8988
rect 22022 -9132 22086 -9068
rect 22022 -9212 22086 -9148
rect 22022 -9292 22086 -9228
rect 22022 -9372 22086 -9308
rect 28341 -3292 28405 -3228
rect 28341 -3372 28405 -3308
rect 28341 -3452 28405 -3388
rect 28341 -3532 28405 -3468
rect 28341 -3612 28405 -3548
rect 28341 -3692 28405 -3628
rect 28341 -3772 28405 -3708
rect 28341 -3852 28405 -3788
rect 28341 -3932 28405 -3868
rect 28341 -4012 28405 -3948
rect 28341 -4092 28405 -4028
rect 28341 -4172 28405 -4108
rect 28341 -4252 28405 -4188
rect 28341 -4332 28405 -4268
rect 28341 -4412 28405 -4348
rect 28341 -4492 28405 -4428
rect 28341 -4572 28405 -4508
rect 28341 -4652 28405 -4588
rect 28341 -4732 28405 -4668
rect 28341 -4812 28405 -4748
rect 28341 -4892 28405 -4828
rect 28341 -4972 28405 -4908
rect 28341 -5052 28405 -4988
rect 28341 -5132 28405 -5068
rect 28341 -5212 28405 -5148
rect 28341 -5292 28405 -5228
rect 28341 -5372 28405 -5308
rect 28341 -5452 28405 -5388
rect 28341 -5532 28405 -5468
rect 28341 -5612 28405 -5548
rect 28341 -5692 28405 -5628
rect 28341 -5772 28405 -5708
rect 28341 -5852 28405 -5788
rect 28341 -5932 28405 -5868
rect 28341 -6012 28405 -5948
rect 28341 -6092 28405 -6028
rect 28341 -6172 28405 -6108
rect 28341 -6252 28405 -6188
rect 28341 -6332 28405 -6268
rect 28341 -6412 28405 -6348
rect 28341 -6492 28405 -6428
rect 28341 -6572 28405 -6508
rect 28341 -6652 28405 -6588
rect 28341 -6732 28405 -6668
rect 28341 -6812 28405 -6748
rect 28341 -6892 28405 -6828
rect 28341 -6972 28405 -6908
rect 28341 -7052 28405 -6988
rect 28341 -7132 28405 -7068
rect 28341 -7212 28405 -7148
rect 28341 -7292 28405 -7228
rect 28341 -7372 28405 -7308
rect 28341 -7452 28405 -7388
rect 28341 -7532 28405 -7468
rect 28341 -7612 28405 -7548
rect 28341 -7692 28405 -7628
rect 28341 -7772 28405 -7708
rect 28341 -7852 28405 -7788
rect 28341 -7932 28405 -7868
rect 28341 -8012 28405 -7948
rect 28341 -8092 28405 -8028
rect 28341 -8172 28405 -8108
rect 28341 -8252 28405 -8188
rect 28341 -8332 28405 -8268
rect 28341 -8412 28405 -8348
rect 28341 -8492 28405 -8428
rect 28341 -8572 28405 -8508
rect 28341 -8652 28405 -8588
rect 28341 -8732 28405 -8668
rect 28341 -8812 28405 -8748
rect 28341 -8892 28405 -8828
rect 28341 -8972 28405 -8908
rect 28341 -9052 28405 -8988
rect 28341 -9132 28405 -9068
rect 28341 -9212 28405 -9148
rect 28341 -9292 28405 -9228
rect 28341 -9372 28405 -9308
rect 34660 -3292 34724 -3228
rect 34660 -3372 34724 -3308
rect 34660 -3452 34724 -3388
rect 34660 -3532 34724 -3468
rect 34660 -3612 34724 -3548
rect 34660 -3692 34724 -3628
rect 34660 -3772 34724 -3708
rect 34660 -3852 34724 -3788
rect 34660 -3932 34724 -3868
rect 34660 -4012 34724 -3948
rect 34660 -4092 34724 -4028
rect 34660 -4172 34724 -4108
rect 34660 -4252 34724 -4188
rect 34660 -4332 34724 -4268
rect 34660 -4412 34724 -4348
rect 34660 -4492 34724 -4428
rect 34660 -4572 34724 -4508
rect 34660 -4652 34724 -4588
rect 34660 -4732 34724 -4668
rect 34660 -4812 34724 -4748
rect 34660 -4892 34724 -4828
rect 34660 -4972 34724 -4908
rect 34660 -5052 34724 -4988
rect 34660 -5132 34724 -5068
rect 34660 -5212 34724 -5148
rect 34660 -5292 34724 -5228
rect 34660 -5372 34724 -5308
rect 34660 -5452 34724 -5388
rect 34660 -5532 34724 -5468
rect 34660 -5612 34724 -5548
rect 34660 -5692 34724 -5628
rect 34660 -5772 34724 -5708
rect 34660 -5852 34724 -5788
rect 34660 -5932 34724 -5868
rect 34660 -6012 34724 -5948
rect 34660 -6092 34724 -6028
rect 34660 -6172 34724 -6108
rect 34660 -6252 34724 -6188
rect 34660 -6332 34724 -6268
rect 34660 -6412 34724 -6348
rect 34660 -6492 34724 -6428
rect 34660 -6572 34724 -6508
rect 34660 -6652 34724 -6588
rect 34660 -6732 34724 -6668
rect 34660 -6812 34724 -6748
rect 34660 -6892 34724 -6828
rect 34660 -6972 34724 -6908
rect 34660 -7052 34724 -6988
rect 34660 -7132 34724 -7068
rect 34660 -7212 34724 -7148
rect 34660 -7292 34724 -7228
rect 34660 -7372 34724 -7308
rect 34660 -7452 34724 -7388
rect 34660 -7532 34724 -7468
rect 34660 -7612 34724 -7548
rect 34660 -7692 34724 -7628
rect 34660 -7772 34724 -7708
rect 34660 -7852 34724 -7788
rect 34660 -7932 34724 -7868
rect 34660 -8012 34724 -7948
rect 34660 -8092 34724 -8028
rect 34660 -8172 34724 -8108
rect 34660 -8252 34724 -8188
rect 34660 -8332 34724 -8268
rect 34660 -8412 34724 -8348
rect 34660 -8492 34724 -8428
rect 34660 -8572 34724 -8508
rect 34660 -8652 34724 -8588
rect 34660 -8732 34724 -8668
rect 34660 -8812 34724 -8748
rect 34660 -8892 34724 -8828
rect 34660 -8972 34724 -8908
rect 34660 -9052 34724 -8988
rect 34660 -9132 34724 -9068
rect 34660 -9212 34724 -9148
rect 34660 -9292 34724 -9228
rect 34660 -9372 34724 -9308
rect 40979 -3292 41043 -3228
rect 40979 -3372 41043 -3308
rect 40979 -3452 41043 -3388
rect 40979 -3532 41043 -3468
rect 40979 -3612 41043 -3548
rect 40979 -3692 41043 -3628
rect 40979 -3772 41043 -3708
rect 40979 -3852 41043 -3788
rect 40979 -3932 41043 -3868
rect 40979 -4012 41043 -3948
rect 40979 -4092 41043 -4028
rect 40979 -4172 41043 -4108
rect 40979 -4252 41043 -4188
rect 40979 -4332 41043 -4268
rect 40979 -4412 41043 -4348
rect 40979 -4492 41043 -4428
rect 40979 -4572 41043 -4508
rect 40979 -4652 41043 -4588
rect 40979 -4732 41043 -4668
rect 40979 -4812 41043 -4748
rect 40979 -4892 41043 -4828
rect 40979 -4972 41043 -4908
rect 40979 -5052 41043 -4988
rect 40979 -5132 41043 -5068
rect 40979 -5212 41043 -5148
rect 40979 -5292 41043 -5228
rect 40979 -5372 41043 -5308
rect 40979 -5452 41043 -5388
rect 40979 -5532 41043 -5468
rect 40979 -5612 41043 -5548
rect 40979 -5692 41043 -5628
rect 40979 -5772 41043 -5708
rect 40979 -5852 41043 -5788
rect 40979 -5932 41043 -5868
rect 40979 -6012 41043 -5948
rect 40979 -6092 41043 -6028
rect 40979 -6172 41043 -6108
rect 40979 -6252 41043 -6188
rect 40979 -6332 41043 -6268
rect 40979 -6412 41043 -6348
rect 40979 -6492 41043 -6428
rect 40979 -6572 41043 -6508
rect 40979 -6652 41043 -6588
rect 40979 -6732 41043 -6668
rect 40979 -6812 41043 -6748
rect 40979 -6892 41043 -6828
rect 40979 -6972 41043 -6908
rect 40979 -7052 41043 -6988
rect 40979 -7132 41043 -7068
rect 40979 -7212 41043 -7148
rect 40979 -7292 41043 -7228
rect 40979 -7372 41043 -7308
rect 40979 -7452 41043 -7388
rect 40979 -7532 41043 -7468
rect 40979 -7612 41043 -7548
rect 40979 -7692 41043 -7628
rect 40979 -7772 41043 -7708
rect 40979 -7852 41043 -7788
rect 40979 -7932 41043 -7868
rect 40979 -8012 41043 -7948
rect 40979 -8092 41043 -8028
rect 40979 -8172 41043 -8108
rect 40979 -8252 41043 -8188
rect 40979 -8332 41043 -8268
rect 40979 -8412 41043 -8348
rect 40979 -8492 41043 -8428
rect 40979 -8572 41043 -8508
rect 40979 -8652 41043 -8588
rect 40979 -8732 41043 -8668
rect 40979 -8812 41043 -8748
rect 40979 -8892 41043 -8828
rect 40979 -8972 41043 -8908
rect 40979 -9052 41043 -8988
rect 40979 -9132 41043 -9068
rect 40979 -9212 41043 -9148
rect 40979 -9292 41043 -9228
rect 40979 -9372 41043 -9308
rect 47298 -3292 47362 -3228
rect 47298 -3372 47362 -3308
rect 47298 -3452 47362 -3388
rect 47298 -3532 47362 -3468
rect 47298 -3612 47362 -3548
rect 47298 -3692 47362 -3628
rect 47298 -3772 47362 -3708
rect 47298 -3852 47362 -3788
rect 47298 -3932 47362 -3868
rect 47298 -4012 47362 -3948
rect 47298 -4092 47362 -4028
rect 47298 -4172 47362 -4108
rect 47298 -4252 47362 -4188
rect 47298 -4332 47362 -4268
rect 47298 -4412 47362 -4348
rect 47298 -4492 47362 -4428
rect 47298 -4572 47362 -4508
rect 47298 -4652 47362 -4588
rect 47298 -4732 47362 -4668
rect 47298 -4812 47362 -4748
rect 47298 -4892 47362 -4828
rect 47298 -4972 47362 -4908
rect 47298 -5052 47362 -4988
rect 47298 -5132 47362 -5068
rect 47298 -5212 47362 -5148
rect 47298 -5292 47362 -5228
rect 47298 -5372 47362 -5308
rect 47298 -5452 47362 -5388
rect 47298 -5532 47362 -5468
rect 47298 -5612 47362 -5548
rect 47298 -5692 47362 -5628
rect 47298 -5772 47362 -5708
rect 47298 -5852 47362 -5788
rect 47298 -5932 47362 -5868
rect 47298 -6012 47362 -5948
rect 47298 -6092 47362 -6028
rect 47298 -6172 47362 -6108
rect 47298 -6252 47362 -6188
rect 47298 -6332 47362 -6268
rect 47298 -6412 47362 -6348
rect 47298 -6492 47362 -6428
rect 47298 -6572 47362 -6508
rect 47298 -6652 47362 -6588
rect 47298 -6732 47362 -6668
rect 47298 -6812 47362 -6748
rect 47298 -6892 47362 -6828
rect 47298 -6972 47362 -6908
rect 47298 -7052 47362 -6988
rect 47298 -7132 47362 -7068
rect 47298 -7212 47362 -7148
rect 47298 -7292 47362 -7228
rect 47298 -7372 47362 -7308
rect 47298 -7452 47362 -7388
rect 47298 -7532 47362 -7468
rect 47298 -7612 47362 -7548
rect 47298 -7692 47362 -7628
rect 47298 -7772 47362 -7708
rect 47298 -7852 47362 -7788
rect 47298 -7932 47362 -7868
rect 47298 -8012 47362 -7948
rect 47298 -8092 47362 -8028
rect 47298 -8172 47362 -8108
rect 47298 -8252 47362 -8188
rect 47298 -8332 47362 -8268
rect 47298 -8412 47362 -8348
rect 47298 -8492 47362 -8428
rect 47298 -8572 47362 -8508
rect 47298 -8652 47362 -8588
rect 47298 -8732 47362 -8668
rect 47298 -8812 47362 -8748
rect 47298 -8892 47362 -8828
rect 47298 -8972 47362 -8908
rect 47298 -9052 47362 -8988
rect 47298 -9132 47362 -9068
rect 47298 -9212 47362 -9148
rect 47298 -9292 47362 -9228
rect 47298 -9372 47362 -9308
rect -41168 -9592 -41104 -9528
rect -41168 -9672 -41104 -9608
rect -41168 -9752 -41104 -9688
rect -41168 -9832 -41104 -9768
rect -41168 -9912 -41104 -9848
rect -41168 -9992 -41104 -9928
rect -41168 -10072 -41104 -10008
rect -41168 -10152 -41104 -10088
rect -41168 -10232 -41104 -10168
rect -41168 -10312 -41104 -10248
rect -41168 -10392 -41104 -10328
rect -41168 -10472 -41104 -10408
rect -41168 -10552 -41104 -10488
rect -41168 -10632 -41104 -10568
rect -41168 -10712 -41104 -10648
rect -41168 -10792 -41104 -10728
rect -41168 -10872 -41104 -10808
rect -41168 -10952 -41104 -10888
rect -41168 -11032 -41104 -10968
rect -41168 -11112 -41104 -11048
rect -41168 -11192 -41104 -11128
rect -41168 -11272 -41104 -11208
rect -41168 -11352 -41104 -11288
rect -41168 -11432 -41104 -11368
rect -41168 -11512 -41104 -11448
rect -41168 -11592 -41104 -11528
rect -41168 -11672 -41104 -11608
rect -41168 -11752 -41104 -11688
rect -41168 -11832 -41104 -11768
rect -41168 -11912 -41104 -11848
rect -41168 -11992 -41104 -11928
rect -41168 -12072 -41104 -12008
rect -41168 -12152 -41104 -12088
rect -41168 -12232 -41104 -12168
rect -41168 -12312 -41104 -12248
rect -41168 -12392 -41104 -12328
rect -41168 -12472 -41104 -12408
rect -41168 -12552 -41104 -12488
rect -41168 -12632 -41104 -12568
rect -41168 -12712 -41104 -12648
rect -41168 -12792 -41104 -12728
rect -41168 -12872 -41104 -12808
rect -41168 -12952 -41104 -12888
rect -41168 -13032 -41104 -12968
rect -41168 -13112 -41104 -13048
rect -41168 -13192 -41104 -13128
rect -41168 -13272 -41104 -13208
rect -41168 -13352 -41104 -13288
rect -41168 -13432 -41104 -13368
rect -41168 -13512 -41104 -13448
rect -41168 -13592 -41104 -13528
rect -41168 -13672 -41104 -13608
rect -41168 -13752 -41104 -13688
rect -41168 -13832 -41104 -13768
rect -41168 -13912 -41104 -13848
rect -41168 -13992 -41104 -13928
rect -41168 -14072 -41104 -14008
rect -41168 -14152 -41104 -14088
rect -41168 -14232 -41104 -14168
rect -41168 -14312 -41104 -14248
rect -41168 -14392 -41104 -14328
rect -41168 -14472 -41104 -14408
rect -41168 -14552 -41104 -14488
rect -41168 -14632 -41104 -14568
rect -41168 -14712 -41104 -14648
rect -41168 -14792 -41104 -14728
rect -41168 -14872 -41104 -14808
rect -41168 -14952 -41104 -14888
rect -41168 -15032 -41104 -14968
rect -41168 -15112 -41104 -15048
rect -41168 -15192 -41104 -15128
rect -41168 -15272 -41104 -15208
rect -41168 -15352 -41104 -15288
rect -41168 -15432 -41104 -15368
rect -41168 -15512 -41104 -15448
rect -41168 -15592 -41104 -15528
rect -41168 -15672 -41104 -15608
rect -34849 -9592 -34785 -9528
rect -34849 -9672 -34785 -9608
rect -34849 -9752 -34785 -9688
rect -34849 -9832 -34785 -9768
rect -34849 -9912 -34785 -9848
rect -34849 -9992 -34785 -9928
rect -34849 -10072 -34785 -10008
rect -34849 -10152 -34785 -10088
rect -34849 -10232 -34785 -10168
rect -34849 -10312 -34785 -10248
rect -34849 -10392 -34785 -10328
rect -34849 -10472 -34785 -10408
rect -34849 -10552 -34785 -10488
rect -34849 -10632 -34785 -10568
rect -34849 -10712 -34785 -10648
rect -34849 -10792 -34785 -10728
rect -34849 -10872 -34785 -10808
rect -34849 -10952 -34785 -10888
rect -34849 -11032 -34785 -10968
rect -34849 -11112 -34785 -11048
rect -34849 -11192 -34785 -11128
rect -34849 -11272 -34785 -11208
rect -34849 -11352 -34785 -11288
rect -34849 -11432 -34785 -11368
rect -34849 -11512 -34785 -11448
rect -34849 -11592 -34785 -11528
rect -34849 -11672 -34785 -11608
rect -34849 -11752 -34785 -11688
rect -34849 -11832 -34785 -11768
rect -34849 -11912 -34785 -11848
rect -34849 -11992 -34785 -11928
rect -34849 -12072 -34785 -12008
rect -34849 -12152 -34785 -12088
rect -34849 -12232 -34785 -12168
rect -34849 -12312 -34785 -12248
rect -34849 -12392 -34785 -12328
rect -34849 -12472 -34785 -12408
rect -34849 -12552 -34785 -12488
rect -34849 -12632 -34785 -12568
rect -34849 -12712 -34785 -12648
rect -34849 -12792 -34785 -12728
rect -34849 -12872 -34785 -12808
rect -34849 -12952 -34785 -12888
rect -34849 -13032 -34785 -12968
rect -34849 -13112 -34785 -13048
rect -34849 -13192 -34785 -13128
rect -34849 -13272 -34785 -13208
rect -34849 -13352 -34785 -13288
rect -34849 -13432 -34785 -13368
rect -34849 -13512 -34785 -13448
rect -34849 -13592 -34785 -13528
rect -34849 -13672 -34785 -13608
rect -34849 -13752 -34785 -13688
rect -34849 -13832 -34785 -13768
rect -34849 -13912 -34785 -13848
rect -34849 -13992 -34785 -13928
rect -34849 -14072 -34785 -14008
rect -34849 -14152 -34785 -14088
rect -34849 -14232 -34785 -14168
rect -34849 -14312 -34785 -14248
rect -34849 -14392 -34785 -14328
rect -34849 -14472 -34785 -14408
rect -34849 -14552 -34785 -14488
rect -34849 -14632 -34785 -14568
rect -34849 -14712 -34785 -14648
rect -34849 -14792 -34785 -14728
rect -34849 -14872 -34785 -14808
rect -34849 -14952 -34785 -14888
rect -34849 -15032 -34785 -14968
rect -34849 -15112 -34785 -15048
rect -34849 -15192 -34785 -15128
rect -34849 -15272 -34785 -15208
rect -34849 -15352 -34785 -15288
rect -34849 -15432 -34785 -15368
rect -34849 -15512 -34785 -15448
rect -34849 -15592 -34785 -15528
rect -34849 -15672 -34785 -15608
rect -28530 -9592 -28466 -9528
rect -28530 -9672 -28466 -9608
rect -28530 -9752 -28466 -9688
rect -28530 -9832 -28466 -9768
rect -28530 -9912 -28466 -9848
rect -28530 -9992 -28466 -9928
rect -28530 -10072 -28466 -10008
rect -28530 -10152 -28466 -10088
rect -28530 -10232 -28466 -10168
rect -28530 -10312 -28466 -10248
rect -28530 -10392 -28466 -10328
rect -28530 -10472 -28466 -10408
rect -28530 -10552 -28466 -10488
rect -28530 -10632 -28466 -10568
rect -28530 -10712 -28466 -10648
rect -28530 -10792 -28466 -10728
rect -28530 -10872 -28466 -10808
rect -28530 -10952 -28466 -10888
rect -28530 -11032 -28466 -10968
rect -28530 -11112 -28466 -11048
rect -28530 -11192 -28466 -11128
rect -28530 -11272 -28466 -11208
rect -28530 -11352 -28466 -11288
rect -28530 -11432 -28466 -11368
rect -28530 -11512 -28466 -11448
rect -28530 -11592 -28466 -11528
rect -28530 -11672 -28466 -11608
rect -28530 -11752 -28466 -11688
rect -28530 -11832 -28466 -11768
rect -28530 -11912 -28466 -11848
rect -28530 -11992 -28466 -11928
rect -28530 -12072 -28466 -12008
rect -28530 -12152 -28466 -12088
rect -28530 -12232 -28466 -12168
rect -28530 -12312 -28466 -12248
rect -28530 -12392 -28466 -12328
rect -28530 -12472 -28466 -12408
rect -28530 -12552 -28466 -12488
rect -28530 -12632 -28466 -12568
rect -28530 -12712 -28466 -12648
rect -28530 -12792 -28466 -12728
rect -28530 -12872 -28466 -12808
rect -28530 -12952 -28466 -12888
rect -28530 -13032 -28466 -12968
rect -28530 -13112 -28466 -13048
rect -28530 -13192 -28466 -13128
rect -28530 -13272 -28466 -13208
rect -28530 -13352 -28466 -13288
rect -28530 -13432 -28466 -13368
rect -28530 -13512 -28466 -13448
rect -28530 -13592 -28466 -13528
rect -28530 -13672 -28466 -13608
rect -28530 -13752 -28466 -13688
rect -28530 -13832 -28466 -13768
rect -28530 -13912 -28466 -13848
rect -28530 -13992 -28466 -13928
rect -28530 -14072 -28466 -14008
rect -28530 -14152 -28466 -14088
rect -28530 -14232 -28466 -14168
rect -28530 -14312 -28466 -14248
rect -28530 -14392 -28466 -14328
rect -28530 -14472 -28466 -14408
rect -28530 -14552 -28466 -14488
rect -28530 -14632 -28466 -14568
rect -28530 -14712 -28466 -14648
rect -28530 -14792 -28466 -14728
rect -28530 -14872 -28466 -14808
rect -28530 -14952 -28466 -14888
rect -28530 -15032 -28466 -14968
rect -28530 -15112 -28466 -15048
rect -28530 -15192 -28466 -15128
rect -28530 -15272 -28466 -15208
rect -28530 -15352 -28466 -15288
rect -28530 -15432 -28466 -15368
rect -28530 -15512 -28466 -15448
rect -28530 -15592 -28466 -15528
rect -28530 -15672 -28466 -15608
rect -22211 -9592 -22147 -9528
rect -22211 -9672 -22147 -9608
rect -22211 -9752 -22147 -9688
rect -22211 -9832 -22147 -9768
rect -22211 -9912 -22147 -9848
rect -22211 -9992 -22147 -9928
rect -22211 -10072 -22147 -10008
rect -22211 -10152 -22147 -10088
rect -22211 -10232 -22147 -10168
rect -22211 -10312 -22147 -10248
rect -22211 -10392 -22147 -10328
rect -22211 -10472 -22147 -10408
rect -22211 -10552 -22147 -10488
rect -22211 -10632 -22147 -10568
rect -22211 -10712 -22147 -10648
rect -22211 -10792 -22147 -10728
rect -22211 -10872 -22147 -10808
rect -22211 -10952 -22147 -10888
rect -22211 -11032 -22147 -10968
rect -22211 -11112 -22147 -11048
rect -22211 -11192 -22147 -11128
rect -22211 -11272 -22147 -11208
rect -22211 -11352 -22147 -11288
rect -22211 -11432 -22147 -11368
rect -22211 -11512 -22147 -11448
rect -22211 -11592 -22147 -11528
rect -22211 -11672 -22147 -11608
rect -22211 -11752 -22147 -11688
rect -22211 -11832 -22147 -11768
rect -22211 -11912 -22147 -11848
rect -22211 -11992 -22147 -11928
rect -22211 -12072 -22147 -12008
rect -22211 -12152 -22147 -12088
rect -22211 -12232 -22147 -12168
rect -22211 -12312 -22147 -12248
rect -22211 -12392 -22147 -12328
rect -22211 -12472 -22147 -12408
rect -22211 -12552 -22147 -12488
rect -22211 -12632 -22147 -12568
rect -22211 -12712 -22147 -12648
rect -22211 -12792 -22147 -12728
rect -22211 -12872 -22147 -12808
rect -22211 -12952 -22147 -12888
rect -22211 -13032 -22147 -12968
rect -22211 -13112 -22147 -13048
rect -22211 -13192 -22147 -13128
rect -22211 -13272 -22147 -13208
rect -22211 -13352 -22147 -13288
rect -22211 -13432 -22147 -13368
rect -22211 -13512 -22147 -13448
rect -22211 -13592 -22147 -13528
rect -22211 -13672 -22147 -13608
rect -22211 -13752 -22147 -13688
rect -22211 -13832 -22147 -13768
rect -22211 -13912 -22147 -13848
rect -22211 -13992 -22147 -13928
rect -22211 -14072 -22147 -14008
rect -22211 -14152 -22147 -14088
rect -22211 -14232 -22147 -14168
rect -22211 -14312 -22147 -14248
rect -22211 -14392 -22147 -14328
rect -22211 -14472 -22147 -14408
rect -22211 -14552 -22147 -14488
rect -22211 -14632 -22147 -14568
rect -22211 -14712 -22147 -14648
rect -22211 -14792 -22147 -14728
rect -22211 -14872 -22147 -14808
rect -22211 -14952 -22147 -14888
rect -22211 -15032 -22147 -14968
rect -22211 -15112 -22147 -15048
rect -22211 -15192 -22147 -15128
rect -22211 -15272 -22147 -15208
rect -22211 -15352 -22147 -15288
rect -22211 -15432 -22147 -15368
rect -22211 -15512 -22147 -15448
rect -22211 -15592 -22147 -15528
rect -22211 -15672 -22147 -15608
rect -15892 -9592 -15828 -9528
rect -15892 -9672 -15828 -9608
rect -15892 -9752 -15828 -9688
rect -15892 -9832 -15828 -9768
rect -15892 -9912 -15828 -9848
rect -15892 -9992 -15828 -9928
rect -15892 -10072 -15828 -10008
rect -15892 -10152 -15828 -10088
rect -15892 -10232 -15828 -10168
rect -15892 -10312 -15828 -10248
rect -15892 -10392 -15828 -10328
rect -15892 -10472 -15828 -10408
rect -15892 -10552 -15828 -10488
rect -15892 -10632 -15828 -10568
rect -15892 -10712 -15828 -10648
rect -15892 -10792 -15828 -10728
rect -15892 -10872 -15828 -10808
rect -15892 -10952 -15828 -10888
rect -15892 -11032 -15828 -10968
rect -15892 -11112 -15828 -11048
rect -15892 -11192 -15828 -11128
rect -15892 -11272 -15828 -11208
rect -15892 -11352 -15828 -11288
rect -15892 -11432 -15828 -11368
rect -15892 -11512 -15828 -11448
rect -15892 -11592 -15828 -11528
rect -15892 -11672 -15828 -11608
rect -15892 -11752 -15828 -11688
rect -15892 -11832 -15828 -11768
rect -15892 -11912 -15828 -11848
rect -15892 -11992 -15828 -11928
rect -15892 -12072 -15828 -12008
rect -15892 -12152 -15828 -12088
rect -15892 -12232 -15828 -12168
rect -15892 -12312 -15828 -12248
rect -15892 -12392 -15828 -12328
rect -15892 -12472 -15828 -12408
rect -15892 -12552 -15828 -12488
rect -15892 -12632 -15828 -12568
rect -15892 -12712 -15828 -12648
rect -15892 -12792 -15828 -12728
rect -15892 -12872 -15828 -12808
rect -15892 -12952 -15828 -12888
rect -15892 -13032 -15828 -12968
rect -15892 -13112 -15828 -13048
rect -15892 -13192 -15828 -13128
rect -15892 -13272 -15828 -13208
rect -15892 -13352 -15828 -13288
rect -15892 -13432 -15828 -13368
rect -15892 -13512 -15828 -13448
rect -15892 -13592 -15828 -13528
rect -15892 -13672 -15828 -13608
rect -15892 -13752 -15828 -13688
rect -15892 -13832 -15828 -13768
rect -15892 -13912 -15828 -13848
rect -15892 -13992 -15828 -13928
rect -15892 -14072 -15828 -14008
rect -15892 -14152 -15828 -14088
rect -15892 -14232 -15828 -14168
rect -15892 -14312 -15828 -14248
rect -15892 -14392 -15828 -14328
rect -15892 -14472 -15828 -14408
rect -15892 -14552 -15828 -14488
rect -15892 -14632 -15828 -14568
rect -15892 -14712 -15828 -14648
rect -15892 -14792 -15828 -14728
rect -15892 -14872 -15828 -14808
rect -15892 -14952 -15828 -14888
rect -15892 -15032 -15828 -14968
rect -15892 -15112 -15828 -15048
rect -15892 -15192 -15828 -15128
rect -15892 -15272 -15828 -15208
rect -15892 -15352 -15828 -15288
rect -15892 -15432 -15828 -15368
rect -15892 -15512 -15828 -15448
rect -15892 -15592 -15828 -15528
rect -15892 -15672 -15828 -15608
rect -9573 -9592 -9509 -9528
rect -9573 -9672 -9509 -9608
rect -9573 -9752 -9509 -9688
rect -9573 -9832 -9509 -9768
rect -9573 -9912 -9509 -9848
rect -9573 -9992 -9509 -9928
rect -9573 -10072 -9509 -10008
rect -9573 -10152 -9509 -10088
rect -9573 -10232 -9509 -10168
rect -9573 -10312 -9509 -10248
rect -9573 -10392 -9509 -10328
rect -9573 -10472 -9509 -10408
rect -9573 -10552 -9509 -10488
rect -9573 -10632 -9509 -10568
rect -9573 -10712 -9509 -10648
rect -9573 -10792 -9509 -10728
rect -9573 -10872 -9509 -10808
rect -9573 -10952 -9509 -10888
rect -9573 -11032 -9509 -10968
rect -9573 -11112 -9509 -11048
rect -9573 -11192 -9509 -11128
rect -9573 -11272 -9509 -11208
rect -9573 -11352 -9509 -11288
rect -9573 -11432 -9509 -11368
rect -9573 -11512 -9509 -11448
rect -9573 -11592 -9509 -11528
rect -9573 -11672 -9509 -11608
rect -9573 -11752 -9509 -11688
rect -9573 -11832 -9509 -11768
rect -9573 -11912 -9509 -11848
rect -9573 -11992 -9509 -11928
rect -9573 -12072 -9509 -12008
rect -9573 -12152 -9509 -12088
rect -9573 -12232 -9509 -12168
rect -9573 -12312 -9509 -12248
rect -9573 -12392 -9509 -12328
rect -9573 -12472 -9509 -12408
rect -9573 -12552 -9509 -12488
rect -9573 -12632 -9509 -12568
rect -9573 -12712 -9509 -12648
rect -9573 -12792 -9509 -12728
rect -9573 -12872 -9509 -12808
rect -9573 -12952 -9509 -12888
rect -9573 -13032 -9509 -12968
rect -9573 -13112 -9509 -13048
rect -9573 -13192 -9509 -13128
rect -9573 -13272 -9509 -13208
rect -9573 -13352 -9509 -13288
rect -9573 -13432 -9509 -13368
rect -9573 -13512 -9509 -13448
rect -9573 -13592 -9509 -13528
rect -9573 -13672 -9509 -13608
rect -9573 -13752 -9509 -13688
rect -9573 -13832 -9509 -13768
rect -9573 -13912 -9509 -13848
rect -9573 -13992 -9509 -13928
rect -9573 -14072 -9509 -14008
rect -9573 -14152 -9509 -14088
rect -9573 -14232 -9509 -14168
rect -9573 -14312 -9509 -14248
rect -9573 -14392 -9509 -14328
rect -9573 -14472 -9509 -14408
rect -9573 -14552 -9509 -14488
rect -9573 -14632 -9509 -14568
rect -9573 -14712 -9509 -14648
rect -9573 -14792 -9509 -14728
rect -9573 -14872 -9509 -14808
rect -9573 -14952 -9509 -14888
rect -9573 -15032 -9509 -14968
rect -9573 -15112 -9509 -15048
rect -9573 -15192 -9509 -15128
rect -9573 -15272 -9509 -15208
rect -9573 -15352 -9509 -15288
rect -9573 -15432 -9509 -15368
rect -9573 -15512 -9509 -15448
rect -9573 -15592 -9509 -15528
rect -9573 -15672 -9509 -15608
rect -3254 -9592 -3190 -9528
rect -3254 -9672 -3190 -9608
rect -3254 -9752 -3190 -9688
rect -3254 -9832 -3190 -9768
rect -3254 -9912 -3190 -9848
rect -3254 -9992 -3190 -9928
rect -3254 -10072 -3190 -10008
rect -3254 -10152 -3190 -10088
rect -3254 -10232 -3190 -10168
rect -3254 -10312 -3190 -10248
rect -3254 -10392 -3190 -10328
rect -3254 -10472 -3190 -10408
rect -3254 -10552 -3190 -10488
rect -3254 -10632 -3190 -10568
rect -3254 -10712 -3190 -10648
rect -3254 -10792 -3190 -10728
rect -3254 -10872 -3190 -10808
rect -3254 -10952 -3190 -10888
rect -3254 -11032 -3190 -10968
rect -3254 -11112 -3190 -11048
rect -3254 -11192 -3190 -11128
rect -3254 -11272 -3190 -11208
rect -3254 -11352 -3190 -11288
rect -3254 -11432 -3190 -11368
rect -3254 -11512 -3190 -11448
rect -3254 -11592 -3190 -11528
rect -3254 -11672 -3190 -11608
rect -3254 -11752 -3190 -11688
rect -3254 -11832 -3190 -11768
rect -3254 -11912 -3190 -11848
rect -3254 -11992 -3190 -11928
rect -3254 -12072 -3190 -12008
rect -3254 -12152 -3190 -12088
rect -3254 -12232 -3190 -12168
rect -3254 -12312 -3190 -12248
rect -3254 -12392 -3190 -12328
rect -3254 -12472 -3190 -12408
rect -3254 -12552 -3190 -12488
rect -3254 -12632 -3190 -12568
rect -3254 -12712 -3190 -12648
rect -3254 -12792 -3190 -12728
rect -3254 -12872 -3190 -12808
rect -3254 -12952 -3190 -12888
rect -3254 -13032 -3190 -12968
rect -3254 -13112 -3190 -13048
rect -3254 -13192 -3190 -13128
rect -3254 -13272 -3190 -13208
rect -3254 -13352 -3190 -13288
rect -3254 -13432 -3190 -13368
rect -3254 -13512 -3190 -13448
rect -3254 -13592 -3190 -13528
rect -3254 -13672 -3190 -13608
rect -3254 -13752 -3190 -13688
rect -3254 -13832 -3190 -13768
rect -3254 -13912 -3190 -13848
rect -3254 -13992 -3190 -13928
rect -3254 -14072 -3190 -14008
rect -3254 -14152 -3190 -14088
rect -3254 -14232 -3190 -14168
rect -3254 -14312 -3190 -14248
rect -3254 -14392 -3190 -14328
rect -3254 -14472 -3190 -14408
rect -3254 -14552 -3190 -14488
rect -3254 -14632 -3190 -14568
rect -3254 -14712 -3190 -14648
rect -3254 -14792 -3190 -14728
rect -3254 -14872 -3190 -14808
rect -3254 -14952 -3190 -14888
rect -3254 -15032 -3190 -14968
rect -3254 -15112 -3190 -15048
rect -3254 -15192 -3190 -15128
rect -3254 -15272 -3190 -15208
rect -3254 -15352 -3190 -15288
rect -3254 -15432 -3190 -15368
rect -3254 -15512 -3190 -15448
rect -3254 -15592 -3190 -15528
rect -3254 -15672 -3190 -15608
rect 3065 -9592 3129 -9528
rect 3065 -9672 3129 -9608
rect 3065 -9752 3129 -9688
rect 3065 -9832 3129 -9768
rect 3065 -9912 3129 -9848
rect 3065 -9992 3129 -9928
rect 3065 -10072 3129 -10008
rect 3065 -10152 3129 -10088
rect 3065 -10232 3129 -10168
rect 3065 -10312 3129 -10248
rect 3065 -10392 3129 -10328
rect 3065 -10472 3129 -10408
rect 3065 -10552 3129 -10488
rect 3065 -10632 3129 -10568
rect 3065 -10712 3129 -10648
rect 3065 -10792 3129 -10728
rect 3065 -10872 3129 -10808
rect 3065 -10952 3129 -10888
rect 3065 -11032 3129 -10968
rect 3065 -11112 3129 -11048
rect 3065 -11192 3129 -11128
rect 3065 -11272 3129 -11208
rect 3065 -11352 3129 -11288
rect 3065 -11432 3129 -11368
rect 3065 -11512 3129 -11448
rect 3065 -11592 3129 -11528
rect 3065 -11672 3129 -11608
rect 3065 -11752 3129 -11688
rect 3065 -11832 3129 -11768
rect 3065 -11912 3129 -11848
rect 3065 -11992 3129 -11928
rect 3065 -12072 3129 -12008
rect 3065 -12152 3129 -12088
rect 3065 -12232 3129 -12168
rect 3065 -12312 3129 -12248
rect 3065 -12392 3129 -12328
rect 3065 -12472 3129 -12408
rect 3065 -12552 3129 -12488
rect 3065 -12632 3129 -12568
rect 3065 -12712 3129 -12648
rect 3065 -12792 3129 -12728
rect 3065 -12872 3129 -12808
rect 3065 -12952 3129 -12888
rect 3065 -13032 3129 -12968
rect 3065 -13112 3129 -13048
rect 3065 -13192 3129 -13128
rect 3065 -13272 3129 -13208
rect 3065 -13352 3129 -13288
rect 3065 -13432 3129 -13368
rect 3065 -13512 3129 -13448
rect 3065 -13592 3129 -13528
rect 3065 -13672 3129 -13608
rect 3065 -13752 3129 -13688
rect 3065 -13832 3129 -13768
rect 3065 -13912 3129 -13848
rect 3065 -13992 3129 -13928
rect 3065 -14072 3129 -14008
rect 3065 -14152 3129 -14088
rect 3065 -14232 3129 -14168
rect 3065 -14312 3129 -14248
rect 3065 -14392 3129 -14328
rect 3065 -14472 3129 -14408
rect 3065 -14552 3129 -14488
rect 3065 -14632 3129 -14568
rect 3065 -14712 3129 -14648
rect 3065 -14792 3129 -14728
rect 3065 -14872 3129 -14808
rect 3065 -14952 3129 -14888
rect 3065 -15032 3129 -14968
rect 3065 -15112 3129 -15048
rect 3065 -15192 3129 -15128
rect 3065 -15272 3129 -15208
rect 3065 -15352 3129 -15288
rect 3065 -15432 3129 -15368
rect 3065 -15512 3129 -15448
rect 3065 -15592 3129 -15528
rect 3065 -15672 3129 -15608
rect 9384 -9592 9448 -9528
rect 9384 -9672 9448 -9608
rect 9384 -9752 9448 -9688
rect 9384 -9832 9448 -9768
rect 9384 -9912 9448 -9848
rect 9384 -9992 9448 -9928
rect 9384 -10072 9448 -10008
rect 9384 -10152 9448 -10088
rect 9384 -10232 9448 -10168
rect 9384 -10312 9448 -10248
rect 9384 -10392 9448 -10328
rect 9384 -10472 9448 -10408
rect 9384 -10552 9448 -10488
rect 9384 -10632 9448 -10568
rect 9384 -10712 9448 -10648
rect 9384 -10792 9448 -10728
rect 9384 -10872 9448 -10808
rect 9384 -10952 9448 -10888
rect 9384 -11032 9448 -10968
rect 9384 -11112 9448 -11048
rect 9384 -11192 9448 -11128
rect 9384 -11272 9448 -11208
rect 9384 -11352 9448 -11288
rect 9384 -11432 9448 -11368
rect 9384 -11512 9448 -11448
rect 9384 -11592 9448 -11528
rect 9384 -11672 9448 -11608
rect 9384 -11752 9448 -11688
rect 9384 -11832 9448 -11768
rect 9384 -11912 9448 -11848
rect 9384 -11992 9448 -11928
rect 9384 -12072 9448 -12008
rect 9384 -12152 9448 -12088
rect 9384 -12232 9448 -12168
rect 9384 -12312 9448 -12248
rect 9384 -12392 9448 -12328
rect 9384 -12472 9448 -12408
rect 9384 -12552 9448 -12488
rect 9384 -12632 9448 -12568
rect 9384 -12712 9448 -12648
rect 9384 -12792 9448 -12728
rect 9384 -12872 9448 -12808
rect 9384 -12952 9448 -12888
rect 9384 -13032 9448 -12968
rect 9384 -13112 9448 -13048
rect 9384 -13192 9448 -13128
rect 9384 -13272 9448 -13208
rect 9384 -13352 9448 -13288
rect 9384 -13432 9448 -13368
rect 9384 -13512 9448 -13448
rect 9384 -13592 9448 -13528
rect 9384 -13672 9448 -13608
rect 9384 -13752 9448 -13688
rect 9384 -13832 9448 -13768
rect 9384 -13912 9448 -13848
rect 9384 -13992 9448 -13928
rect 9384 -14072 9448 -14008
rect 9384 -14152 9448 -14088
rect 9384 -14232 9448 -14168
rect 9384 -14312 9448 -14248
rect 9384 -14392 9448 -14328
rect 9384 -14472 9448 -14408
rect 9384 -14552 9448 -14488
rect 9384 -14632 9448 -14568
rect 9384 -14712 9448 -14648
rect 9384 -14792 9448 -14728
rect 9384 -14872 9448 -14808
rect 9384 -14952 9448 -14888
rect 9384 -15032 9448 -14968
rect 9384 -15112 9448 -15048
rect 9384 -15192 9448 -15128
rect 9384 -15272 9448 -15208
rect 9384 -15352 9448 -15288
rect 9384 -15432 9448 -15368
rect 9384 -15512 9448 -15448
rect 9384 -15592 9448 -15528
rect 9384 -15672 9448 -15608
rect 15703 -9592 15767 -9528
rect 15703 -9672 15767 -9608
rect 15703 -9752 15767 -9688
rect 15703 -9832 15767 -9768
rect 15703 -9912 15767 -9848
rect 15703 -9992 15767 -9928
rect 15703 -10072 15767 -10008
rect 15703 -10152 15767 -10088
rect 15703 -10232 15767 -10168
rect 15703 -10312 15767 -10248
rect 15703 -10392 15767 -10328
rect 15703 -10472 15767 -10408
rect 15703 -10552 15767 -10488
rect 15703 -10632 15767 -10568
rect 15703 -10712 15767 -10648
rect 15703 -10792 15767 -10728
rect 15703 -10872 15767 -10808
rect 15703 -10952 15767 -10888
rect 15703 -11032 15767 -10968
rect 15703 -11112 15767 -11048
rect 15703 -11192 15767 -11128
rect 15703 -11272 15767 -11208
rect 15703 -11352 15767 -11288
rect 15703 -11432 15767 -11368
rect 15703 -11512 15767 -11448
rect 15703 -11592 15767 -11528
rect 15703 -11672 15767 -11608
rect 15703 -11752 15767 -11688
rect 15703 -11832 15767 -11768
rect 15703 -11912 15767 -11848
rect 15703 -11992 15767 -11928
rect 15703 -12072 15767 -12008
rect 15703 -12152 15767 -12088
rect 15703 -12232 15767 -12168
rect 15703 -12312 15767 -12248
rect 15703 -12392 15767 -12328
rect 15703 -12472 15767 -12408
rect 15703 -12552 15767 -12488
rect 15703 -12632 15767 -12568
rect 15703 -12712 15767 -12648
rect 15703 -12792 15767 -12728
rect 15703 -12872 15767 -12808
rect 15703 -12952 15767 -12888
rect 15703 -13032 15767 -12968
rect 15703 -13112 15767 -13048
rect 15703 -13192 15767 -13128
rect 15703 -13272 15767 -13208
rect 15703 -13352 15767 -13288
rect 15703 -13432 15767 -13368
rect 15703 -13512 15767 -13448
rect 15703 -13592 15767 -13528
rect 15703 -13672 15767 -13608
rect 15703 -13752 15767 -13688
rect 15703 -13832 15767 -13768
rect 15703 -13912 15767 -13848
rect 15703 -13992 15767 -13928
rect 15703 -14072 15767 -14008
rect 15703 -14152 15767 -14088
rect 15703 -14232 15767 -14168
rect 15703 -14312 15767 -14248
rect 15703 -14392 15767 -14328
rect 15703 -14472 15767 -14408
rect 15703 -14552 15767 -14488
rect 15703 -14632 15767 -14568
rect 15703 -14712 15767 -14648
rect 15703 -14792 15767 -14728
rect 15703 -14872 15767 -14808
rect 15703 -14952 15767 -14888
rect 15703 -15032 15767 -14968
rect 15703 -15112 15767 -15048
rect 15703 -15192 15767 -15128
rect 15703 -15272 15767 -15208
rect 15703 -15352 15767 -15288
rect 15703 -15432 15767 -15368
rect 15703 -15512 15767 -15448
rect 15703 -15592 15767 -15528
rect 15703 -15672 15767 -15608
rect 22022 -9592 22086 -9528
rect 22022 -9672 22086 -9608
rect 22022 -9752 22086 -9688
rect 22022 -9832 22086 -9768
rect 22022 -9912 22086 -9848
rect 22022 -9992 22086 -9928
rect 22022 -10072 22086 -10008
rect 22022 -10152 22086 -10088
rect 22022 -10232 22086 -10168
rect 22022 -10312 22086 -10248
rect 22022 -10392 22086 -10328
rect 22022 -10472 22086 -10408
rect 22022 -10552 22086 -10488
rect 22022 -10632 22086 -10568
rect 22022 -10712 22086 -10648
rect 22022 -10792 22086 -10728
rect 22022 -10872 22086 -10808
rect 22022 -10952 22086 -10888
rect 22022 -11032 22086 -10968
rect 22022 -11112 22086 -11048
rect 22022 -11192 22086 -11128
rect 22022 -11272 22086 -11208
rect 22022 -11352 22086 -11288
rect 22022 -11432 22086 -11368
rect 22022 -11512 22086 -11448
rect 22022 -11592 22086 -11528
rect 22022 -11672 22086 -11608
rect 22022 -11752 22086 -11688
rect 22022 -11832 22086 -11768
rect 22022 -11912 22086 -11848
rect 22022 -11992 22086 -11928
rect 22022 -12072 22086 -12008
rect 22022 -12152 22086 -12088
rect 22022 -12232 22086 -12168
rect 22022 -12312 22086 -12248
rect 22022 -12392 22086 -12328
rect 22022 -12472 22086 -12408
rect 22022 -12552 22086 -12488
rect 22022 -12632 22086 -12568
rect 22022 -12712 22086 -12648
rect 22022 -12792 22086 -12728
rect 22022 -12872 22086 -12808
rect 22022 -12952 22086 -12888
rect 22022 -13032 22086 -12968
rect 22022 -13112 22086 -13048
rect 22022 -13192 22086 -13128
rect 22022 -13272 22086 -13208
rect 22022 -13352 22086 -13288
rect 22022 -13432 22086 -13368
rect 22022 -13512 22086 -13448
rect 22022 -13592 22086 -13528
rect 22022 -13672 22086 -13608
rect 22022 -13752 22086 -13688
rect 22022 -13832 22086 -13768
rect 22022 -13912 22086 -13848
rect 22022 -13992 22086 -13928
rect 22022 -14072 22086 -14008
rect 22022 -14152 22086 -14088
rect 22022 -14232 22086 -14168
rect 22022 -14312 22086 -14248
rect 22022 -14392 22086 -14328
rect 22022 -14472 22086 -14408
rect 22022 -14552 22086 -14488
rect 22022 -14632 22086 -14568
rect 22022 -14712 22086 -14648
rect 22022 -14792 22086 -14728
rect 22022 -14872 22086 -14808
rect 22022 -14952 22086 -14888
rect 22022 -15032 22086 -14968
rect 22022 -15112 22086 -15048
rect 22022 -15192 22086 -15128
rect 22022 -15272 22086 -15208
rect 22022 -15352 22086 -15288
rect 22022 -15432 22086 -15368
rect 22022 -15512 22086 -15448
rect 22022 -15592 22086 -15528
rect 22022 -15672 22086 -15608
rect 28341 -9592 28405 -9528
rect 28341 -9672 28405 -9608
rect 28341 -9752 28405 -9688
rect 28341 -9832 28405 -9768
rect 28341 -9912 28405 -9848
rect 28341 -9992 28405 -9928
rect 28341 -10072 28405 -10008
rect 28341 -10152 28405 -10088
rect 28341 -10232 28405 -10168
rect 28341 -10312 28405 -10248
rect 28341 -10392 28405 -10328
rect 28341 -10472 28405 -10408
rect 28341 -10552 28405 -10488
rect 28341 -10632 28405 -10568
rect 28341 -10712 28405 -10648
rect 28341 -10792 28405 -10728
rect 28341 -10872 28405 -10808
rect 28341 -10952 28405 -10888
rect 28341 -11032 28405 -10968
rect 28341 -11112 28405 -11048
rect 28341 -11192 28405 -11128
rect 28341 -11272 28405 -11208
rect 28341 -11352 28405 -11288
rect 28341 -11432 28405 -11368
rect 28341 -11512 28405 -11448
rect 28341 -11592 28405 -11528
rect 28341 -11672 28405 -11608
rect 28341 -11752 28405 -11688
rect 28341 -11832 28405 -11768
rect 28341 -11912 28405 -11848
rect 28341 -11992 28405 -11928
rect 28341 -12072 28405 -12008
rect 28341 -12152 28405 -12088
rect 28341 -12232 28405 -12168
rect 28341 -12312 28405 -12248
rect 28341 -12392 28405 -12328
rect 28341 -12472 28405 -12408
rect 28341 -12552 28405 -12488
rect 28341 -12632 28405 -12568
rect 28341 -12712 28405 -12648
rect 28341 -12792 28405 -12728
rect 28341 -12872 28405 -12808
rect 28341 -12952 28405 -12888
rect 28341 -13032 28405 -12968
rect 28341 -13112 28405 -13048
rect 28341 -13192 28405 -13128
rect 28341 -13272 28405 -13208
rect 28341 -13352 28405 -13288
rect 28341 -13432 28405 -13368
rect 28341 -13512 28405 -13448
rect 28341 -13592 28405 -13528
rect 28341 -13672 28405 -13608
rect 28341 -13752 28405 -13688
rect 28341 -13832 28405 -13768
rect 28341 -13912 28405 -13848
rect 28341 -13992 28405 -13928
rect 28341 -14072 28405 -14008
rect 28341 -14152 28405 -14088
rect 28341 -14232 28405 -14168
rect 28341 -14312 28405 -14248
rect 28341 -14392 28405 -14328
rect 28341 -14472 28405 -14408
rect 28341 -14552 28405 -14488
rect 28341 -14632 28405 -14568
rect 28341 -14712 28405 -14648
rect 28341 -14792 28405 -14728
rect 28341 -14872 28405 -14808
rect 28341 -14952 28405 -14888
rect 28341 -15032 28405 -14968
rect 28341 -15112 28405 -15048
rect 28341 -15192 28405 -15128
rect 28341 -15272 28405 -15208
rect 28341 -15352 28405 -15288
rect 28341 -15432 28405 -15368
rect 28341 -15512 28405 -15448
rect 28341 -15592 28405 -15528
rect 28341 -15672 28405 -15608
rect 34660 -9592 34724 -9528
rect 34660 -9672 34724 -9608
rect 34660 -9752 34724 -9688
rect 34660 -9832 34724 -9768
rect 34660 -9912 34724 -9848
rect 34660 -9992 34724 -9928
rect 34660 -10072 34724 -10008
rect 34660 -10152 34724 -10088
rect 34660 -10232 34724 -10168
rect 34660 -10312 34724 -10248
rect 34660 -10392 34724 -10328
rect 34660 -10472 34724 -10408
rect 34660 -10552 34724 -10488
rect 34660 -10632 34724 -10568
rect 34660 -10712 34724 -10648
rect 34660 -10792 34724 -10728
rect 34660 -10872 34724 -10808
rect 34660 -10952 34724 -10888
rect 34660 -11032 34724 -10968
rect 34660 -11112 34724 -11048
rect 34660 -11192 34724 -11128
rect 34660 -11272 34724 -11208
rect 34660 -11352 34724 -11288
rect 34660 -11432 34724 -11368
rect 34660 -11512 34724 -11448
rect 34660 -11592 34724 -11528
rect 34660 -11672 34724 -11608
rect 34660 -11752 34724 -11688
rect 34660 -11832 34724 -11768
rect 34660 -11912 34724 -11848
rect 34660 -11992 34724 -11928
rect 34660 -12072 34724 -12008
rect 34660 -12152 34724 -12088
rect 34660 -12232 34724 -12168
rect 34660 -12312 34724 -12248
rect 34660 -12392 34724 -12328
rect 34660 -12472 34724 -12408
rect 34660 -12552 34724 -12488
rect 34660 -12632 34724 -12568
rect 34660 -12712 34724 -12648
rect 34660 -12792 34724 -12728
rect 34660 -12872 34724 -12808
rect 34660 -12952 34724 -12888
rect 34660 -13032 34724 -12968
rect 34660 -13112 34724 -13048
rect 34660 -13192 34724 -13128
rect 34660 -13272 34724 -13208
rect 34660 -13352 34724 -13288
rect 34660 -13432 34724 -13368
rect 34660 -13512 34724 -13448
rect 34660 -13592 34724 -13528
rect 34660 -13672 34724 -13608
rect 34660 -13752 34724 -13688
rect 34660 -13832 34724 -13768
rect 34660 -13912 34724 -13848
rect 34660 -13992 34724 -13928
rect 34660 -14072 34724 -14008
rect 34660 -14152 34724 -14088
rect 34660 -14232 34724 -14168
rect 34660 -14312 34724 -14248
rect 34660 -14392 34724 -14328
rect 34660 -14472 34724 -14408
rect 34660 -14552 34724 -14488
rect 34660 -14632 34724 -14568
rect 34660 -14712 34724 -14648
rect 34660 -14792 34724 -14728
rect 34660 -14872 34724 -14808
rect 34660 -14952 34724 -14888
rect 34660 -15032 34724 -14968
rect 34660 -15112 34724 -15048
rect 34660 -15192 34724 -15128
rect 34660 -15272 34724 -15208
rect 34660 -15352 34724 -15288
rect 34660 -15432 34724 -15368
rect 34660 -15512 34724 -15448
rect 34660 -15592 34724 -15528
rect 34660 -15672 34724 -15608
rect 40979 -9592 41043 -9528
rect 40979 -9672 41043 -9608
rect 40979 -9752 41043 -9688
rect 40979 -9832 41043 -9768
rect 40979 -9912 41043 -9848
rect 40979 -9992 41043 -9928
rect 40979 -10072 41043 -10008
rect 40979 -10152 41043 -10088
rect 40979 -10232 41043 -10168
rect 40979 -10312 41043 -10248
rect 40979 -10392 41043 -10328
rect 40979 -10472 41043 -10408
rect 40979 -10552 41043 -10488
rect 40979 -10632 41043 -10568
rect 40979 -10712 41043 -10648
rect 40979 -10792 41043 -10728
rect 40979 -10872 41043 -10808
rect 40979 -10952 41043 -10888
rect 40979 -11032 41043 -10968
rect 40979 -11112 41043 -11048
rect 40979 -11192 41043 -11128
rect 40979 -11272 41043 -11208
rect 40979 -11352 41043 -11288
rect 40979 -11432 41043 -11368
rect 40979 -11512 41043 -11448
rect 40979 -11592 41043 -11528
rect 40979 -11672 41043 -11608
rect 40979 -11752 41043 -11688
rect 40979 -11832 41043 -11768
rect 40979 -11912 41043 -11848
rect 40979 -11992 41043 -11928
rect 40979 -12072 41043 -12008
rect 40979 -12152 41043 -12088
rect 40979 -12232 41043 -12168
rect 40979 -12312 41043 -12248
rect 40979 -12392 41043 -12328
rect 40979 -12472 41043 -12408
rect 40979 -12552 41043 -12488
rect 40979 -12632 41043 -12568
rect 40979 -12712 41043 -12648
rect 40979 -12792 41043 -12728
rect 40979 -12872 41043 -12808
rect 40979 -12952 41043 -12888
rect 40979 -13032 41043 -12968
rect 40979 -13112 41043 -13048
rect 40979 -13192 41043 -13128
rect 40979 -13272 41043 -13208
rect 40979 -13352 41043 -13288
rect 40979 -13432 41043 -13368
rect 40979 -13512 41043 -13448
rect 40979 -13592 41043 -13528
rect 40979 -13672 41043 -13608
rect 40979 -13752 41043 -13688
rect 40979 -13832 41043 -13768
rect 40979 -13912 41043 -13848
rect 40979 -13992 41043 -13928
rect 40979 -14072 41043 -14008
rect 40979 -14152 41043 -14088
rect 40979 -14232 41043 -14168
rect 40979 -14312 41043 -14248
rect 40979 -14392 41043 -14328
rect 40979 -14472 41043 -14408
rect 40979 -14552 41043 -14488
rect 40979 -14632 41043 -14568
rect 40979 -14712 41043 -14648
rect 40979 -14792 41043 -14728
rect 40979 -14872 41043 -14808
rect 40979 -14952 41043 -14888
rect 40979 -15032 41043 -14968
rect 40979 -15112 41043 -15048
rect 40979 -15192 41043 -15128
rect 40979 -15272 41043 -15208
rect 40979 -15352 41043 -15288
rect 40979 -15432 41043 -15368
rect 40979 -15512 41043 -15448
rect 40979 -15592 41043 -15528
rect 40979 -15672 41043 -15608
rect 47298 -9592 47362 -9528
rect 47298 -9672 47362 -9608
rect 47298 -9752 47362 -9688
rect 47298 -9832 47362 -9768
rect 47298 -9912 47362 -9848
rect 47298 -9992 47362 -9928
rect 47298 -10072 47362 -10008
rect 47298 -10152 47362 -10088
rect 47298 -10232 47362 -10168
rect 47298 -10312 47362 -10248
rect 47298 -10392 47362 -10328
rect 47298 -10472 47362 -10408
rect 47298 -10552 47362 -10488
rect 47298 -10632 47362 -10568
rect 47298 -10712 47362 -10648
rect 47298 -10792 47362 -10728
rect 47298 -10872 47362 -10808
rect 47298 -10952 47362 -10888
rect 47298 -11032 47362 -10968
rect 47298 -11112 47362 -11048
rect 47298 -11192 47362 -11128
rect 47298 -11272 47362 -11208
rect 47298 -11352 47362 -11288
rect 47298 -11432 47362 -11368
rect 47298 -11512 47362 -11448
rect 47298 -11592 47362 -11528
rect 47298 -11672 47362 -11608
rect 47298 -11752 47362 -11688
rect 47298 -11832 47362 -11768
rect 47298 -11912 47362 -11848
rect 47298 -11992 47362 -11928
rect 47298 -12072 47362 -12008
rect 47298 -12152 47362 -12088
rect 47298 -12232 47362 -12168
rect 47298 -12312 47362 -12248
rect 47298 -12392 47362 -12328
rect 47298 -12472 47362 -12408
rect 47298 -12552 47362 -12488
rect 47298 -12632 47362 -12568
rect 47298 -12712 47362 -12648
rect 47298 -12792 47362 -12728
rect 47298 -12872 47362 -12808
rect 47298 -12952 47362 -12888
rect 47298 -13032 47362 -12968
rect 47298 -13112 47362 -13048
rect 47298 -13192 47362 -13128
rect 47298 -13272 47362 -13208
rect 47298 -13352 47362 -13288
rect 47298 -13432 47362 -13368
rect 47298 -13512 47362 -13448
rect 47298 -13592 47362 -13528
rect 47298 -13672 47362 -13608
rect 47298 -13752 47362 -13688
rect 47298 -13832 47362 -13768
rect 47298 -13912 47362 -13848
rect 47298 -13992 47362 -13928
rect 47298 -14072 47362 -14008
rect 47298 -14152 47362 -14088
rect 47298 -14232 47362 -14168
rect 47298 -14312 47362 -14248
rect 47298 -14392 47362 -14328
rect 47298 -14472 47362 -14408
rect 47298 -14552 47362 -14488
rect 47298 -14632 47362 -14568
rect 47298 -14712 47362 -14648
rect 47298 -14792 47362 -14728
rect 47298 -14872 47362 -14808
rect 47298 -14952 47362 -14888
rect 47298 -15032 47362 -14968
rect 47298 -15112 47362 -15048
rect 47298 -15192 47362 -15128
rect 47298 -15272 47362 -15208
rect 47298 -15352 47362 -15288
rect 47298 -15432 47362 -15368
rect 47298 -15512 47362 -15448
rect 47298 -15592 47362 -15528
rect 47298 -15672 47362 -15608
rect -41168 -15892 -41104 -15828
rect -41168 -15972 -41104 -15908
rect -41168 -16052 -41104 -15988
rect -41168 -16132 -41104 -16068
rect -41168 -16212 -41104 -16148
rect -41168 -16292 -41104 -16228
rect -41168 -16372 -41104 -16308
rect -41168 -16452 -41104 -16388
rect -41168 -16532 -41104 -16468
rect -41168 -16612 -41104 -16548
rect -41168 -16692 -41104 -16628
rect -41168 -16772 -41104 -16708
rect -41168 -16852 -41104 -16788
rect -41168 -16932 -41104 -16868
rect -41168 -17012 -41104 -16948
rect -41168 -17092 -41104 -17028
rect -41168 -17172 -41104 -17108
rect -41168 -17252 -41104 -17188
rect -41168 -17332 -41104 -17268
rect -41168 -17412 -41104 -17348
rect -41168 -17492 -41104 -17428
rect -41168 -17572 -41104 -17508
rect -41168 -17652 -41104 -17588
rect -41168 -17732 -41104 -17668
rect -41168 -17812 -41104 -17748
rect -41168 -17892 -41104 -17828
rect -41168 -17972 -41104 -17908
rect -41168 -18052 -41104 -17988
rect -41168 -18132 -41104 -18068
rect -41168 -18212 -41104 -18148
rect -41168 -18292 -41104 -18228
rect -41168 -18372 -41104 -18308
rect -41168 -18452 -41104 -18388
rect -41168 -18532 -41104 -18468
rect -41168 -18612 -41104 -18548
rect -41168 -18692 -41104 -18628
rect -41168 -18772 -41104 -18708
rect -41168 -18852 -41104 -18788
rect -41168 -18932 -41104 -18868
rect -41168 -19012 -41104 -18948
rect -41168 -19092 -41104 -19028
rect -41168 -19172 -41104 -19108
rect -41168 -19252 -41104 -19188
rect -41168 -19332 -41104 -19268
rect -41168 -19412 -41104 -19348
rect -41168 -19492 -41104 -19428
rect -41168 -19572 -41104 -19508
rect -41168 -19652 -41104 -19588
rect -41168 -19732 -41104 -19668
rect -41168 -19812 -41104 -19748
rect -41168 -19892 -41104 -19828
rect -41168 -19972 -41104 -19908
rect -41168 -20052 -41104 -19988
rect -41168 -20132 -41104 -20068
rect -41168 -20212 -41104 -20148
rect -41168 -20292 -41104 -20228
rect -41168 -20372 -41104 -20308
rect -41168 -20452 -41104 -20388
rect -41168 -20532 -41104 -20468
rect -41168 -20612 -41104 -20548
rect -41168 -20692 -41104 -20628
rect -41168 -20772 -41104 -20708
rect -41168 -20852 -41104 -20788
rect -41168 -20932 -41104 -20868
rect -41168 -21012 -41104 -20948
rect -41168 -21092 -41104 -21028
rect -41168 -21172 -41104 -21108
rect -41168 -21252 -41104 -21188
rect -41168 -21332 -41104 -21268
rect -41168 -21412 -41104 -21348
rect -41168 -21492 -41104 -21428
rect -41168 -21572 -41104 -21508
rect -41168 -21652 -41104 -21588
rect -41168 -21732 -41104 -21668
rect -41168 -21812 -41104 -21748
rect -41168 -21892 -41104 -21828
rect -41168 -21972 -41104 -21908
rect -34849 -15892 -34785 -15828
rect -34849 -15972 -34785 -15908
rect -34849 -16052 -34785 -15988
rect -34849 -16132 -34785 -16068
rect -34849 -16212 -34785 -16148
rect -34849 -16292 -34785 -16228
rect -34849 -16372 -34785 -16308
rect -34849 -16452 -34785 -16388
rect -34849 -16532 -34785 -16468
rect -34849 -16612 -34785 -16548
rect -34849 -16692 -34785 -16628
rect -34849 -16772 -34785 -16708
rect -34849 -16852 -34785 -16788
rect -34849 -16932 -34785 -16868
rect -34849 -17012 -34785 -16948
rect -34849 -17092 -34785 -17028
rect -34849 -17172 -34785 -17108
rect -34849 -17252 -34785 -17188
rect -34849 -17332 -34785 -17268
rect -34849 -17412 -34785 -17348
rect -34849 -17492 -34785 -17428
rect -34849 -17572 -34785 -17508
rect -34849 -17652 -34785 -17588
rect -34849 -17732 -34785 -17668
rect -34849 -17812 -34785 -17748
rect -34849 -17892 -34785 -17828
rect -34849 -17972 -34785 -17908
rect -34849 -18052 -34785 -17988
rect -34849 -18132 -34785 -18068
rect -34849 -18212 -34785 -18148
rect -34849 -18292 -34785 -18228
rect -34849 -18372 -34785 -18308
rect -34849 -18452 -34785 -18388
rect -34849 -18532 -34785 -18468
rect -34849 -18612 -34785 -18548
rect -34849 -18692 -34785 -18628
rect -34849 -18772 -34785 -18708
rect -34849 -18852 -34785 -18788
rect -34849 -18932 -34785 -18868
rect -34849 -19012 -34785 -18948
rect -34849 -19092 -34785 -19028
rect -34849 -19172 -34785 -19108
rect -34849 -19252 -34785 -19188
rect -34849 -19332 -34785 -19268
rect -34849 -19412 -34785 -19348
rect -34849 -19492 -34785 -19428
rect -34849 -19572 -34785 -19508
rect -34849 -19652 -34785 -19588
rect -34849 -19732 -34785 -19668
rect -34849 -19812 -34785 -19748
rect -34849 -19892 -34785 -19828
rect -34849 -19972 -34785 -19908
rect -34849 -20052 -34785 -19988
rect -34849 -20132 -34785 -20068
rect -34849 -20212 -34785 -20148
rect -34849 -20292 -34785 -20228
rect -34849 -20372 -34785 -20308
rect -34849 -20452 -34785 -20388
rect -34849 -20532 -34785 -20468
rect -34849 -20612 -34785 -20548
rect -34849 -20692 -34785 -20628
rect -34849 -20772 -34785 -20708
rect -34849 -20852 -34785 -20788
rect -34849 -20932 -34785 -20868
rect -34849 -21012 -34785 -20948
rect -34849 -21092 -34785 -21028
rect -34849 -21172 -34785 -21108
rect -34849 -21252 -34785 -21188
rect -34849 -21332 -34785 -21268
rect -34849 -21412 -34785 -21348
rect -34849 -21492 -34785 -21428
rect -34849 -21572 -34785 -21508
rect -34849 -21652 -34785 -21588
rect -34849 -21732 -34785 -21668
rect -34849 -21812 -34785 -21748
rect -34849 -21892 -34785 -21828
rect -34849 -21972 -34785 -21908
rect -28530 -15892 -28466 -15828
rect -28530 -15972 -28466 -15908
rect -28530 -16052 -28466 -15988
rect -28530 -16132 -28466 -16068
rect -28530 -16212 -28466 -16148
rect -28530 -16292 -28466 -16228
rect -28530 -16372 -28466 -16308
rect -28530 -16452 -28466 -16388
rect -28530 -16532 -28466 -16468
rect -28530 -16612 -28466 -16548
rect -28530 -16692 -28466 -16628
rect -28530 -16772 -28466 -16708
rect -28530 -16852 -28466 -16788
rect -28530 -16932 -28466 -16868
rect -28530 -17012 -28466 -16948
rect -28530 -17092 -28466 -17028
rect -28530 -17172 -28466 -17108
rect -28530 -17252 -28466 -17188
rect -28530 -17332 -28466 -17268
rect -28530 -17412 -28466 -17348
rect -28530 -17492 -28466 -17428
rect -28530 -17572 -28466 -17508
rect -28530 -17652 -28466 -17588
rect -28530 -17732 -28466 -17668
rect -28530 -17812 -28466 -17748
rect -28530 -17892 -28466 -17828
rect -28530 -17972 -28466 -17908
rect -28530 -18052 -28466 -17988
rect -28530 -18132 -28466 -18068
rect -28530 -18212 -28466 -18148
rect -28530 -18292 -28466 -18228
rect -28530 -18372 -28466 -18308
rect -28530 -18452 -28466 -18388
rect -28530 -18532 -28466 -18468
rect -28530 -18612 -28466 -18548
rect -28530 -18692 -28466 -18628
rect -28530 -18772 -28466 -18708
rect -28530 -18852 -28466 -18788
rect -28530 -18932 -28466 -18868
rect -28530 -19012 -28466 -18948
rect -28530 -19092 -28466 -19028
rect -28530 -19172 -28466 -19108
rect -28530 -19252 -28466 -19188
rect -28530 -19332 -28466 -19268
rect -28530 -19412 -28466 -19348
rect -28530 -19492 -28466 -19428
rect -28530 -19572 -28466 -19508
rect -28530 -19652 -28466 -19588
rect -28530 -19732 -28466 -19668
rect -28530 -19812 -28466 -19748
rect -28530 -19892 -28466 -19828
rect -28530 -19972 -28466 -19908
rect -28530 -20052 -28466 -19988
rect -28530 -20132 -28466 -20068
rect -28530 -20212 -28466 -20148
rect -28530 -20292 -28466 -20228
rect -28530 -20372 -28466 -20308
rect -28530 -20452 -28466 -20388
rect -28530 -20532 -28466 -20468
rect -28530 -20612 -28466 -20548
rect -28530 -20692 -28466 -20628
rect -28530 -20772 -28466 -20708
rect -28530 -20852 -28466 -20788
rect -28530 -20932 -28466 -20868
rect -28530 -21012 -28466 -20948
rect -28530 -21092 -28466 -21028
rect -28530 -21172 -28466 -21108
rect -28530 -21252 -28466 -21188
rect -28530 -21332 -28466 -21268
rect -28530 -21412 -28466 -21348
rect -28530 -21492 -28466 -21428
rect -28530 -21572 -28466 -21508
rect -28530 -21652 -28466 -21588
rect -28530 -21732 -28466 -21668
rect -28530 -21812 -28466 -21748
rect -28530 -21892 -28466 -21828
rect -28530 -21972 -28466 -21908
rect -22211 -15892 -22147 -15828
rect -22211 -15972 -22147 -15908
rect -22211 -16052 -22147 -15988
rect -22211 -16132 -22147 -16068
rect -22211 -16212 -22147 -16148
rect -22211 -16292 -22147 -16228
rect -22211 -16372 -22147 -16308
rect -22211 -16452 -22147 -16388
rect -22211 -16532 -22147 -16468
rect -22211 -16612 -22147 -16548
rect -22211 -16692 -22147 -16628
rect -22211 -16772 -22147 -16708
rect -22211 -16852 -22147 -16788
rect -22211 -16932 -22147 -16868
rect -22211 -17012 -22147 -16948
rect -22211 -17092 -22147 -17028
rect -22211 -17172 -22147 -17108
rect -22211 -17252 -22147 -17188
rect -22211 -17332 -22147 -17268
rect -22211 -17412 -22147 -17348
rect -22211 -17492 -22147 -17428
rect -22211 -17572 -22147 -17508
rect -22211 -17652 -22147 -17588
rect -22211 -17732 -22147 -17668
rect -22211 -17812 -22147 -17748
rect -22211 -17892 -22147 -17828
rect -22211 -17972 -22147 -17908
rect -22211 -18052 -22147 -17988
rect -22211 -18132 -22147 -18068
rect -22211 -18212 -22147 -18148
rect -22211 -18292 -22147 -18228
rect -22211 -18372 -22147 -18308
rect -22211 -18452 -22147 -18388
rect -22211 -18532 -22147 -18468
rect -22211 -18612 -22147 -18548
rect -22211 -18692 -22147 -18628
rect -22211 -18772 -22147 -18708
rect -22211 -18852 -22147 -18788
rect -22211 -18932 -22147 -18868
rect -22211 -19012 -22147 -18948
rect -22211 -19092 -22147 -19028
rect -22211 -19172 -22147 -19108
rect -22211 -19252 -22147 -19188
rect -22211 -19332 -22147 -19268
rect -22211 -19412 -22147 -19348
rect -22211 -19492 -22147 -19428
rect -22211 -19572 -22147 -19508
rect -22211 -19652 -22147 -19588
rect -22211 -19732 -22147 -19668
rect -22211 -19812 -22147 -19748
rect -22211 -19892 -22147 -19828
rect -22211 -19972 -22147 -19908
rect -22211 -20052 -22147 -19988
rect -22211 -20132 -22147 -20068
rect -22211 -20212 -22147 -20148
rect -22211 -20292 -22147 -20228
rect -22211 -20372 -22147 -20308
rect -22211 -20452 -22147 -20388
rect -22211 -20532 -22147 -20468
rect -22211 -20612 -22147 -20548
rect -22211 -20692 -22147 -20628
rect -22211 -20772 -22147 -20708
rect -22211 -20852 -22147 -20788
rect -22211 -20932 -22147 -20868
rect -22211 -21012 -22147 -20948
rect -22211 -21092 -22147 -21028
rect -22211 -21172 -22147 -21108
rect -22211 -21252 -22147 -21188
rect -22211 -21332 -22147 -21268
rect -22211 -21412 -22147 -21348
rect -22211 -21492 -22147 -21428
rect -22211 -21572 -22147 -21508
rect -22211 -21652 -22147 -21588
rect -22211 -21732 -22147 -21668
rect -22211 -21812 -22147 -21748
rect -22211 -21892 -22147 -21828
rect -22211 -21972 -22147 -21908
rect -15892 -15892 -15828 -15828
rect -15892 -15972 -15828 -15908
rect -15892 -16052 -15828 -15988
rect -15892 -16132 -15828 -16068
rect -15892 -16212 -15828 -16148
rect -15892 -16292 -15828 -16228
rect -15892 -16372 -15828 -16308
rect -15892 -16452 -15828 -16388
rect -15892 -16532 -15828 -16468
rect -15892 -16612 -15828 -16548
rect -15892 -16692 -15828 -16628
rect -15892 -16772 -15828 -16708
rect -15892 -16852 -15828 -16788
rect -15892 -16932 -15828 -16868
rect -15892 -17012 -15828 -16948
rect -15892 -17092 -15828 -17028
rect -15892 -17172 -15828 -17108
rect -15892 -17252 -15828 -17188
rect -15892 -17332 -15828 -17268
rect -15892 -17412 -15828 -17348
rect -15892 -17492 -15828 -17428
rect -15892 -17572 -15828 -17508
rect -15892 -17652 -15828 -17588
rect -15892 -17732 -15828 -17668
rect -15892 -17812 -15828 -17748
rect -15892 -17892 -15828 -17828
rect -15892 -17972 -15828 -17908
rect -15892 -18052 -15828 -17988
rect -15892 -18132 -15828 -18068
rect -15892 -18212 -15828 -18148
rect -15892 -18292 -15828 -18228
rect -15892 -18372 -15828 -18308
rect -15892 -18452 -15828 -18388
rect -15892 -18532 -15828 -18468
rect -15892 -18612 -15828 -18548
rect -15892 -18692 -15828 -18628
rect -15892 -18772 -15828 -18708
rect -15892 -18852 -15828 -18788
rect -15892 -18932 -15828 -18868
rect -15892 -19012 -15828 -18948
rect -15892 -19092 -15828 -19028
rect -15892 -19172 -15828 -19108
rect -15892 -19252 -15828 -19188
rect -15892 -19332 -15828 -19268
rect -15892 -19412 -15828 -19348
rect -15892 -19492 -15828 -19428
rect -15892 -19572 -15828 -19508
rect -15892 -19652 -15828 -19588
rect -15892 -19732 -15828 -19668
rect -15892 -19812 -15828 -19748
rect -15892 -19892 -15828 -19828
rect -15892 -19972 -15828 -19908
rect -15892 -20052 -15828 -19988
rect -15892 -20132 -15828 -20068
rect -15892 -20212 -15828 -20148
rect -15892 -20292 -15828 -20228
rect -15892 -20372 -15828 -20308
rect -15892 -20452 -15828 -20388
rect -15892 -20532 -15828 -20468
rect -15892 -20612 -15828 -20548
rect -15892 -20692 -15828 -20628
rect -15892 -20772 -15828 -20708
rect -15892 -20852 -15828 -20788
rect -15892 -20932 -15828 -20868
rect -15892 -21012 -15828 -20948
rect -15892 -21092 -15828 -21028
rect -15892 -21172 -15828 -21108
rect -15892 -21252 -15828 -21188
rect -15892 -21332 -15828 -21268
rect -15892 -21412 -15828 -21348
rect -15892 -21492 -15828 -21428
rect -15892 -21572 -15828 -21508
rect -15892 -21652 -15828 -21588
rect -15892 -21732 -15828 -21668
rect -15892 -21812 -15828 -21748
rect -15892 -21892 -15828 -21828
rect -15892 -21972 -15828 -21908
rect -9573 -15892 -9509 -15828
rect -9573 -15972 -9509 -15908
rect -9573 -16052 -9509 -15988
rect -9573 -16132 -9509 -16068
rect -9573 -16212 -9509 -16148
rect -9573 -16292 -9509 -16228
rect -9573 -16372 -9509 -16308
rect -9573 -16452 -9509 -16388
rect -9573 -16532 -9509 -16468
rect -9573 -16612 -9509 -16548
rect -9573 -16692 -9509 -16628
rect -9573 -16772 -9509 -16708
rect -9573 -16852 -9509 -16788
rect -9573 -16932 -9509 -16868
rect -9573 -17012 -9509 -16948
rect -9573 -17092 -9509 -17028
rect -9573 -17172 -9509 -17108
rect -9573 -17252 -9509 -17188
rect -9573 -17332 -9509 -17268
rect -9573 -17412 -9509 -17348
rect -9573 -17492 -9509 -17428
rect -9573 -17572 -9509 -17508
rect -9573 -17652 -9509 -17588
rect -9573 -17732 -9509 -17668
rect -9573 -17812 -9509 -17748
rect -9573 -17892 -9509 -17828
rect -9573 -17972 -9509 -17908
rect -9573 -18052 -9509 -17988
rect -9573 -18132 -9509 -18068
rect -9573 -18212 -9509 -18148
rect -9573 -18292 -9509 -18228
rect -9573 -18372 -9509 -18308
rect -9573 -18452 -9509 -18388
rect -9573 -18532 -9509 -18468
rect -9573 -18612 -9509 -18548
rect -9573 -18692 -9509 -18628
rect -9573 -18772 -9509 -18708
rect -9573 -18852 -9509 -18788
rect -9573 -18932 -9509 -18868
rect -9573 -19012 -9509 -18948
rect -9573 -19092 -9509 -19028
rect -9573 -19172 -9509 -19108
rect -9573 -19252 -9509 -19188
rect -9573 -19332 -9509 -19268
rect -9573 -19412 -9509 -19348
rect -9573 -19492 -9509 -19428
rect -9573 -19572 -9509 -19508
rect -9573 -19652 -9509 -19588
rect -9573 -19732 -9509 -19668
rect -9573 -19812 -9509 -19748
rect -9573 -19892 -9509 -19828
rect -9573 -19972 -9509 -19908
rect -9573 -20052 -9509 -19988
rect -9573 -20132 -9509 -20068
rect -9573 -20212 -9509 -20148
rect -9573 -20292 -9509 -20228
rect -9573 -20372 -9509 -20308
rect -9573 -20452 -9509 -20388
rect -9573 -20532 -9509 -20468
rect -9573 -20612 -9509 -20548
rect -9573 -20692 -9509 -20628
rect -9573 -20772 -9509 -20708
rect -9573 -20852 -9509 -20788
rect -9573 -20932 -9509 -20868
rect -9573 -21012 -9509 -20948
rect -9573 -21092 -9509 -21028
rect -9573 -21172 -9509 -21108
rect -9573 -21252 -9509 -21188
rect -9573 -21332 -9509 -21268
rect -9573 -21412 -9509 -21348
rect -9573 -21492 -9509 -21428
rect -9573 -21572 -9509 -21508
rect -9573 -21652 -9509 -21588
rect -9573 -21732 -9509 -21668
rect -9573 -21812 -9509 -21748
rect -9573 -21892 -9509 -21828
rect -9573 -21972 -9509 -21908
rect -3254 -15892 -3190 -15828
rect -3254 -15972 -3190 -15908
rect -3254 -16052 -3190 -15988
rect -3254 -16132 -3190 -16068
rect -3254 -16212 -3190 -16148
rect -3254 -16292 -3190 -16228
rect -3254 -16372 -3190 -16308
rect -3254 -16452 -3190 -16388
rect -3254 -16532 -3190 -16468
rect -3254 -16612 -3190 -16548
rect -3254 -16692 -3190 -16628
rect -3254 -16772 -3190 -16708
rect -3254 -16852 -3190 -16788
rect -3254 -16932 -3190 -16868
rect -3254 -17012 -3190 -16948
rect -3254 -17092 -3190 -17028
rect -3254 -17172 -3190 -17108
rect -3254 -17252 -3190 -17188
rect -3254 -17332 -3190 -17268
rect -3254 -17412 -3190 -17348
rect -3254 -17492 -3190 -17428
rect -3254 -17572 -3190 -17508
rect -3254 -17652 -3190 -17588
rect -3254 -17732 -3190 -17668
rect -3254 -17812 -3190 -17748
rect -3254 -17892 -3190 -17828
rect -3254 -17972 -3190 -17908
rect -3254 -18052 -3190 -17988
rect -3254 -18132 -3190 -18068
rect -3254 -18212 -3190 -18148
rect -3254 -18292 -3190 -18228
rect -3254 -18372 -3190 -18308
rect -3254 -18452 -3190 -18388
rect -3254 -18532 -3190 -18468
rect -3254 -18612 -3190 -18548
rect -3254 -18692 -3190 -18628
rect -3254 -18772 -3190 -18708
rect -3254 -18852 -3190 -18788
rect -3254 -18932 -3190 -18868
rect -3254 -19012 -3190 -18948
rect -3254 -19092 -3190 -19028
rect -3254 -19172 -3190 -19108
rect -3254 -19252 -3190 -19188
rect -3254 -19332 -3190 -19268
rect -3254 -19412 -3190 -19348
rect -3254 -19492 -3190 -19428
rect -3254 -19572 -3190 -19508
rect -3254 -19652 -3190 -19588
rect -3254 -19732 -3190 -19668
rect -3254 -19812 -3190 -19748
rect -3254 -19892 -3190 -19828
rect -3254 -19972 -3190 -19908
rect -3254 -20052 -3190 -19988
rect -3254 -20132 -3190 -20068
rect -3254 -20212 -3190 -20148
rect -3254 -20292 -3190 -20228
rect -3254 -20372 -3190 -20308
rect -3254 -20452 -3190 -20388
rect -3254 -20532 -3190 -20468
rect -3254 -20612 -3190 -20548
rect -3254 -20692 -3190 -20628
rect -3254 -20772 -3190 -20708
rect -3254 -20852 -3190 -20788
rect -3254 -20932 -3190 -20868
rect -3254 -21012 -3190 -20948
rect -3254 -21092 -3190 -21028
rect -3254 -21172 -3190 -21108
rect -3254 -21252 -3190 -21188
rect -3254 -21332 -3190 -21268
rect -3254 -21412 -3190 -21348
rect -3254 -21492 -3190 -21428
rect -3254 -21572 -3190 -21508
rect -3254 -21652 -3190 -21588
rect -3254 -21732 -3190 -21668
rect -3254 -21812 -3190 -21748
rect -3254 -21892 -3190 -21828
rect -3254 -21972 -3190 -21908
rect 3065 -15892 3129 -15828
rect 3065 -15972 3129 -15908
rect 3065 -16052 3129 -15988
rect 3065 -16132 3129 -16068
rect 3065 -16212 3129 -16148
rect 3065 -16292 3129 -16228
rect 3065 -16372 3129 -16308
rect 3065 -16452 3129 -16388
rect 3065 -16532 3129 -16468
rect 3065 -16612 3129 -16548
rect 3065 -16692 3129 -16628
rect 3065 -16772 3129 -16708
rect 3065 -16852 3129 -16788
rect 3065 -16932 3129 -16868
rect 3065 -17012 3129 -16948
rect 3065 -17092 3129 -17028
rect 3065 -17172 3129 -17108
rect 3065 -17252 3129 -17188
rect 3065 -17332 3129 -17268
rect 3065 -17412 3129 -17348
rect 3065 -17492 3129 -17428
rect 3065 -17572 3129 -17508
rect 3065 -17652 3129 -17588
rect 3065 -17732 3129 -17668
rect 3065 -17812 3129 -17748
rect 3065 -17892 3129 -17828
rect 3065 -17972 3129 -17908
rect 3065 -18052 3129 -17988
rect 3065 -18132 3129 -18068
rect 3065 -18212 3129 -18148
rect 3065 -18292 3129 -18228
rect 3065 -18372 3129 -18308
rect 3065 -18452 3129 -18388
rect 3065 -18532 3129 -18468
rect 3065 -18612 3129 -18548
rect 3065 -18692 3129 -18628
rect 3065 -18772 3129 -18708
rect 3065 -18852 3129 -18788
rect 3065 -18932 3129 -18868
rect 3065 -19012 3129 -18948
rect 3065 -19092 3129 -19028
rect 3065 -19172 3129 -19108
rect 3065 -19252 3129 -19188
rect 3065 -19332 3129 -19268
rect 3065 -19412 3129 -19348
rect 3065 -19492 3129 -19428
rect 3065 -19572 3129 -19508
rect 3065 -19652 3129 -19588
rect 3065 -19732 3129 -19668
rect 3065 -19812 3129 -19748
rect 3065 -19892 3129 -19828
rect 3065 -19972 3129 -19908
rect 3065 -20052 3129 -19988
rect 3065 -20132 3129 -20068
rect 3065 -20212 3129 -20148
rect 3065 -20292 3129 -20228
rect 3065 -20372 3129 -20308
rect 3065 -20452 3129 -20388
rect 3065 -20532 3129 -20468
rect 3065 -20612 3129 -20548
rect 3065 -20692 3129 -20628
rect 3065 -20772 3129 -20708
rect 3065 -20852 3129 -20788
rect 3065 -20932 3129 -20868
rect 3065 -21012 3129 -20948
rect 3065 -21092 3129 -21028
rect 3065 -21172 3129 -21108
rect 3065 -21252 3129 -21188
rect 3065 -21332 3129 -21268
rect 3065 -21412 3129 -21348
rect 3065 -21492 3129 -21428
rect 3065 -21572 3129 -21508
rect 3065 -21652 3129 -21588
rect 3065 -21732 3129 -21668
rect 3065 -21812 3129 -21748
rect 3065 -21892 3129 -21828
rect 3065 -21972 3129 -21908
rect 9384 -15892 9448 -15828
rect 9384 -15972 9448 -15908
rect 9384 -16052 9448 -15988
rect 9384 -16132 9448 -16068
rect 9384 -16212 9448 -16148
rect 9384 -16292 9448 -16228
rect 9384 -16372 9448 -16308
rect 9384 -16452 9448 -16388
rect 9384 -16532 9448 -16468
rect 9384 -16612 9448 -16548
rect 9384 -16692 9448 -16628
rect 9384 -16772 9448 -16708
rect 9384 -16852 9448 -16788
rect 9384 -16932 9448 -16868
rect 9384 -17012 9448 -16948
rect 9384 -17092 9448 -17028
rect 9384 -17172 9448 -17108
rect 9384 -17252 9448 -17188
rect 9384 -17332 9448 -17268
rect 9384 -17412 9448 -17348
rect 9384 -17492 9448 -17428
rect 9384 -17572 9448 -17508
rect 9384 -17652 9448 -17588
rect 9384 -17732 9448 -17668
rect 9384 -17812 9448 -17748
rect 9384 -17892 9448 -17828
rect 9384 -17972 9448 -17908
rect 9384 -18052 9448 -17988
rect 9384 -18132 9448 -18068
rect 9384 -18212 9448 -18148
rect 9384 -18292 9448 -18228
rect 9384 -18372 9448 -18308
rect 9384 -18452 9448 -18388
rect 9384 -18532 9448 -18468
rect 9384 -18612 9448 -18548
rect 9384 -18692 9448 -18628
rect 9384 -18772 9448 -18708
rect 9384 -18852 9448 -18788
rect 9384 -18932 9448 -18868
rect 9384 -19012 9448 -18948
rect 9384 -19092 9448 -19028
rect 9384 -19172 9448 -19108
rect 9384 -19252 9448 -19188
rect 9384 -19332 9448 -19268
rect 9384 -19412 9448 -19348
rect 9384 -19492 9448 -19428
rect 9384 -19572 9448 -19508
rect 9384 -19652 9448 -19588
rect 9384 -19732 9448 -19668
rect 9384 -19812 9448 -19748
rect 9384 -19892 9448 -19828
rect 9384 -19972 9448 -19908
rect 9384 -20052 9448 -19988
rect 9384 -20132 9448 -20068
rect 9384 -20212 9448 -20148
rect 9384 -20292 9448 -20228
rect 9384 -20372 9448 -20308
rect 9384 -20452 9448 -20388
rect 9384 -20532 9448 -20468
rect 9384 -20612 9448 -20548
rect 9384 -20692 9448 -20628
rect 9384 -20772 9448 -20708
rect 9384 -20852 9448 -20788
rect 9384 -20932 9448 -20868
rect 9384 -21012 9448 -20948
rect 9384 -21092 9448 -21028
rect 9384 -21172 9448 -21108
rect 9384 -21252 9448 -21188
rect 9384 -21332 9448 -21268
rect 9384 -21412 9448 -21348
rect 9384 -21492 9448 -21428
rect 9384 -21572 9448 -21508
rect 9384 -21652 9448 -21588
rect 9384 -21732 9448 -21668
rect 9384 -21812 9448 -21748
rect 9384 -21892 9448 -21828
rect 9384 -21972 9448 -21908
rect 15703 -15892 15767 -15828
rect 15703 -15972 15767 -15908
rect 15703 -16052 15767 -15988
rect 15703 -16132 15767 -16068
rect 15703 -16212 15767 -16148
rect 15703 -16292 15767 -16228
rect 15703 -16372 15767 -16308
rect 15703 -16452 15767 -16388
rect 15703 -16532 15767 -16468
rect 15703 -16612 15767 -16548
rect 15703 -16692 15767 -16628
rect 15703 -16772 15767 -16708
rect 15703 -16852 15767 -16788
rect 15703 -16932 15767 -16868
rect 15703 -17012 15767 -16948
rect 15703 -17092 15767 -17028
rect 15703 -17172 15767 -17108
rect 15703 -17252 15767 -17188
rect 15703 -17332 15767 -17268
rect 15703 -17412 15767 -17348
rect 15703 -17492 15767 -17428
rect 15703 -17572 15767 -17508
rect 15703 -17652 15767 -17588
rect 15703 -17732 15767 -17668
rect 15703 -17812 15767 -17748
rect 15703 -17892 15767 -17828
rect 15703 -17972 15767 -17908
rect 15703 -18052 15767 -17988
rect 15703 -18132 15767 -18068
rect 15703 -18212 15767 -18148
rect 15703 -18292 15767 -18228
rect 15703 -18372 15767 -18308
rect 15703 -18452 15767 -18388
rect 15703 -18532 15767 -18468
rect 15703 -18612 15767 -18548
rect 15703 -18692 15767 -18628
rect 15703 -18772 15767 -18708
rect 15703 -18852 15767 -18788
rect 15703 -18932 15767 -18868
rect 15703 -19012 15767 -18948
rect 15703 -19092 15767 -19028
rect 15703 -19172 15767 -19108
rect 15703 -19252 15767 -19188
rect 15703 -19332 15767 -19268
rect 15703 -19412 15767 -19348
rect 15703 -19492 15767 -19428
rect 15703 -19572 15767 -19508
rect 15703 -19652 15767 -19588
rect 15703 -19732 15767 -19668
rect 15703 -19812 15767 -19748
rect 15703 -19892 15767 -19828
rect 15703 -19972 15767 -19908
rect 15703 -20052 15767 -19988
rect 15703 -20132 15767 -20068
rect 15703 -20212 15767 -20148
rect 15703 -20292 15767 -20228
rect 15703 -20372 15767 -20308
rect 15703 -20452 15767 -20388
rect 15703 -20532 15767 -20468
rect 15703 -20612 15767 -20548
rect 15703 -20692 15767 -20628
rect 15703 -20772 15767 -20708
rect 15703 -20852 15767 -20788
rect 15703 -20932 15767 -20868
rect 15703 -21012 15767 -20948
rect 15703 -21092 15767 -21028
rect 15703 -21172 15767 -21108
rect 15703 -21252 15767 -21188
rect 15703 -21332 15767 -21268
rect 15703 -21412 15767 -21348
rect 15703 -21492 15767 -21428
rect 15703 -21572 15767 -21508
rect 15703 -21652 15767 -21588
rect 15703 -21732 15767 -21668
rect 15703 -21812 15767 -21748
rect 15703 -21892 15767 -21828
rect 15703 -21972 15767 -21908
rect 22022 -15892 22086 -15828
rect 22022 -15972 22086 -15908
rect 22022 -16052 22086 -15988
rect 22022 -16132 22086 -16068
rect 22022 -16212 22086 -16148
rect 22022 -16292 22086 -16228
rect 22022 -16372 22086 -16308
rect 22022 -16452 22086 -16388
rect 22022 -16532 22086 -16468
rect 22022 -16612 22086 -16548
rect 22022 -16692 22086 -16628
rect 22022 -16772 22086 -16708
rect 22022 -16852 22086 -16788
rect 22022 -16932 22086 -16868
rect 22022 -17012 22086 -16948
rect 22022 -17092 22086 -17028
rect 22022 -17172 22086 -17108
rect 22022 -17252 22086 -17188
rect 22022 -17332 22086 -17268
rect 22022 -17412 22086 -17348
rect 22022 -17492 22086 -17428
rect 22022 -17572 22086 -17508
rect 22022 -17652 22086 -17588
rect 22022 -17732 22086 -17668
rect 22022 -17812 22086 -17748
rect 22022 -17892 22086 -17828
rect 22022 -17972 22086 -17908
rect 22022 -18052 22086 -17988
rect 22022 -18132 22086 -18068
rect 22022 -18212 22086 -18148
rect 22022 -18292 22086 -18228
rect 22022 -18372 22086 -18308
rect 22022 -18452 22086 -18388
rect 22022 -18532 22086 -18468
rect 22022 -18612 22086 -18548
rect 22022 -18692 22086 -18628
rect 22022 -18772 22086 -18708
rect 22022 -18852 22086 -18788
rect 22022 -18932 22086 -18868
rect 22022 -19012 22086 -18948
rect 22022 -19092 22086 -19028
rect 22022 -19172 22086 -19108
rect 22022 -19252 22086 -19188
rect 22022 -19332 22086 -19268
rect 22022 -19412 22086 -19348
rect 22022 -19492 22086 -19428
rect 22022 -19572 22086 -19508
rect 22022 -19652 22086 -19588
rect 22022 -19732 22086 -19668
rect 22022 -19812 22086 -19748
rect 22022 -19892 22086 -19828
rect 22022 -19972 22086 -19908
rect 22022 -20052 22086 -19988
rect 22022 -20132 22086 -20068
rect 22022 -20212 22086 -20148
rect 22022 -20292 22086 -20228
rect 22022 -20372 22086 -20308
rect 22022 -20452 22086 -20388
rect 22022 -20532 22086 -20468
rect 22022 -20612 22086 -20548
rect 22022 -20692 22086 -20628
rect 22022 -20772 22086 -20708
rect 22022 -20852 22086 -20788
rect 22022 -20932 22086 -20868
rect 22022 -21012 22086 -20948
rect 22022 -21092 22086 -21028
rect 22022 -21172 22086 -21108
rect 22022 -21252 22086 -21188
rect 22022 -21332 22086 -21268
rect 22022 -21412 22086 -21348
rect 22022 -21492 22086 -21428
rect 22022 -21572 22086 -21508
rect 22022 -21652 22086 -21588
rect 22022 -21732 22086 -21668
rect 22022 -21812 22086 -21748
rect 22022 -21892 22086 -21828
rect 22022 -21972 22086 -21908
rect 28341 -15892 28405 -15828
rect 28341 -15972 28405 -15908
rect 28341 -16052 28405 -15988
rect 28341 -16132 28405 -16068
rect 28341 -16212 28405 -16148
rect 28341 -16292 28405 -16228
rect 28341 -16372 28405 -16308
rect 28341 -16452 28405 -16388
rect 28341 -16532 28405 -16468
rect 28341 -16612 28405 -16548
rect 28341 -16692 28405 -16628
rect 28341 -16772 28405 -16708
rect 28341 -16852 28405 -16788
rect 28341 -16932 28405 -16868
rect 28341 -17012 28405 -16948
rect 28341 -17092 28405 -17028
rect 28341 -17172 28405 -17108
rect 28341 -17252 28405 -17188
rect 28341 -17332 28405 -17268
rect 28341 -17412 28405 -17348
rect 28341 -17492 28405 -17428
rect 28341 -17572 28405 -17508
rect 28341 -17652 28405 -17588
rect 28341 -17732 28405 -17668
rect 28341 -17812 28405 -17748
rect 28341 -17892 28405 -17828
rect 28341 -17972 28405 -17908
rect 28341 -18052 28405 -17988
rect 28341 -18132 28405 -18068
rect 28341 -18212 28405 -18148
rect 28341 -18292 28405 -18228
rect 28341 -18372 28405 -18308
rect 28341 -18452 28405 -18388
rect 28341 -18532 28405 -18468
rect 28341 -18612 28405 -18548
rect 28341 -18692 28405 -18628
rect 28341 -18772 28405 -18708
rect 28341 -18852 28405 -18788
rect 28341 -18932 28405 -18868
rect 28341 -19012 28405 -18948
rect 28341 -19092 28405 -19028
rect 28341 -19172 28405 -19108
rect 28341 -19252 28405 -19188
rect 28341 -19332 28405 -19268
rect 28341 -19412 28405 -19348
rect 28341 -19492 28405 -19428
rect 28341 -19572 28405 -19508
rect 28341 -19652 28405 -19588
rect 28341 -19732 28405 -19668
rect 28341 -19812 28405 -19748
rect 28341 -19892 28405 -19828
rect 28341 -19972 28405 -19908
rect 28341 -20052 28405 -19988
rect 28341 -20132 28405 -20068
rect 28341 -20212 28405 -20148
rect 28341 -20292 28405 -20228
rect 28341 -20372 28405 -20308
rect 28341 -20452 28405 -20388
rect 28341 -20532 28405 -20468
rect 28341 -20612 28405 -20548
rect 28341 -20692 28405 -20628
rect 28341 -20772 28405 -20708
rect 28341 -20852 28405 -20788
rect 28341 -20932 28405 -20868
rect 28341 -21012 28405 -20948
rect 28341 -21092 28405 -21028
rect 28341 -21172 28405 -21108
rect 28341 -21252 28405 -21188
rect 28341 -21332 28405 -21268
rect 28341 -21412 28405 -21348
rect 28341 -21492 28405 -21428
rect 28341 -21572 28405 -21508
rect 28341 -21652 28405 -21588
rect 28341 -21732 28405 -21668
rect 28341 -21812 28405 -21748
rect 28341 -21892 28405 -21828
rect 28341 -21972 28405 -21908
rect 34660 -15892 34724 -15828
rect 34660 -15972 34724 -15908
rect 34660 -16052 34724 -15988
rect 34660 -16132 34724 -16068
rect 34660 -16212 34724 -16148
rect 34660 -16292 34724 -16228
rect 34660 -16372 34724 -16308
rect 34660 -16452 34724 -16388
rect 34660 -16532 34724 -16468
rect 34660 -16612 34724 -16548
rect 34660 -16692 34724 -16628
rect 34660 -16772 34724 -16708
rect 34660 -16852 34724 -16788
rect 34660 -16932 34724 -16868
rect 34660 -17012 34724 -16948
rect 34660 -17092 34724 -17028
rect 34660 -17172 34724 -17108
rect 34660 -17252 34724 -17188
rect 34660 -17332 34724 -17268
rect 34660 -17412 34724 -17348
rect 34660 -17492 34724 -17428
rect 34660 -17572 34724 -17508
rect 34660 -17652 34724 -17588
rect 34660 -17732 34724 -17668
rect 34660 -17812 34724 -17748
rect 34660 -17892 34724 -17828
rect 34660 -17972 34724 -17908
rect 34660 -18052 34724 -17988
rect 34660 -18132 34724 -18068
rect 34660 -18212 34724 -18148
rect 34660 -18292 34724 -18228
rect 34660 -18372 34724 -18308
rect 34660 -18452 34724 -18388
rect 34660 -18532 34724 -18468
rect 34660 -18612 34724 -18548
rect 34660 -18692 34724 -18628
rect 34660 -18772 34724 -18708
rect 34660 -18852 34724 -18788
rect 34660 -18932 34724 -18868
rect 34660 -19012 34724 -18948
rect 34660 -19092 34724 -19028
rect 34660 -19172 34724 -19108
rect 34660 -19252 34724 -19188
rect 34660 -19332 34724 -19268
rect 34660 -19412 34724 -19348
rect 34660 -19492 34724 -19428
rect 34660 -19572 34724 -19508
rect 34660 -19652 34724 -19588
rect 34660 -19732 34724 -19668
rect 34660 -19812 34724 -19748
rect 34660 -19892 34724 -19828
rect 34660 -19972 34724 -19908
rect 34660 -20052 34724 -19988
rect 34660 -20132 34724 -20068
rect 34660 -20212 34724 -20148
rect 34660 -20292 34724 -20228
rect 34660 -20372 34724 -20308
rect 34660 -20452 34724 -20388
rect 34660 -20532 34724 -20468
rect 34660 -20612 34724 -20548
rect 34660 -20692 34724 -20628
rect 34660 -20772 34724 -20708
rect 34660 -20852 34724 -20788
rect 34660 -20932 34724 -20868
rect 34660 -21012 34724 -20948
rect 34660 -21092 34724 -21028
rect 34660 -21172 34724 -21108
rect 34660 -21252 34724 -21188
rect 34660 -21332 34724 -21268
rect 34660 -21412 34724 -21348
rect 34660 -21492 34724 -21428
rect 34660 -21572 34724 -21508
rect 34660 -21652 34724 -21588
rect 34660 -21732 34724 -21668
rect 34660 -21812 34724 -21748
rect 34660 -21892 34724 -21828
rect 34660 -21972 34724 -21908
rect 40979 -15892 41043 -15828
rect 40979 -15972 41043 -15908
rect 40979 -16052 41043 -15988
rect 40979 -16132 41043 -16068
rect 40979 -16212 41043 -16148
rect 40979 -16292 41043 -16228
rect 40979 -16372 41043 -16308
rect 40979 -16452 41043 -16388
rect 40979 -16532 41043 -16468
rect 40979 -16612 41043 -16548
rect 40979 -16692 41043 -16628
rect 40979 -16772 41043 -16708
rect 40979 -16852 41043 -16788
rect 40979 -16932 41043 -16868
rect 40979 -17012 41043 -16948
rect 40979 -17092 41043 -17028
rect 40979 -17172 41043 -17108
rect 40979 -17252 41043 -17188
rect 40979 -17332 41043 -17268
rect 40979 -17412 41043 -17348
rect 40979 -17492 41043 -17428
rect 40979 -17572 41043 -17508
rect 40979 -17652 41043 -17588
rect 40979 -17732 41043 -17668
rect 40979 -17812 41043 -17748
rect 40979 -17892 41043 -17828
rect 40979 -17972 41043 -17908
rect 40979 -18052 41043 -17988
rect 40979 -18132 41043 -18068
rect 40979 -18212 41043 -18148
rect 40979 -18292 41043 -18228
rect 40979 -18372 41043 -18308
rect 40979 -18452 41043 -18388
rect 40979 -18532 41043 -18468
rect 40979 -18612 41043 -18548
rect 40979 -18692 41043 -18628
rect 40979 -18772 41043 -18708
rect 40979 -18852 41043 -18788
rect 40979 -18932 41043 -18868
rect 40979 -19012 41043 -18948
rect 40979 -19092 41043 -19028
rect 40979 -19172 41043 -19108
rect 40979 -19252 41043 -19188
rect 40979 -19332 41043 -19268
rect 40979 -19412 41043 -19348
rect 40979 -19492 41043 -19428
rect 40979 -19572 41043 -19508
rect 40979 -19652 41043 -19588
rect 40979 -19732 41043 -19668
rect 40979 -19812 41043 -19748
rect 40979 -19892 41043 -19828
rect 40979 -19972 41043 -19908
rect 40979 -20052 41043 -19988
rect 40979 -20132 41043 -20068
rect 40979 -20212 41043 -20148
rect 40979 -20292 41043 -20228
rect 40979 -20372 41043 -20308
rect 40979 -20452 41043 -20388
rect 40979 -20532 41043 -20468
rect 40979 -20612 41043 -20548
rect 40979 -20692 41043 -20628
rect 40979 -20772 41043 -20708
rect 40979 -20852 41043 -20788
rect 40979 -20932 41043 -20868
rect 40979 -21012 41043 -20948
rect 40979 -21092 41043 -21028
rect 40979 -21172 41043 -21108
rect 40979 -21252 41043 -21188
rect 40979 -21332 41043 -21268
rect 40979 -21412 41043 -21348
rect 40979 -21492 41043 -21428
rect 40979 -21572 41043 -21508
rect 40979 -21652 41043 -21588
rect 40979 -21732 41043 -21668
rect 40979 -21812 41043 -21748
rect 40979 -21892 41043 -21828
rect 40979 -21972 41043 -21908
rect 47298 -15892 47362 -15828
rect 47298 -15972 47362 -15908
rect 47298 -16052 47362 -15988
rect 47298 -16132 47362 -16068
rect 47298 -16212 47362 -16148
rect 47298 -16292 47362 -16228
rect 47298 -16372 47362 -16308
rect 47298 -16452 47362 -16388
rect 47298 -16532 47362 -16468
rect 47298 -16612 47362 -16548
rect 47298 -16692 47362 -16628
rect 47298 -16772 47362 -16708
rect 47298 -16852 47362 -16788
rect 47298 -16932 47362 -16868
rect 47298 -17012 47362 -16948
rect 47298 -17092 47362 -17028
rect 47298 -17172 47362 -17108
rect 47298 -17252 47362 -17188
rect 47298 -17332 47362 -17268
rect 47298 -17412 47362 -17348
rect 47298 -17492 47362 -17428
rect 47298 -17572 47362 -17508
rect 47298 -17652 47362 -17588
rect 47298 -17732 47362 -17668
rect 47298 -17812 47362 -17748
rect 47298 -17892 47362 -17828
rect 47298 -17972 47362 -17908
rect 47298 -18052 47362 -17988
rect 47298 -18132 47362 -18068
rect 47298 -18212 47362 -18148
rect 47298 -18292 47362 -18228
rect 47298 -18372 47362 -18308
rect 47298 -18452 47362 -18388
rect 47298 -18532 47362 -18468
rect 47298 -18612 47362 -18548
rect 47298 -18692 47362 -18628
rect 47298 -18772 47362 -18708
rect 47298 -18852 47362 -18788
rect 47298 -18932 47362 -18868
rect 47298 -19012 47362 -18948
rect 47298 -19092 47362 -19028
rect 47298 -19172 47362 -19108
rect 47298 -19252 47362 -19188
rect 47298 -19332 47362 -19268
rect 47298 -19412 47362 -19348
rect 47298 -19492 47362 -19428
rect 47298 -19572 47362 -19508
rect 47298 -19652 47362 -19588
rect 47298 -19732 47362 -19668
rect 47298 -19812 47362 -19748
rect 47298 -19892 47362 -19828
rect 47298 -19972 47362 -19908
rect 47298 -20052 47362 -19988
rect 47298 -20132 47362 -20068
rect 47298 -20212 47362 -20148
rect 47298 -20292 47362 -20228
rect 47298 -20372 47362 -20308
rect 47298 -20452 47362 -20388
rect 47298 -20532 47362 -20468
rect 47298 -20612 47362 -20548
rect 47298 -20692 47362 -20628
rect 47298 -20772 47362 -20708
rect 47298 -20852 47362 -20788
rect 47298 -20932 47362 -20868
rect 47298 -21012 47362 -20948
rect 47298 -21092 47362 -21028
rect 47298 -21172 47362 -21108
rect 47298 -21252 47362 -21188
rect 47298 -21332 47362 -21268
rect 47298 -21412 47362 -21348
rect 47298 -21492 47362 -21428
rect 47298 -21572 47362 -21508
rect 47298 -21652 47362 -21588
rect 47298 -21732 47362 -21668
rect 47298 -21812 47362 -21748
rect 47298 -21892 47362 -21828
rect 47298 -21972 47362 -21908
rect -41168 -22192 -41104 -22128
rect -41168 -22272 -41104 -22208
rect -41168 -22352 -41104 -22288
rect -41168 -22432 -41104 -22368
rect -41168 -22512 -41104 -22448
rect -41168 -22592 -41104 -22528
rect -41168 -22672 -41104 -22608
rect -41168 -22752 -41104 -22688
rect -41168 -22832 -41104 -22768
rect -41168 -22912 -41104 -22848
rect -41168 -22992 -41104 -22928
rect -41168 -23072 -41104 -23008
rect -41168 -23152 -41104 -23088
rect -41168 -23232 -41104 -23168
rect -41168 -23312 -41104 -23248
rect -41168 -23392 -41104 -23328
rect -41168 -23472 -41104 -23408
rect -41168 -23552 -41104 -23488
rect -41168 -23632 -41104 -23568
rect -41168 -23712 -41104 -23648
rect -41168 -23792 -41104 -23728
rect -41168 -23872 -41104 -23808
rect -41168 -23952 -41104 -23888
rect -41168 -24032 -41104 -23968
rect -41168 -24112 -41104 -24048
rect -41168 -24192 -41104 -24128
rect -41168 -24272 -41104 -24208
rect -41168 -24352 -41104 -24288
rect -41168 -24432 -41104 -24368
rect -41168 -24512 -41104 -24448
rect -41168 -24592 -41104 -24528
rect -41168 -24672 -41104 -24608
rect -41168 -24752 -41104 -24688
rect -41168 -24832 -41104 -24768
rect -41168 -24912 -41104 -24848
rect -41168 -24992 -41104 -24928
rect -41168 -25072 -41104 -25008
rect -41168 -25152 -41104 -25088
rect -41168 -25232 -41104 -25168
rect -41168 -25312 -41104 -25248
rect -41168 -25392 -41104 -25328
rect -41168 -25472 -41104 -25408
rect -41168 -25552 -41104 -25488
rect -41168 -25632 -41104 -25568
rect -41168 -25712 -41104 -25648
rect -41168 -25792 -41104 -25728
rect -41168 -25872 -41104 -25808
rect -41168 -25952 -41104 -25888
rect -41168 -26032 -41104 -25968
rect -41168 -26112 -41104 -26048
rect -41168 -26192 -41104 -26128
rect -41168 -26272 -41104 -26208
rect -41168 -26352 -41104 -26288
rect -41168 -26432 -41104 -26368
rect -41168 -26512 -41104 -26448
rect -41168 -26592 -41104 -26528
rect -41168 -26672 -41104 -26608
rect -41168 -26752 -41104 -26688
rect -41168 -26832 -41104 -26768
rect -41168 -26912 -41104 -26848
rect -41168 -26992 -41104 -26928
rect -41168 -27072 -41104 -27008
rect -41168 -27152 -41104 -27088
rect -41168 -27232 -41104 -27168
rect -41168 -27312 -41104 -27248
rect -41168 -27392 -41104 -27328
rect -41168 -27472 -41104 -27408
rect -41168 -27552 -41104 -27488
rect -41168 -27632 -41104 -27568
rect -41168 -27712 -41104 -27648
rect -41168 -27792 -41104 -27728
rect -41168 -27872 -41104 -27808
rect -41168 -27952 -41104 -27888
rect -41168 -28032 -41104 -27968
rect -41168 -28112 -41104 -28048
rect -41168 -28192 -41104 -28128
rect -41168 -28272 -41104 -28208
rect -34849 -22192 -34785 -22128
rect -34849 -22272 -34785 -22208
rect -34849 -22352 -34785 -22288
rect -34849 -22432 -34785 -22368
rect -34849 -22512 -34785 -22448
rect -34849 -22592 -34785 -22528
rect -34849 -22672 -34785 -22608
rect -34849 -22752 -34785 -22688
rect -34849 -22832 -34785 -22768
rect -34849 -22912 -34785 -22848
rect -34849 -22992 -34785 -22928
rect -34849 -23072 -34785 -23008
rect -34849 -23152 -34785 -23088
rect -34849 -23232 -34785 -23168
rect -34849 -23312 -34785 -23248
rect -34849 -23392 -34785 -23328
rect -34849 -23472 -34785 -23408
rect -34849 -23552 -34785 -23488
rect -34849 -23632 -34785 -23568
rect -34849 -23712 -34785 -23648
rect -34849 -23792 -34785 -23728
rect -34849 -23872 -34785 -23808
rect -34849 -23952 -34785 -23888
rect -34849 -24032 -34785 -23968
rect -34849 -24112 -34785 -24048
rect -34849 -24192 -34785 -24128
rect -34849 -24272 -34785 -24208
rect -34849 -24352 -34785 -24288
rect -34849 -24432 -34785 -24368
rect -34849 -24512 -34785 -24448
rect -34849 -24592 -34785 -24528
rect -34849 -24672 -34785 -24608
rect -34849 -24752 -34785 -24688
rect -34849 -24832 -34785 -24768
rect -34849 -24912 -34785 -24848
rect -34849 -24992 -34785 -24928
rect -34849 -25072 -34785 -25008
rect -34849 -25152 -34785 -25088
rect -34849 -25232 -34785 -25168
rect -34849 -25312 -34785 -25248
rect -34849 -25392 -34785 -25328
rect -34849 -25472 -34785 -25408
rect -34849 -25552 -34785 -25488
rect -34849 -25632 -34785 -25568
rect -34849 -25712 -34785 -25648
rect -34849 -25792 -34785 -25728
rect -34849 -25872 -34785 -25808
rect -34849 -25952 -34785 -25888
rect -34849 -26032 -34785 -25968
rect -34849 -26112 -34785 -26048
rect -34849 -26192 -34785 -26128
rect -34849 -26272 -34785 -26208
rect -34849 -26352 -34785 -26288
rect -34849 -26432 -34785 -26368
rect -34849 -26512 -34785 -26448
rect -34849 -26592 -34785 -26528
rect -34849 -26672 -34785 -26608
rect -34849 -26752 -34785 -26688
rect -34849 -26832 -34785 -26768
rect -34849 -26912 -34785 -26848
rect -34849 -26992 -34785 -26928
rect -34849 -27072 -34785 -27008
rect -34849 -27152 -34785 -27088
rect -34849 -27232 -34785 -27168
rect -34849 -27312 -34785 -27248
rect -34849 -27392 -34785 -27328
rect -34849 -27472 -34785 -27408
rect -34849 -27552 -34785 -27488
rect -34849 -27632 -34785 -27568
rect -34849 -27712 -34785 -27648
rect -34849 -27792 -34785 -27728
rect -34849 -27872 -34785 -27808
rect -34849 -27952 -34785 -27888
rect -34849 -28032 -34785 -27968
rect -34849 -28112 -34785 -28048
rect -34849 -28192 -34785 -28128
rect -34849 -28272 -34785 -28208
rect -28530 -22192 -28466 -22128
rect -28530 -22272 -28466 -22208
rect -28530 -22352 -28466 -22288
rect -28530 -22432 -28466 -22368
rect -28530 -22512 -28466 -22448
rect -28530 -22592 -28466 -22528
rect -28530 -22672 -28466 -22608
rect -28530 -22752 -28466 -22688
rect -28530 -22832 -28466 -22768
rect -28530 -22912 -28466 -22848
rect -28530 -22992 -28466 -22928
rect -28530 -23072 -28466 -23008
rect -28530 -23152 -28466 -23088
rect -28530 -23232 -28466 -23168
rect -28530 -23312 -28466 -23248
rect -28530 -23392 -28466 -23328
rect -28530 -23472 -28466 -23408
rect -28530 -23552 -28466 -23488
rect -28530 -23632 -28466 -23568
rect -28530 -23712 -28466 -23648
rect -28530 -23792 -28466 -23728
rect -28530 -23872 -28466 -23808
rect -28530 -23952 -28466 -23888
rect -28530 -24032 -28466 -23968
rect -28530 -24112 -28466 -24048
rect -28530 -24192 -28466 -24128
rect -28530 -24272 -28466 -24208
rect -28530 -24352 -28466 -24288
rect -28530 -24432 -28466 -24368
rect -28530 -24512 -28466 -24448
rect -28530 -24592 -28466 -24528
rect -28530 -24672 -28466 -24608
rect -28530 -24752 -28466 -24688
rect -28530 -24832 -28466 -24768
rect -28530 -24912 -28466 -24848
rect -28530 -24992 -28466 -24928
rect -28530 -25072 -28466 -25008
rect -28530 -25152 -28466 -25088
rect -28530 -25232 -28466 -25168
rect -28530 -25312 -28466 -25248
rect -28530 -25392 -28466 -25328
rect -28530 -25472 -28466 -25408
rect -28530 -25552 -28466 -25488
rect -28530 -25632 -28466 -25568
rect -28530 -25712 -28466 -25648
rect -28530 -25792 -28466 -25728
rect -28530 -25872 -28466 -25808
rect -28530 -25952 -28466 -25888
rect -28530 -26032 -28466 -25968
rect -28530 -26112 -28466 -26048
rect -28530 -26192 -28466 -26128
rect -28530 -26272 -28466 -26208
rect -28530 -26352 -28466 -26288
rect -28530 -26432 -28466 -26368
rect -28530 -26512 -28466 -26448
rect -28530 -26592 -28466 -26528
rect -28530 -26672 -28466 -26608
rect -28530 -26752 -28466 -26688
rect -28530 -26832 -28466 -26768
rect -28530 -26912 -28466 -26848
rect -28530 -26992 -28466 -26928
rect -28530 -27072 -28466 -27008
rect -28530 -27152 -28466 -27088
rect -28530 -27232 -28466 -27168
rect -28530 -27312 -28466 -27248
rect -28530 -27392 -28466 -27328
rect -28530 -27472 -28466 -27408
rect -28530 -27552 -28466 -27488
rect -28530 -27632 -28466 -27568
rect -28530 -27712 -28466 -27648
rect -28530 -27792 -28466 -27728
rect -28530 -27872 -28466 -27808
rect -28530 -27952 -28466 -27888
rect -28530 -28032 -28466 -27968
rect -28530 -28112 -28466 -28048
rect -28530 -28192 -28466 -28128
rect -28530 -28272 -28466 -28208
rect -22211 -22192 -22147 -22128
rect -22211 -22272 -22147 -22208
rect -22211 -22352 -22147 -22288
rect -22211 -22432 -22147 -22368
rect -22211 -22512 -22147 -22448
rect -22211 -22592 -22147 -22528
rect -22211 -22672 -22147 -22608
rect -22211 -22752 -22147 -22688
rect -22211 -22832 -22147 -22768
rect -22211 -22912 -22147 -22848
rect -22211 -22992 -22147 -22928
rect -22211 -23072 -22147 -23008
rect -22211 -23152 -22147 -23088
rect -22211 -23232 -22147 -23168
rect -22211 -23312 -22147 -23248
rect -22211 -23392 -22147 -23328
rect -22211 -23472 -22147 -23408
rect -22211 -23552 -22147 -23488
rect -22211 -23632 -22147 -23568
rect -22211 -23712 -22147 -23648
rect -22211 -23792 -22147 -23728
rect -22211 -23872 -22147 -23808
rect -22211 -23952 -22147 -23888
rect -22211 -24032 -22147 -23968
rect -22211 -24112 -22147 -24048
rect -22211 -24192 -22147 -24128
rect -22211 -24272 -22147 -24208
rect -22211 -24352 -22147 -24288
rect -22211 -24432 -22147 -24368
rect -22211 -24512 -22147 -24448
rect -22211 -24592 -22147 -24528
rect -22211 -24672 -22147 -24608
rect -22211 -24752 -22147 -24688
rect -22211 -24832 -22147 -24768
rect -22211 -24912 -22147 -24848
rect -22211 -24992 -22147 -24928
rect -22211 -25072 -22147 -25008
rect -22211 -25152 -22147 -25088
rect -22211 -25232 -22147 -25168
rect -22211 -25312 -22147 -25248
rect -22211 -25392 -22147 -25328
rect -22211 -25472 -22147 -25408
rect -22211 -25552 -22147 -25488
rect -22211 -25632 -22147 -25568
rect -22211 -25712 -22147 -25648
rect -22211 -25792 -22147 -25728
rect -22211 -25872 -22147 -25808
rect -22211 -25952 -22147 -25888
rect -22211 -26032 -22147 -25968
rect -22211 -26112 -22147 -26048
rect -22211 -26192 -22147 -26128
rect -22211 -26272 -22147 -26208
rect -22211 -26352 -22147 -26288
rect -22211 -26432 -22147 -26368
rect -22211 -26512 -22147 -26448
rect -22211 -26592 -22147 -26528
rect -22211 -26672 -22147 -26608
rect -22211 -26752 -22147 -26688
rect -22211 -26832 -22147 -26768
rect -22211 -26912 -22147 -26848
rect -22211 -26992 -22147 -26928
rect -22211 -27072 -22147 -27008
rect -22211 -27152 -22147 -27088
rect -22211 -27232 -22147 -27168
rect -22211 -27312 -22147 -27248
rect -22211 -27392 -22147 -27328
rect -22211 -27472 -22147 -27408
rect -22211 -27552 -22147 -27488
rect -22211 -27632 -22147 -27568
rect -22211 -27712 -22147 -27648
rect -22211 -27792 -22147 -27728
rect -22211 -27872 -22147 -27808
rect -22211 -27952 -22147 -27888
rect -22211 -28032 -22147 -27968
rect -22211 -28112 -22147 -28048
rect -22211 -28192 -22147 -28128
rect -22211 -28272 -22147 -28208
rect -15892 -22192 -15828 -22128
rect -15892 -22272 -15828 -22208
rect -15892 -22352 -15828 -22288
rect -15892 -22432 -15828 -22368
rect -15892 -22512 -15828 -22448
rect -15892 -22592 -15828 -22528
rect -15892 -22672 -15828 -22608
rect -15892 -22752 -15828 -22688
rect -15892 -22832 -15828 -22768
rect -15892 -22912 -15828 -22848
rect -15892 -22992 -15828 -22928
rect -15892 -23072 -15828 -23008
rect -15892 -23152 -15828 -23088
rect -15892 -23232 -15828 -23168
rect -15892 -23312 -15828 -23248
rect -15892 -23392 -15828 -23328
rect -15892 -23472 -15828 -23408
rect -15892 -23552 -15828 -23488
rect -15892 -23632 -15828 -23568
rect -15892 -23712 -15828 -23648
rect -15892 -23792 -15828 -23728
rect -15892 -23872 -15828 -23808
rect -15892 -23952 -15828 -23888
rect -15892 -24032 -15828 -23968
rect -15892 -24112 -15828 -24048
rect -15892 -24192 -15828 -24128
rect -15892 -24272 -15828 -24208
rect -15892 -24352 -15828 -24288
rect -15892 -24432 -15828 -24368
rect -15892 -24512 -15828 -24448
rect -15892 -24592 -15828 -24528
rect -15892 -24672 -15828 -24608
rect -15892 -24752 -15828 -24688
rect -15892 -24832 -15828 -24768
rect -15892 -24912 -15828 -24848
rect -15892 -24992 -15828 -24928
rect -15892 -25072 -15828 -25008
rect -15892 -25152 -15828 -25088
rect -15892 -25232 -15828 -25168
rect -15892 -25312 -15828 -25248
rect -15892 -25392 -15828 -25328
rect -15892 -25472 -15828 -25408
rect -15892 -25552 -15828 -25488
rect -15892 -25632 -15828 -25568
rect -15892 -25712 -15828 -25648
rect -15892 -25792 -15828 -25728
rect -15892 -25872 -15828 -25808
rect -15892 -25952 -15828 -25888
rect -15892 -26032 -15828 -25968
rect -15892 -26112 -15828 -26048
rect -15892 -26192 -15828 -26128
rect -15892 -26272 -15828 -26208
rect -15892 -26352 -15828 -26288
rect -15892 -26432 -15828 -26368
rect -15892 -26512 -15828 -26448
rect -15892 -26592 -15828 -26528
rect -15892 -26672 -15828 -26608
rect -15892 -26752 -15828 -26688
rect -15892 -26832 -15828 -26768
rect -15892 -26912 -15828 -26848
rect -15892 -26992 -15828 -26928
rect -15892 -27072 -15828 -27008
rect -15892 -27152 -15828 -27088
rect -15892 -27232 -15828 -27168
rect -15892 -27312 -15828 -27248
rect -15892 -27392 -15828 -27328
rect -15892 -27472 -15828 -27408
rect -15892 -27552 -15828 -27488
rect -15892 -27632 -15828 -27568
rect -15892 -27712 -15828 -27648
rect -15892 -27792 -15828 -27728
rect -15892 -27872 -15828 -27808
rect -15892 -27952 -15828 -27888
rect -15892 -28032 -15828 -27968
rect -15892 -28112 -15828 -28048
rect -15892 -28192 -15828 -28128
rect -15892 -28272 -15828 -28208
rect -9573 -22192 -9509 -22128
rect -9573 -22272 -9509 -22208
rect -9573 -22352 -9509 -22288
rect -9573 -22432 -9509 -22368
rect -9573 -22512 -9509 -22448
rect -9573 -22592 -9509 -22528
rect -9573 -22672 -9509 -22608
rect -9573 -22752 -9509 -22688
rect -9573 -22832 -9509 -22768
rect -9573 -22912 -9509 -22848
rect -9573 -22992 -9509 -22928
rect -9573 -23072 -9509 -23008
rect -9573 -23152 -9509 -23088
rect -9573 -23232 -9509 -23168
rect -9573 -23312 -9509 -23248
rect -9573 -23392 -9509 -23328
rect -9573 -23472 -9509 -23408
rect -9573 -23552 -9509 -23488
rect -9573 -23632 -9509 -23568
rect -9573 -23712 -9509 -23648
rect -9573 -23792 -9509 -23728
rect -9573 -23872 -9509 -23808
rect -9573 -23952 -9509 -23888
rect -9573 -24032 -9509 -23968
rect -9573 -24112 -9509 -24048
rect -9573 -24192 -9509 -24128
rect -9573 -24272 -9509 -24208
rect -9573 -24352 -9509 -24288
rect -9573 -24432 -9509 -24368
rect -9573 -24512 -9509 -24448
rect -9573 -24592 -9509 -24528
rect -9573 -24672 -9509 -24608
rect -9573 -24752 -9509 -24688
rect -9573 -24832 -9509 -24768
rect -9573 -24912 -9509 -24848
rect -9573 -24992 -9509 -24928
rect -9573 -25072 -9509 -25008
rect -9573 -25152 -9509 -25088
rect -9573 -25232 -9509 -25168
rect -9573 -25312 -9509 -25248
rect -9573 -25392 -9509 -25328
rect -9573 -25472 -9509 -25408
rect -9573 -25552 -9509 -25488
rect -9573 -25632 -9509 -25568
rect -9573 -25712 -9509 -25648
rect -9573 -25792 -9509 -25728
rect -9573 -25872 -9509 -25808
rect -9573 -25952 -9509 -25888
rect -9573 -26032 -9509 -25968
rect -9573 -26112 -9509 -26048
rect -9573 -26192 -9509 -26128
rect -9573 -26272 -9509 -26208
rect -9573 -26352 -9509 -26288
rect -9573 -26432 -9509 -26368
rect -9573 -26512 -9509 -26448
rect -9573 -26592 -9509 -26528
rect -9573 -26672 -9509 -26608
rect -9573 -26752 -9509 -26688
rect -9573 -26832 -9509 -26768
rect -9573 -26912 -9509 -26848
rect -9573 -26992 -9509 -26928
rect -9573 -27072 -9509 -27008
rect -9573 -27152 -9509 -27088
rect -9573 -27232 -9509 -27168
rect -9573 -27312 -9509 -27248
rect -9573 -27392 -9509 -27328
rect -9573 -27472 -9509 -27408
rect -9573 -27552 -9509 -27488
rect -9573 -27632 -9509 -27568
rect -9573 -27712 -9509 -27648
rect -9573 -27792 -9509 -27728
rect -9573 -27872 -9509 -27808
rect -9573 -27952 -9509 -27888
rect -9573 -28032 -9509 -27968
rect -9573 -28112 -9509 -28048
rect -9573 -28192 -9509 -28128
rect -9573 -28272 -9509 -28208
rect -3254 -22192 -3190 -22128
rect -3254 -22272 -3190 -22208
rect -3254 -22352 -3190 -22288
rect -3254 -22432 -3190 -22368
rect -3254 -22512 -3190 -22448
rect -3254 -22592 -3190 -22528
rect -3254 -22672 -3190 -22608
rect -3254 -22752 -3190 -22688
rect -3254 -22832 -3190 -22768
rect -3254 -22912 -3190 -22848
rect -3254 -22992 -3190 -22928
rect -3254 -23072 -3190 -23008
rect -3254 -23152 -3190 -23088
rect -3254 -23232 -3190 -23168
rect -3254 -23312 -3190 -23248
rect -3254 -23392 -3190 -23328
rect -3254 -23472 -3190 -23408
rect -3254 -23552 -3190 -23488
rect -3254 -23632 -3190 -23568
rect -3254 -23712 -3190 -23648
rect -3254 -23792 -3190 -23728
rect -3254 -23872 -3190 -23808
rect -3254 -23952 -3190 -23888
rect -3254 -24032 -3190 -23968
rect -3254 -24112 -3190 -24048
rect -3254 -24192 -3190 -24128
rect -3254 -24272 -3190 -24208
rect -3254 -24352 -3190 -24288
rect -3254 -24432 -3190 -24368
rect -3254 -24512 -3190 -24448
rect -3254 -24592 -3190 -24528
rect -3254 -24672 -3190 -24608
rect -3254 -24752 -3190 -24688
rect -3254 -24832 -3190 -24768
rect -3254 -24912 -3190 -24848
rect -3254 -24992 -3190 -24928
rect -3254 -25072 -3190 -25008
rect -3254 -25152 -3190 -25088
rect -3254 -25232 -3190 -25168
rect -3254 -25312 -3190 -25248
rect -3254 -25392 -3190 -25328
rect -3254 -25472 -3190 -25408
rect -3254 -25552 -3190 -25488
rect -3254 -25632 -3190 -25568
rect -3254 -25712 -3190 -25648
rect -3254 -25792 -3190 -25728
rect -3254 -25872 -3190 -25808
rect -3254 -25952 -3190 -25888
rect -3254 -26032 -3190 -25968
rect -3254 -26112 -3190 -26048
rect -3254 -26192 -3190 -26128
rect -3254 -26272 -3190 -26208
rect -3254 -26352 -3190 -26288
rect -3254 -26432 -3190 -26368
rect -3254 -26512 -3190 -26448
rect -3254 -26592 -3190 -26528
rect -3254 -26672 -3190 -26608
rect -3254 -26752 -3190 -26688
rect -3254 -26832 -3190 -26768
rect -3254 -26912 -3190 -26848
rect -3254 -26992 -3190 -26928
rect -3254 -27072 -3190 -27008
rect -3254 -27152 -3190 -27088
rect -3254 -27232 -3190 -27168
rect -3254 -27312 -3190 -27248
rect -3254 -27392 -3190 -27328
rect -3254 -27472 -3190 -27408
rect -3254 -27552 -3190 -27488
rect -3254 -27632 -3190 -27568
rect -3254 -27712 -3190 -27648
rect -3254 -27792 -3190 -27728
rect -3254 -27872 -3190 -27808
rect -3254 -27952 -3190 -27888
rect -3254 -28032 -3190 -27968
rect -3254 -28112 -3190 -28048
rect -3254 -28192 -3190 -28128
rect -3254 -28272 -3190 -28208
rect 3065 -22192 3129 -22128
rect 3065 -22272 3129 -22208
rect 3065 -22352 3129 -22288
rect 3065 -22432 3129 -22368
rect 3065 -22512 3129 -22448
rect 3065 -22592 3129 -22528
rect 3065 -22672 3129 -22608
rect 3065 -22752 3129 -22688
rect 3065 -22832 3129 -22768
rect 3065 -22912 3129 -22848
rect 3065 -22992 3129 -22928
rect 3065 -23072 3129 -23008
rect 3065 -23152 3129 -23088
rect 3065 -23232 3129 -23168
rect 3065 -23312 3129 -23248
rect 3065 -23392 3129 -23328
rect 3065 -23472 3129 -23408
rect 3065 -23552 3129 -23488
rect 3065 -23632 3129 -23568
rect 3065 -23712 3129 -23648
rect 3065 -23792 3129 -23728
rect 3065 -23872 3129 -23808
rect 3065 -23952 3129 -23888
rect 3065 -24032 3129 -23968
rect 3065 -24112 3129 -24048
rect 3065 -24192 3129 -24128
rect 3065 -24272 3129 -24208
rect 3065 -24352 3129 -24288
rect 3065 -24432 3129 -24368
rect 3065 -24512 3129 -24448
rect 3065 -24592 3129 -24528
rect 3065 -24672 3129 -24608
rect 3065 -24752 3129 -24688
rect 3065 -24832 3129 -24768
rect 3065 -24912 3129 -24848
rect 3065 -24992 3129 -24928
rect 3065 -25072 3129 -25008
rect 3065 -25152 3129 -25088
rect 3065 -25232 3129 -25168
rect 3065 -25312 3129 -25248
rect 3065 -25392 3129 -25328
rect 3065 -25472 3129 -25408
rect 3065 -25552 3129 -25488
rect 3065 -25632 3129 -25568
rect 3065 -25712 3129 -25648
rect 3065 -25792 3129 -25728
rect 3065 -25872 3129 -25808
rect 3065 -25952 3129 -25888
rect 3065 -26032 3129 -25968
rect 3065 -26112 3129 -26048
rect 3065 -26192 3129 -26128
rect 3065 -26272 3129 -26208
rect 3065 -26352 3129 -26288
rect 3065 -26432 3129 -26368
rect 3065 -26512 3129 -26448
rect 3065 -26592 3129 -26528
rect 3065 -26672 3129 -26608
rect 3065 -26752 3129 -26688
rect 3065 -26832 3129 -26768
rect 3065 -26912 3129 -26848
rect 3065 -26992 3129 -26928
rect 3065 -27072 3129 -27008
rect 3065 -27152 3129 -27088
rect 3065 -27232 3129 -27168
rect 3065 -27312 3129 -27248
rect 3065 -27392 3129 -27328
rect 3065 -27472 3129 -27408
rect 3065 -27552 3129 -27488
rect 3065 -27632 3129 -27568
rect 3065 -27712 3129 -27648
rect 3065 -27792 3129 -27728
rect 3065 -27872 3129 -27808
rect 3065 -27952 3129 -27888
rect 3065 -28032 3129 -27968
rect 3065 -28112 3129 -28048
rect 3065 -28192 3129 -28128
rect 3065 -28272 3129 -28208
rect 9384 -22192 9448 -22128
rect 9384 -22272 9448 -22208
rect 9384 -22352 9448 -22288
rect 9384 -22432 9448 -22368
rect 9384 -22512 9448 -22448
rect 9384 -22592 9448 -22528
rect 9384 -22672 9448 -22608
rect 9384 -22752 9448 -22688
rect 9384 -22832 9448 -22768
rect 9384 -22912 9448 -22848
rect 9384 -22992 9448 -22928
rect 9384 -23072 9448 -23008
rect 9384 -23152 9448 -23088
rect 9384 -23232 9448 -23168
rect 9384 -23312 9448 -23248
rect 9384 -23392 9448 -23328
rect 9384 -23472 9448 -23408
rect 9384 -23552 9448 -23488
rect 9384 -23632 9448 -23568
rect 9384 -23712 9448 -23648
rect 9384 -23792 9448 -23728
rect 9384 -23872 9448 -23808
rect 9384 -23952 9448 -23888
rect 9384 -24032 9448 -23968
rect 9384 -24112 9448 -24048
rect 9384 -24192 9448 -24128
rect 9384 -24272 9448 -24208
rect 9384 -24352 9448 -24288
rect 9384 -24432 9448 -24368
rect 9384 -24512 9448 -24448
rect 9384 -24592 9448 -24528
rect 9384 -24672 9448 -24608
rect 9384 -24752 9448 -24688
rect 9384 -24832 9448 -24768
rect 9384 -24912 9448 -24848
rect 9384 -24992 9448 -24928
rect 9384 -25072 9448 -25008
rect 9384 -25152 9448 -25088
rect 9384 -25232 9448 -25168
rect 9384 -25312 9448 -25248
rect 9384 -25392 9448 -25328
rect 9384 -25472 9448 -25408
rect 9384 -25552 9448 -25488
rect 9384 -25632 9448 -25568
rect 9384 -25712 9448 -25648
rect 9384 -25792 9448 -25728
rect 9384 -25872 9448 -25808
rect 9384 -25952 9448 -25888
rect 9384 -26032 9448 -25968
rect 9384 -26112 9448 -26048
rect 9384 -26192 9448 -26128
rect 9384 -26272 9448 -26208
rect 9384 -26352 9448 -26288
rect 9384 -26432 9448 -26368
rect 9384 -26512 9448 -26448
rect 9384 -26592 9448 -26528
rect 9384 -26672 9448 -26608
rect 9384 -26752 9448 -26688
rect 9384 -26832 9448 -26768
rect 9384 -26912 9448 -26848
rect 9384 -26992 9448 -26928
rect 9384 -27072 9448 -27008
rect 9384 -27152 9448 -27088
rect 9384 -27232 9448 -27168
rect 9384 -27312 9448 -27248
rect 9384 -27392 9448 -27328
rect 9384 -27472 9448 -27408
rect 9384 -27552 9448 -27488
rect 9384 -27632 9448 -27568
rect 9384 -27712 9448 -27648
rect 9384 -27792 9448 -27728
rect 9384 -27872 9448 -27808
rect 9384 -27952 9448 -27888
rect 9384 -28032 9448 -27968
rect 9384 -28112 9448 -28048
rect 9384 -28192 9448 -28128
rect 9384 -28272 9448 -28208
rect 15703 -22192 15767 -22128
rect 15703 -22272 15767 -22208
rect 15703 -22352 15767 -22288
rect 15703 -22432 15767 -22368
rect 15703 -22512 15767 -22448
rect 15703 -22592 15767 -22528
rect 15703 -22672 15767 -22608
rect 15703 -22752 15767 -22688
rect 15703 -22832 15767 -22768
rect 15703 -22912 15767 -22848
rect 15703 -22992 15767 -22928
rect 15703 -23072 15767 -23008
rect 15703 -23152 15767 -23088
rect 15703 -23232 15767 -23168
rect 15703 -23312 15767 -23248
rect 15703 -23392 15767 -23328
rect 15703 -23472 15767 -23408
rect 15703 -23552 15767 -23488
rect 15703 -23632 15767 -23568
rect 15703 -23712 15767 -23648
rect 15703 -23792 15767 -23728
rect 15703 -23872 15767 -23808
rect 15703 -23952 15767 -23888
rect 15703 -24032 15767 -23968
rect 15703 -24112 15767 -24048
rect 15703 -24192 15767 -24128
rect 15703 -24272 15767 -24208
rect 15703 -24352 15767 -24288
rect 15703 -24432 15767 -24368
rect 15703 -24512 15767 -24448
rect 15703 -24592 15767 -24528
rect 15703 -24672 15767 -24608
rect 15703 -24752 15767 -24688
rect 15703 -24832 15767 -24768
rect 15703 -24912 15767 -24848
rect 15703 -24992 15767 -24928
rect 15703 -25072 15767 -25008
rect 15703 -25152 15767 -25088
rect 15703 -25232 15767 -25168
rect 15703 -25312 15767 -25248
rect 15703 -25392 15767 -25328
rect 15703 -25472 15767 -25408
rect 15703 -25552 15767 -25488
rect 15703 -25632 15767 -25568
rect 15703 -25712 15767 -25648
rect 15703 -25792 15767 -25728
rect 15703 -25872 15767 -25808
rect 15703 -25952 15767 -25888
rect 15703 -26032 15767 -25968
rect 15703 -26112 15767 -26048
rect 15703 -26192 15767 -26128
rect 15703 -26272 15767 -26208
rect 15703 -26352 15767 -26288
rect 15703 -26432 15767 -26368
rect 15703 -26512 15767 -26448
rect 15703 -26592 15767 -26528
rect 15703 -26672 15767 -26608
rect 15703 -26752 15767 -26688
rect 15703 -26832 15767 -26768
rect 15703 -26912 15767 -26848
rect 15703 -26992 15767 -26928
rect 15703 -27072 15767 -27008
rect 15703 -27152 15767 -27088
rect 15703 -27232 15767 -27168
rect 15703 -27312 15767 -27248
rect 15703 -27392 15767 -27328
rect 15703 -27472 15767 -27408
rect 15703 -27552 15767 -27488
rect 15703 -27632 15767 -27568
rect 15703 -27712 15767 -27648
rect 15703 -27792 15767 -27728
rect 15703 -27872 15767 -27808
rect 15703 -27952 15767 -27888
rect 15703 -28032 15767 -27968
rect 15703 -28112 15767 -28048
rect 15703 -28192 15767 -28128
rect 15703 -28272 15767 -28208
rect 22022 -22192 22086 -22128
rect 22022 -22272 22086 -22208
rect 22022 -22352 22086 -22288
rect 22022 -22432 22086 -22368
rect 22022 -22512 22086 -22448
rect 22022 -22592 22086 -22528
rect 22022 -22672 22086 -22608
rect 22022 -22752 22086 -22688
rect 22022 -22832 22086 -22768
rect 22022 -22912 22086 -22848
rect 22022 -22992 22086 -22928
rect 22022 -23072 22086 -23008
rect 22022 -23152 22086 -23088
rect 22022 -23232 22086 -23168
rect 22022 -23312 22086 -23248
rect 22022 -23392 22086 -23328
rect 22022 -23472 22086 -23408
rect 22022 -23552 22086 -23488
rect 22022 -23632 22086 -23568
rect 22022 -23712 22086 -23648
rect 22022 -23792 22086 -23728
rect 22022 -23872 22086 -23808
rect 22022 -23952 22086 -23888
rect 22022 -24032 22086 -23968
rect 22022 -24112 22086 -24048
rect 22022 -24192 22086 -24128
rect 22022 -24272 22086 -24208
rect 22022 -24352 22086 -24288
rect 22022 -24432 22086 -24368
rect 22022 -24512 22086 -24448
rect 22022 -24592 22086 -24528
rect 22022 -24672 22086 -24608
rect 22022 -24752 22086 -24688
rect 22022 -24832 22086 -24768
rect 22022 -24912 22086 -24848
rect 22022 -24992 22086 -24928
rect 22022 -25072 22086 -25008
rect 22022 -25152 22086 -25088
rect 22022 -25232 22086 -25168
rect 22022 -25312 22086 -25248
rect 22022 -25392 22086 -25328
rect 22022 -25472 22086 -25408
rect 22022 -25552 22086 -25488
rect 22022 -25632 22086 -25568
rect 22022 -25712 22086 -25648
rect 22022 -25792 22086 -25728
rect 22022 -25872 22086 -25808
rect 22022 -25952 22086 -25888
rect 22022 -26032 22086 -25968
rect 22022 -26112 22086 -26048
rect 22022 -26192 22086 -26128
rect 22022 -26272 22086 -26208
rect 22022 -26352 22086 -26288
rect 22022 -26432 22086 -26368
rect 22022 -26512 22086 -26448
rect 22022 -26592 22086 -26528
rect 22022 -26672 22086 -26608
rect 22022 -26752 22086 -26688
rect 22022 -26832 22086 -26768
rect 22022 -26912 22086 -26848
rect 22022 -26992 22086 -26928
rect 22022 -27072 22086 -27008
rect 22022 -27152 22086 -27088
rect 22022 -27232 22086 -27168
rect 22022 -27312 22086 -27248
rect 22022 -27392 22086 -27328
rect 22022 -27472 22086 -27408
rect 22022 -27552 22086 -27488
rect 22022 -27632 22086 -27568
rect 22022 -27712 22086 -27648
rect 22022 -27792 22086 -27728
rect 22022 -27872 22086 -27808
rect 22022 -27952 22086 -27888
rect 22022 -28032 22086 -27968
rect 22022 -28112 22086 -28048
rect 22022 -28192 22086 -28128
rect 22022 -28272 22086 -28208
rect 28341 -22192 28405 -22128
rect 28341 -22272 28405 -22208
rect 28341 -22352 28405 -22288
rect 28341 -22432 28405 -22368
rect 28341 -22512 28405 -22448
rect 28341 -22592 28405 -22528
rect 28341 -22672 28405 -22608
rect 28341 -22752 28405 -22688
rect 28341 -22832 28405 -22768
rect 28341 -22912 28405 -22848
rect 28341 -22992 28405 -22928
rect 28341 -23072 28405 -23008
rect 28341 -23152 28405 -23088
rect 28341 -23232 28405 -23168
rect 28341 -23312 28405 -23248
rect 28341 -23392 28405 -23328
rect 28341 -23472 28405 -23408
rect 28341 -23552 28405 -23488
rect 28341 -23632 28405 -23568
rect 28341 -23712 28405 -23648
rect 28341 -23792 28405 -23728
rect 28341 -23872 28405 -23808
rect 28341 -23952 28405 -23888
rect 28341 -24032 28405 -23968
rect 28341 -24112 28405 -24048
rect 28341 -24192 28405 -24128
rect 28341 -24272 28405 -24208
rect 28341 -24352 28405 -24288
rect 28341 -24432 28405 -24368
rect 28341 -24512 28405 -24448
rect 28341 -24592 28405 -24528
rect 28341 -24672 28405 -24608
rect 28341 -24752 28405 -24688
rect 28341 -24832 28405 -24768
rect 28341 -24912 28405 -24848
rect 28341 -24992 28405 -24928
rect 28341 -25072 28405 -25008
rect 28341 -25152 28405 -25088
rect 28341 -25232 28405 -25168
rect 28341 -25312 28405 -25248
rect 28341 -25392 28405 -25328
rect 28341 -25472 28405 -25408
rect 28341 -25552 28405 -25488
rect 28341 -25632 28405 -25568
rect 28341 -25712 28405 -25648
rect 28341 -25792 28405 -25728
rect 28341 -25872 28405 -25808
rect 28341 -25952 28405 -25888
rect 28341 -26032 28405 -25968
rect 28341 -26112 28405 -26048
rect 28341 -26192 28405 -26128
rect 28341 -26272 28405 -26208
rect 28341 -26352 28405 -26288
rect 28341 -26432 28405 -26368
rect 28341 -26512 28405 -26448
rect 28341 -26592 28405 -26528
rect 28341 -26672 28405 -26608
rect 28341 -26752 28405 -26688
rect 28341 -26832 28405 -26768
rect 28341 -26912 28405 -26848
rect 28341 -26992 28405 -26928
rect 28341 -27072 28405 -27008
rect 28341 -27152 28405 -27088
rect 28341 -27232 28405 -27168
rect 28341 -27312 28405 -27248
rect 28341 -27392 28405 -27328
rect 28341 -27472 28405 -27408
rect 28341 -27552 28405 -27488
rect 28341 -27632 28405 -27568
rect 28341 -27712 28405 -27648
rect 28341 -27792 28405 -27728
rect 28341 -27872 28405 -27808
rect 28341 -27952 28405 -27888
rect 28341 -28032 28405 -27968
rect 28341 -28112 28405 -28048
rect 28341 -28192 28405 -28128
rect 28341 -28272 28405 -28208
rect 34660 -22192 34724 -22128
rect 34660 -22272 34724 -22208
rect 34660 -22352 34724 -22288
rect 34660 -22432 34724 -22368
rect 34660 -22512 34724 -22448
rect 34660 -22592 34724 -22528
rect 34660 -22672 34724 -22608
rect 34660 -22752 34724 -22688
rect 34660 -22832 34724 -22768
rect 34660 -22912 34724 -22848
rect 34660 -22992 34724 -22928
rect 34660 -23072 34724 -23008
rect 34660 -23152 34724 -23088
rect 34660 -23232 34724 -23168
rect 34660 -23312 34724 -23248
rect 34660 -23392 34724 -23328
rect 34660 -23472 34724 -23408
rect 34660 -23552 34724 -23488
rect 34660 -23632 34724 -23568
rect 34660 -23712 34724 -23648
rect 34660 -23792 34724 -23728
rect 34660 -23872 34724 -23808
rect 34660 -23952 34724 -23888
rect 34660 -24032 34724 -23968
rect 34660 -24112 34724 -24048
rect 34660 -24192 34724 -24128
rect 34660 -24272 34724 -24208
rect 34660 -24352 34724 -24288
rect 34660 -24432 34724 -24368
rect 34660 -24512 34724 -24448
rect 34660 -24592 34724 -24528
rect 34660 -24672 34724 -24608
rect 34660 -24752 34724 -24688
rect 34660 -24832 34724 -24768
rect 34660 -24912 34724 -24848
rect 34660 -24992 34724 -24928
rect 34660 -25072 34724 -25008
rect 34660 -25152 34724 -25088
rect 34660 -25232 34724 -25168
rect 34660 -25312 34724 -25248
rect 34660 -25392 34724 -25328
rect 34660 -25472 34724 -25408
rect 34660 -25552 34724 -25488
rect 34660 -25632 34724 -25568
rect 34660 -25712 34724 -25648
rect 34660 -25792 34724 -25728
rect 34660 -25872 34724 -25808
rect 34660 -25952 34724 -25888
rect 34660 -26032 34724 -25968
rect 34660 -26112 34724 -26048
rect 34660 -26192 34724 -26128
rect 34660 -26272 34724 -26208
rect 34660 -26352 34724 -26288
rect 34660 -26432 34724 -26368
rect 34660 -26512 34724 -26448
rect 34660 -26592 34724 -26528
rect 34660 -26672 34724 -26608
rect 34660 -26752 34724 -26688
rect 34660 -26832 34724 -26768
rect 34660 -26912 34724 -26848
rect 34660 -26992 34724 -26928
rect 34660 -27072 34724 -27008
rect 34660 -27152 34724 -27088
rect 34660 -27232 34724 -27168
rect 34660 -27312 34724 -27248
rect 34660 -27392 34724 -27328
rect 34660 -27472 34724 -27408
rect 34660 -27552 34724 -27488
rect 34660 -27632 34724 -27568
rect 34660 -27712 34724 -27648
rect 34660 -27792 34724 -27728
rect 34660 -27872 34724 -27808
rect 34660 -27952 34724 -27888
rect 34660 -28032 34724 -27968
rect 34660 -28112 34724 -28048
rect 34660 -28192 34724 -28128
rect 34660 -28272 34724 -28208
rect 40979 -22192 41043 -22128
rect 40979 -22272 41043 -22208
rect 40979 -22352 41043 -22288
rect 40979 -22432 41043 -22368
rect 40979 -22512 41043 -22448
rect 40979 -22592 41043 -22528
rect 40979 -22672 41043 -22608
rect 40979 -22752 41043 -22688
rect 40979 -22832 41043 -22768
rect 40979 -22912 41043 -22848
rect 40979 -22992 41043 -22928
rect 40979 -23072 41043 -23008
rect 40979 -23152 41043 -23088
rect 40979 -23232 41043 -23168
rect 40979 -23312 41043 -23248
rect 40979 -23392 41043 -23328
rect 40979 -23472 41043 -23408
rect 40979 -23552 41043 -23488
rect 40979 -23632 41043 -23568
rect 40979 -23712 41043 -23648
rect 40979 -23792 41043 -23728
rect 40979 -23872 41043 -23808
rect 40979 -23952 41043 -23888
rect 40979 -24032 41043 -23968
rect 40979 -24112 41043 -24048
rect 40979 -24192 41043 -24128
rect 40979 -24272 41043 -24208
rect 40979 -24352 41043 -24288
rect 40979 -24432 41043 -24368
rect 40979 -24512 41043 -24448
rect 40979 -24592 41043 -24528
rect 40979 -24672 41043 -24608
rect 40979 -24752 41043 -24688
rect 40979 -24832 41043 -24768
rect 40979 -24912 41043 -24848
rect 40979 -24992 41043 -24928
rect 40979 -25072 41043 -25008
rect 40979 -25152 41043 -25088
rect 40979 -25232 41043 -25168
rect 40979 -25312 41043 -25248
rect 40979 -25392 41043 -25328
rect 40979 -25472 41043 -25408
rect 40979 -25552 41043 -25488
rect 40979 -25632 41043 -25568
rect 40979 -25712 41043 -25648
rect 40979 -25792 41043 -25728
rect 40979 -25872 41043 -25808
rect 40979 -25952 41043 -25888
rect 40979 -26032 41043 -25968
rect 40979 -26112 41043 -26048
rect 40979 -26192 41043 -26128
rect 40979 -26272 41043 -26208
rect 40979 -26352 41043 -26288
rect 40979 -26432 41043 -26368
rect 40979 -26512 41043 -26448
rect 40979 -26592 41043 -26528
rect 40979 -26672 41043 -26608
rect 40979 -26752 41043 -26688
rect 40979 -26832 41043 -26768
rect 40979 -26912 41043 -26848
rect 40979 -26992 41043 -26928
rect 40979 -27072 41043 -27008
rect 40979 -27152 41043 -27088
rect 40979 -27232 41043 -27168
rect 40979 -27312 41043 -27248
rect 40979 -27392 41043 -27328
rect 40979 -27472 41043 -27408
rect 40979 -27552 41043 -27488
rect 40979 -27632 41043 -27568
rect 40979 -27712 41043 -27648
rect 40979 -27792 41043 -27728
rect 40979 -27872 41043 -27808
rect 40979 -27952 41043 -27888
rect 40979 -28032 41043 -27968
rect 40979 -28112 41043 -28048
rect 40979 -28192 41043 -28128
rect 40979 -28272 41043 -28208
rect 47298 -22192 47362 -22128
rect 47298 -22272 47362 -22208
rect 47298 -22352 47362 -22288
rect 47298 -22432 47362 -22368
rect 47298 -22512 47362 -22448
rect 47298 -22592 47362 -22528
rect 47298 -22672 47362 -22608
rect 47298 -22752 47362 -22688
rect 47298 -22832 47362 -22768
rect 47298 -22912 47362 -22848
rect 47298 -22992 47362 -22928
rect 47298 -23072 47362 -23008
rect 47298 -23152 47362 -23088
rect 47298 -23232 47362 -23168
rect 47298 -23312 47362 -23248
rect 47298 -23392 47362 -23328
rect 47298 -23472 47362 -23408
rect 47298 -23552 47362 -23488
rect 47298 -23632 47362 -23568
rect 47298 -23712 47362 -23648
rect 47298 -23792 47362 -23728
rect 47298 -23872 47362 -23808
rect 47298 -23952 47362 -23888
rect 47298 -24032 47362 -23968
rect 47298 -24112 47362 -24048
rect 47298 -24192 47362 -24128
rect 47298 -24272 47362 -24208
rect 47298 -24352 47362 -24288
rect 47298 -24432 47362 -24368
rect 47298 -24512 47362 -24448
rect 47298 -24592 47362 -24528
rect 47298 -24672 47362 -24608
rect 47298 -24752 47362 -24688
rect 47298 -24832 47362 -24768
rect 47298 -24912 47362 -24848
rect 47298 -24992 47362 -24928
rect 47298 -25072 47362 -25008
rect 47298 -25152 47362 -25088
rect 47298 -25232 47362 -25168
rect 47298 -25312 47362 -25248
rect 47298 -25392 47362 -25328
rect 47298 -25472 47362 -25408
rect 47298 -25552 47362 -25488
rect 47298 -25632 47362 -25568
rect 47298 -25712 47362 -25648
rect 47298 -25792 47362 -25728
rect 47298 -25872 47362 -25808
rect 47298 -25952 47362 -25888
rect 47298 -26032 47362 -25968
rect 47298 -26112 47362 -26048
rect 47298 -26192 47362 -26128
rect 47298 -26272 47362 -26208
rect 47298 -26352 47362 -26288
rect 47298 -26432 47362 -26368
rect 47298 -26512 47362 -26448
rect 47298 -26592 47362 -26528
rect 47298 -26672 47362 -26608
rect 47298 -26752 47362 -26688
rect 47298 -26832 47362 -26768
rect 47298 -26912 47362 -26848
rect 47298 -26992 47362 -26928
rect 47298 -27072 47362 -27008
rect 47298 -27152 47362 -27088
rect 47298 -27232 47362 -27168
rect 47298 -27312 47362 -27248
rect 47298 -27392 47362 -27328
rect 47298 -27472 47362 -27408
rect 47298 -27552 47362 -27488
rect 47298 -27632 47362 -27568
rect 47298 -27712 47362 -27648
rect 47298 -27792 47362 -27728
rect 47298 -27872 47362 -27808
rect 47298 -27952 47362 -27888
rect 47298 -28032 47362 -27968
rect 47298 -28112 47362 -28048
rect 47298 -28192 47362 -28128
rect 47298 -28272 47362 -28208
rect -41168 -28492 -41104 -28428
rect -41168 -28572 -41104 -28508
rect -41168 -28652 -41104 -28588
rect -41168 -28732 -41104 -28668
rect -41168 -28812 -41104 -28748
rect -41168 -28892 -41104 -28828
rect -41168 -28972 -41104 -28908
rect -41168 -29052 -41104 -28988
rect -41168 -29132 -41104 -29068
rect -41168 -29212 -41104 -29148
rect -41168 -29292 -41104 -29228
rect -41168 -29372 -41104 -29308
rect -41168 -29452 -41104 -29388
rect -41168 -29532 -41104 -29468
rect -41168 -29612 -41104 -29548
rect -41168 -29692 -41104 -29628
rect -41168 -29772 -41104 -29708
rect -41168 -29852 -41104 -29788
rect -41168 -29932 -41104 -29868
rect -41168 -30012 -41104 -29948
rect -41168 -30092 -41104 -30028
rect -41168 -30172 -41104 -30108
rect -41168 -30252 -41104 -30188
rect -41168 -30332 -41104 -30268
rect -41168 -30412 -41104 -30348
rect -41168 -30492 -41104 -30428
rect -41168 -30572 -41104 -30508
rect -41168 -30652 -41104 -30588
rect -41168 -30732 -41104 -30668
rect -41168 -30812 -41104 -30748
rect -41168 -30892 -41104 -30828
rect -41168 -30972 -41104 -30908
rect -41168 -31052 -41104 -30988
rect -41168 -31132 -41104 -31068
rect -41168 -31212 -41104 -31148
rect -41168 -31292 -41104 -31228
rect -41168 -31372 -41104 -31308
rect -41168 -31452 -41104 -31388
rect -41168 -31532 -41104 -31468
rect -41168 -31612 -41104 -31548
rect -41168 -31692 -41104 -31628
rect -41168 -31772 -41104 -31708
rect -41168 -31852 -41104 -31788
rect -41168 -31932 -41104 -31868
rect -41168 -32012 -41104 -31948
rect -41168 -32092 -41104 -32028
rect -41168 -32172 -41104 -32108
rect -41168 -32252 -41104 -32188
rect -41168 -32332 -41104 -32268
rect -41168 -32412 -41104 -32348
rect -41168 -32492 -41104 -32428
rect -41168 -32572 -41104 -32508
rect -41168 -32652 -41104 -32588
rect -41168 -32732 -41104 -32668
rect -41168 -32812 -41104 -32748
rect -41168 -32892 -41104 -32828
rect -41168 -32972 -41104 -32908
rect -41168 -33052 -41104 -32988
rect -41168 -33132 -41104 -33068
rect -41168 -33212 -41104 -33148
rect -41168 -33292 -41104 -33228
rect -41168 -33372 -41104 -33308
rect -41168 -33452 -41104 -33388
rect -41168 -33532 -41104 -33468
rect -41168 -33612 -41104 -33548
rect -41168 -33692 -41104 -33628
rect -41168 -33772 -41104 -33708
rect -41168 -33852 -41104 -33788
rect -41168 -33932 -41104 -33868
rect -41168 -34012 -41104 -33948
rect -41168 -34092 -41104 -34028
rect -41168 -34172 -41104 -34108
rect -41168 -34252 -41104 -34188
rect -41168 -34332 -41104 -34268
rect -41168 -34412 -41104 -34348
rect -41168 -34492 -41104 -34428
rect -41168 -34572 -41104 -34508
rect -34849 -28492 -34785 -28428
rect -34849 -28572 -34785 -28508
rect -34849 -28652 -34785 -28588
rect -34849 -28732 -34785 -28668
rect -34849 -28812 -34785 -28748
rect -34849 -28892 -34785 -28828
rect -34849 -28972 -34785 -28908
rect -34849 -29052 -34785 -28988
rect -34849 -29132 -34785 -29068
rect -34849 -29212 -34785 -29148
rect -34849 -29292 -34785 -29228
rect -34849 -29372 -34785 -29308
rect -34849 -29452 -34785 -29388
rect -34849 -29532 -34785 -29468
rect -34849 -29612 -34785 -29548
rect -34849 -29692 -34785 -29628
rect -34849 -29772 -34785 -29708
rect -34849 -29852 -34785 -29788
rect -34849 -29932 -34785 -29868
rect -34849 -30012 -34785 -29948
rect -34849 -30092 -34785 -30028
rect -34849 -30172 -34785 -30108
rect -34849 -30252 -34785 -30188
rect -34849 -30332 -34785 -30268
rect -34849 -30412 -34785 -30348
rect -34849 -30492 -34785 -30428
rect -34849 -30572 -34785 -30508
rect -34849 -30652 -34785 -30588
rect -34849 -30732 -34785 -30668
rect -34849 -30812 -34785 -30748
rect -34849 -30892 -34785 -30828
rect -34849 -30972 -34785 -30908
rect -34849 -31052 -34785 -30988
rect -34849 -31132 -34785 -31068
rect -34849 -31212 -34785 -31148
rect -34849 -31292 -34785 -31228
rect -34849 -31372 -34785 -31308
rect -34849 -31452 -34785 -31388
rect -34849 -31532 -34785 -31468
rect -34849 -31612 -34785 -31548
rect -34849 -31692 -34785 -31628
rect -34849 -31772 -34785 -31708
rect -34849 -31852 -34785 -31788
rect -34849 -31932 -34785 -31868
rect -34849 -32012 -34785 -31948
rect -34849 -32092 -34785 -32028
rect -34849 -32172 -34785 -32108
rect -34849 -32252 -34785 -32188
rect -34849 -32332 -34785 -32268
rect -34849 -32412 -34785 -32348
rect -34849 -32492 -34785 -32428
rect -34849 -32572 -34785 -32508
rect -34849 -32652 -34785 -32588
rect -34849 -32732 -34785 -32668
rect -34849 -32812 -34785 -32748
rect -34849 -32892 -34785 -32828
rect -34849 -32972 -34785 -32908
rect -34849 -33052 -34785 -32988
rect -34849 -33132 -34785 -33068
rect -34849 -33212 -34785 -33148
rect -34849 -33292 -34785 -33228
rect -34849 -33372 -34785 -33308
rect -34849 -33452 -34785 -33388
rect -34849 -33532 -34785 -33468
rect -34849 -33612 -34785 -33548
rect -34849 -33692 -34785 -33628
rect -34849 -33772 -34785 -33708
rect -34849 -33852 -34785 -33788
rect -34849 -33932 -34785 -33868
rect -34849 -34012 -34785 -33948
rect -34849 -34092 -34785 -34028
rect -34849 -34172 -34785 -34108
rect -34849 -34252 -34785 -34188
rect -34849 -34332 -34785 -34268
rect -34849 -34412 -34785 -34348
rect -34849 -34492 -34785 -34428
rect -34849 -34572 -34785 -34508
rect -28530 -28492 -28466 -28428
rect -28530 -28572 -28466 -28508
rect -28530 -28652 -28466 -28588
rect -28530 -28732 -28466 -28668
rect -28530 -28812 -28466 -28748
rect -28530 -28892 -28466 -28828
rect -28530 -28972 -28466 -28908
rect -28530 -29052 -28466 -28988
rect -28530 -29132 -28466 -29068
rect -28530 -29212 -28466 -29148
rect -28530 -29292 -28466 -29228
rect -28530 -29372 -28466 -29308
rect -28530 -29452 -28466 -29388
rect -28530 -29532 -28466 -29468
rect -28530 -29612 -28466 -29548
rect -28530 -29692 -28466 -29628
rect -28530 -29772 -28466 -29708
rect -28530 -29852 -28466 -29788
rect -28530 -29932 -28466 -29868
rect -28530 -30012 -28466 -29948
rect -28530 -30092 -28466 -30028
rect -28530 -30172 -28466 -30108
rect -28530 -30252 -28466 -30188
rect -28530 -30332 -28466 -30268
rect -28530 -30412 -28466 -30348
rect -28530 -30492 -28466 -30428
rect -28530 -30572 -28466 -30508
rect -28530 -30652 -28466 -30588
rect -28530 -30732 -28466 -30668
rect -28530 -30812 -28466 -30748
rect -28530 -30892 -28466 -30828
rect -28530 -30972 -28466 -30908
rect -28530 -31052 -28466 -30988
rect -28530 -31132 -28466 -31068
rect -28530 -31212 -28466 -31148
rect -28530 -31292 -28466 -31228
rect -28530 -31372 -28466 -31308
rect -28530 -31452 -28466 -31388
rect -28530 -31532 -28466 -31468
rect -28530 -31612 -28466 -31548
rect -28530 -31692 -28466 -31628
rect -28530 -31772 -28466 -31708
rect -28530 -31852 -28466 -31788
rect -28530 -31932 -28466 -31868
rect -28530 -32012 -28466 -31948
rect -28530 -32092 -28466 -32028
rect -28530 -32172 -28466 -32108
rect -28530 -32252 -28466 -32188
rect -28530 -32332 -28466 -32268
rect -28530 -32412 -28466 -32348
rect -28530 -32492 -28466 -32428
rect -28530 -32572 -28466 -32508
rect -28530 -32652 -28466 -32588
rect -28530 -32732 -28466 -32668
rect -28530 -32812 -28466 -32748
rect -28530 -32892 -28466 -32828
rect -28530 -32972 -28466 -32908
rect -28530 -33052 -28466 -32988
rect -28530 -33132 -28466 -33068
rect -28530 -33212 -28466 -33148
rect -28530 -33292 -28466 -33228
rect -28530 -33372 -28466 -33308
rect -28530 -33452 -28466 -33388
rect -28530 -33532 -28466 -33468
rect -28530 -33612 -28466 -33548
rect -28530 -33692 -28466 -33628
rect -28530 -33772 -28466 -33708
rect -28530 -33852 -28466 -33788
rect -28530 -33932 -28466 -33868
rect -28530 -34012 -28466 -33948
rect -28530 -34092 -28466 -34028
rect -28530 -34172 -28466 -34108
rect -28530 -34252 -28466 -34188
rect -28530 -34332 -28466 -34268
rect -28530 -34412 -28466 -34348
rect -28530 -34492 -28466 -34428
rect -28530 -34572 -28466 -34508
rect -22211 -28492 -22147 -28428
rect -22211 -28572 -22147 -28508
rect -22211 -28652 -22147 -28588
rect -22211 -28732 -22147 -28668
rect -22211 -28812 -22147 -28748
rect -22211 -28892 -22147 -28828
rect -22211 -28972 -22147 -28908
rect -22211 -29052 -22147 -28988
rect -22211 -29132 -22147 -29068
rect -22211 -29212 -22147 -29148
rect -22211 -29292 -22147 -29228
rect -22211 -29372 -22147 -29308
rect -22211 -29452 -22147 -29388
rect -22211 -29532 -22147 -29468
rect -22211 -29612 -22147 -29548
rect -22211 -29692 -22147 -29628
rect -22211 -29772 -22147 -29708
rect -22211 -29852 -22147 -29788
rect -22211 -29932 -22147 -29868
rect -22211 -30012 -22147 -29948
rect -22211 -30092 -22147 -30028
rect -22211 -30172 -22147 -30108
rect -22211 -30252 -22147 -30188
rect -22211 -30332 -22147 -30268
rect -22211 -30412 -22147 -30348
rect -22211 -30492 -22147 -30428
rect -22211 -30572 -22147 -30508
rect -22211 -30652 -22147 -30588
rect -22211 -30732 -22147 -30668
rect -22211 -30812 -22147 -30748
rect -22211 -30892 -22147 -30828
rect -22211 -30972 -22147 -30908
rect -22211 -31052 -22147 -30988
rect -22211 -31132 -22147 -31068
rect -22211 -31212 -22147 -31148
rect -22211 -31292 -22147 -31228
rect -22211 -31372 -22147 -31308
rect -22211 -31452 -22147 -31388
rect -22211 -31532 -22147 -31468
rect -22211 -31612 -22147 -31548
rect -22211 -31692 -22147 -31628
rect -22211 -31772 -22147 -31708
rect -22211 -31852 -22147 -31788
rect -22211 -31932 -22147 -31868
rect -22211 -32012 -22147 -31948
rect -22211 -32092 -22147 -32028
rect -22211 -32172 -22147 -32108
rect -22211 -32252 -22147 -32188
rect -22211 -32332 -22147 -32268
rect -22211 -32412 -22147 -32348
rect -22211 -32492 -22147 -32428
rect -22211 -32572 -22147 -32508
rect -22211 -32652 -22147 -32588
rect -22211 -32732 -22147 -32668
rect -22211 -32812 -22147 -32748
rect -22211 -32892 -22147 -32828
rect -22211 -32972 -22147 -32908
rect -22211 -33052 -22147 -32988
rect -22211 -33132 -22147 -33068
rect -22211 -33212 -22147 -33148
rect -22211 -33292 -22147 -33228
rect -22211 -33372 -22147 -33308
rect -22211 -33452 -22147 -33388
rect -22211 -33532 -22147 -33468
rect -22211 -33612 -22147 -33548
rect -22211 -33692 -22147 -33628
rect -22211 -33772 -22147 -33708
rect -22211 -33852 -22147 -33788
rect -22211 -33932 -22147 -33868
rect -22211 -34012 -22147 -33948
rect -22211 -34092 -22147 -34028
rect -22211 -34172 -22147 -34108
rect -22211 -34252 -22147 -34188
rect -22211 -34332 -22147 -34268
rect -22211 -34412 -22147 -34348
rect -22211 -34492 -22147 -34428
rect -22211 -34572 -22147 -34508
rect -15892 -28492 -15828 -28428
rect -15892 -28572 -15828 -28508
rect -15892 -28652 -15828 -28588
rect -15892 -28732 -15828 -28668
rect -15892 -28812 -15828 -28748
rect -15892 -28892 -15828 -28828
rect -15892 -28972 -15828 -28908
rect -15892 -29052 -15828 -28988
rect -15892 -29132 -15828 -29068
rect -15892 -29212 -15828 -29148
rect -15892 -29292 -15828 -29228
rect -15892 -29372 -15828 -29308
rect -15892 -29452 -15828 -29388
rect -15892 -29532 -15828 -29468
rect -15892 -29612 -15828 -29548
rect -15892 -29692 -15828 -29628
rect -15892 -29772 -15828 -29708
rect -15892 -29852 -15828 -29788
rect -15892 -29932 -15828 -29868
rect -15892 -30012 -15828 -29948
rect -15892 -30092 -15828 -30028
rect -15892 -30172 -15828 -30108
rect -15892 -30252 -15828 -30188
rect -15892 -30332 -15828 -30268
rect -15892 -30412 -15828 -30348
rect -15892 -30492 -15828 -30428
rect -15892 -30572 -15828 -30508
rect -15892 -30652 -15828 -30588
rect -15892 -30732 -15828 -30668
rect -15892 -30812 -15828 -30748
rect -15892 -30892 -15828 -30828
rect -15892 -30972 -15828 -30908
rect -15892 -31052 -15828 -30988
rect -15892 -31132 -15828 -31068
rect -15892 -31212 -15828 -31148
rect -15892 -31292 -15828 -31228
rect -15892 -31372 -15828 -31308
rect -15892 -31452 -15828 -31388
rect -15892 -31532 -15828 -31468
rect -15892 -31612 -15828 -31548
rect -15892 -31692 -15828 -31628
rect -15892 -31772 -15828 -31708
rect -15892 -31852 -15828 -31788
rect -15892 -31932 -15828 -31868
rect -15892 -32012 -15828 -31948
rect -15892 -32092 -15828 -32028
rect -15892 -32172 -15828 -32108
rect -15892 -32252 -15828 -32188
rect -15892 -32332 -15828 -32268
rect -15892 -32412 -15828 -32348
rect -15892 -32492 -15828 -32428
rect -15892 -32572 -15828 -32508
rect -15892 -32652 -15828 -32588
rect -15892 -32732 -15828 -32668
rect -15892 -32812 -15828 -32748
rect -15892 -32892 -15828 -32828
rect -15892 -32972 -15828 -32908
rect -15892 -33052 -15828 -32988
rect -15892 -33132 -15828 -33068
rect -15892 -33212 -15828 -33148
rect -15892 -33292 -15828 -33228
rect -15892 -33372 -15828 -33308
rect -15892 -33452 -15828 -33388
rect -15892 -33532 -15828 -33468
rect -15892 -33612 -15828 -33548
rect -15892 -33692 -15828 -33628
rect -15892 -33772 -15828 -33708
rect -15892 -33852 -15828 -33788
rect -15892 -33932 -15828 -33868
rect -15892 -34012 -15828 -33948
rect -15892 -34092 -15828 -34028
rect -15892 -34172 -15828 -34108
rect -15892 -34252 -15828 -34188
rect -15892 -34332 -15828 -34268
rect -15892 -34412 -15828 -34348
rect -15892 -34492 -15828 -34428
rect -15892 -34572 -15828 -34508
rect -9573 -28492 -9509 -28428
rect -9573 -28572 -9509 -28508
rect -9573 -28652 -9509 -28588
rect -9573 -28732 -9509 -28668
rect -9573 -28812 -9509 -28748
rect -9573 -28892 -9509 -28828
rect -9573 -28972 -9509 -28908
rect -9573 -29052 -9509 -28988
rect -9573 -29132 -9509 -29068
rect -9573 -29212 -9509 -29148
rect -9573 -29292 -9509 -29228
rect -9573 -29372 -9509 -29308
rect -9573 -29452 -9509 -29388
rect -9573 -29532 -9509 -29468
rect -9573 -29612 -9509 -29548
rect -9573 -29692 -9509 -29628
rect -9573 -29772 -9509 -29708
rect -9573 -29852 -9509 -29788
rect -9573 -29932 -9509 -29868
rect -9573 -30012 -9509 -29948
rect -9573 -30092 -9509 -30028
rect -9573 -30172 -9509 -30108
rect -9573 -30252 -9509 -30188
rect -9573 -30332 -9509 -30268
rect -9573 -30412 -9509 -30348
rect -9573 -30492 -9509 -30428
rect -9573 -30572 -9509 -30508
rect -9573 -30652 -9509 -30588
rect -9573 -30732 -9509 -30668
rect -9573 -30812 -9509 -30748
rect -9573 -30892 -9509 -30828
rect -9573 -30972 -9509 -30908
rect -9573 -31052 -9509 -30988
rect -9573 -31132 -9509 -31068
rect -9573 -31212 -9509 -31148
rect -9573 -31292 -9509 -31228
rect -9573 -31372 -9509 -31308
rect -9573 -31452 -9509 -31388
rect -9573 -31532 -9509 -31468
rect -9573 -31612 -9509 -31548
rect -9573 -31692 -9509 -31628
rect -9573 -31772 -9509 -31708
rect -9573 -31852 -9509 -31788
rect -9573 -31932 -9509 -31868
rect -9573 -32012 -9509 -31948
rect -9573 -32092 -9509 -32028
rect -9573 -32172 -9509 -32108
rect -9573 -32252 -9509 -32188
rect -9573 -32332 -9509 -32268
rect -9573 -32412 -9509 -32348
rect -9573 -32492 -9509 -32428
rect -9573 -32572 -9509 -32508
rect -9573 -32652 -9509 -32588
rect -9573 -32732 -9509 -32668
rect -9573 -32812 -9509 -32748
rect -9573 -32892 -9509 -32828
rect -9573 -32972 -9509 -32908
rect -9573 -33052 -9509 -32988
rect -9573 -33132 -9509 -33068
rect -9573 -33212 -9509 -33148
rect -9573 -33292 -9509 -33228
rect -9573 -33372 -9509 -33308
rect -9573 -33452 -9509 -33388
rect -9573 -33532 -9509 -33468
rect -9573 -33612 -9509 -33548
rect -9573 -33692 -9509 -33628
rect -9573 -33772 -9509 -33708
rect -9573 -33852 -9509 -33788
rect -9573 -33932 -9509 -33868
rect -9573 -34012 -9509 -33948
rect -9573 -34092 -9509 -34028
rect -9573 -34172 -9509 -34108
rect -9573 -34252 -9509 -34188
rect -9573 -34332 -9509 -34268
rect -9573 -34412 -9509 -34348
rect -9573 -34492 -9509 -34428
rect -9573 -34572 -9509 -34508
rect -3254 -28492 -3190 -28428
rect -3254 -28572 -3190 -28508
rect -3254 -28652 -3190 -28588
rect -3254 -28732 -3190 -28668
rect -3254 -28812 -3190 -28748
rect -3254 -28892 -3190 -28828
rect -3254 -28972 -3190 -28908
rect -3254 -29052 -3190 -28988
rect -3254 -29132 -3190 -29068
rect -3254 -29212 -3190 -29148
rect -3254 -29292 -3190 -29228
rect -3254 -29372 -3190 -29308
rect -3254 -29452 -3190 -29388
rect -3254 -29532 -3190 -29468
rect -3254 -29612 -3190 -29548
rect -3254 -29692 -3190 -29628
rect -3254 -29772 -3190 -29708
rect -3254 -29852 -3190 -29788
rect -3254 -29932 -3190 -29868
rect -3254 -30012 -3190 -29948
rect -3254 -30092 -3190 -30028
rect -3254 -30172 -3190 -30108
rect -3254 -30252 -3190 -30188
rect -3254 -30332 -3190 -30268
rect -3254 -30412 -3190 -30348
rect -3254 -30492 -3190 -30428
rect -3254 -30572 -3190 -30508
rect -3254 -30652 -3190 -30588
rect -3254 -30732 -3190 -30668
rect -3254 -30812 -3190 -30748
rect -3254 -30892 -3190 -30828
rect -3254 -30972 -3190 -30908
rect -3254 -31052 -3190 -30988
rect -3254 -31132 -3190 -31068
rect -3254 -31212 -3190 -31148
rect -3254 -31292 -3190 -31228
rect -3254 -31372 -3190 -31308
rect -3254 -31452 -3190 -31388
rect -3254 -31532 -3190 -31468
rect -3254 -31612 -3190 -31548
rect -3254 -31692 -3190 -31628
rect -3254 -31772 -3190 -31708
rect -3254 -31852 -3190 -31788
rect -3254 -31932 -3190 -31868
rect -3254 -32012 -3190 -31948
rect -3254 -32092 -3190 -32028
rect -3254 -32172 -3190 -32108
rect -3254 -32252 -3190 -32188
rect -3254 -32332 -3190 -32268
rect -3254 -32412 -3190 -32348
rect -3254 -32492 -3190 -32428
rect -3254 -32572 -3190 -32508
rect -3254 -32652 -3190 -32588
rect -3254 -32732 -3190 -32668
rect -3254 -32812 -3190 -32748
rect -3254 -32892 -3190 -32828
rect -3254 -32972 -3190 -32908
rect -3254 -33052 -3190 -32988
rect -3254 -33132 -3190 -33068
rect -3254 -33212 -3190 -33148
rect -3254 -33292 -3190 -33228
rect -3254 -33372 -3190 -33308
rect -3254 -33452 -3190 -33388
rect -3254 -33532 -3190 -33468
rect -3254 -33612 -3190 -33548
rect -3254 -33692 -3190 -33628
rect -3254 -33772 -3190 -33708
rect -3254 -33852 -3190 -33788
rect -3254 -33932 -3190 -33868
rect -3254 -34012 -3190 -33948
rect -3254 -34092 -3190 -34028
rect -3254 -34172 -3190 -34108
rect -3254 -34252 -3190 -34188
rect -3254 -34332 -3190 -34268
rect -3254 -34412 -3190 -34348
rect -3254 -34492 -3190 -34428
rect -3254 -34572 -3190 -34508
rect 3065 -28492 3129 -28428
rect 3065 -28572 3129 -28508
rect 3065 -28652 3129 -28588
rect 3065 -28732 3129 -28668
rect 3065 -28812 3129 -28748
rect 3065 -28892 3129 -28828
rect 3065 -28972 3129 -28908
rect 3065 -29052 3129 -28988
rect 3065 -29132 3129 -29068
rect 3065 -29212 3129 -29148
rect 3065 -29292 3129 -29228
rect 3065 -29372 3129 -29308
rect 3065 -29452 3129 -29388
rect 3065 -29532 3129 -29468
rect 3065 -29612 3129 -29548
rect 3065 -29692 3129 -29628
rect 3065 -29772 3129 -29708
rect 3065 -29852 3129 -29788
rect 3065 -29932 3129 -29868
rect 3065 -30012 3129 -29948
rect 3065 -30092 3129 -30028
rect 3065 -30172 3129 -30108
rect 3065 -30252 3129 -30188
rect 3065 -30332 3129 -30268
rect 3065 -30412 3129 -30348
rect 3065 -30492 3129 -30428
rect 3065 -30572 3129 -30508
rect 3065 -30652 3129 -30588
rect 3065 -30732 3129 -30668
rect 3065 -30812 3129 -30748
rect 3065 -30892 3129 -30828
rect 3065 -30972 3129 -30908
rect 3065 -31052 3129 -30988
rect 3065 -31132 3129 -31068
rect 3065 -31212 3129 -31148
rect 3065 -31292 3129 -31228
rect 3065 -31372 3129 -31308
rect 3065 -31452 3129 -31388
rect 3065 -31532 3129 -31468
rect 3065 -31612 3129 -31548
rect 3065 -31692 3129 -31628
rect 3065 -31772 3129 -31708
rect 3065 -31852 3129 -31788
rect 3065 -31932 3129 -31868
rect 3065 -32012 3129 -31948
rect 3065 -32092 3129 -32028
rect 3065 -32172 3129 -32108
rect 3065 -32252 3129 -32188
rect 3065 -32332 3129 -32268
rect 3065 -32412 3129 -32348
rect 3065 -32492 3129 -32428
rect 3065 -32572 3129 -32508
rect 3065 -32652 3129 -32588
rect 3065 -32732 3129 -32668
rect 3065 -32812 3129 -32748
rect 3065 -32892 3129 -32828
rect 3065 -32972 3129 -32908
rect 3065 -33052 3129 -32988
rect 3065 -33132 3129 -33068
rect 3065 -33212 3129 -33148
rect 3065 -33292 3129 -33228
rect 3065 -33372 3129 -33308
rect 3065 -33452 3129 -33388
rect 3065 -33532 3129 -33468
rect 3065 -33612 3129 -33548
rect 3065 -33692 3129 -33628
rect 3065 -33772 3129 -33708
rect 3065 -33852 3129 -33788
rect 3065 -33932 3129 -33868
rect 3065 -34012 3129 -33948
rect 3065 -34092 3129 -34028
rect 3065 -34172 3129 -34108
rect 3065 -34252 3129 -34188
rect 3065 -34332 3129 -34268
rect 3065 -34412 3129 -34348
rect 3065 -34492 3129 -34428
rect 3065 -34572 3129 -34508
rect 9384 -28492 9448 -28428
rect 9384 -28572 9448 -28508
rect 9384 -28652 9448 -28588
rect 9384 -28732 9448 -28668
rect 9384 -28812 9448 -28748
rect 9384 -28892 9448 -28828
rect 9384 -28972 9448 -28908
rect 9384 -29052 9448 -28988
rect 9384 -29132 9448 -29068
rect 9384 -29212 9448 -29148
rect 9384 -29292 9448 -29228
rect 9384 -29372 9448 -29308
rect 9384 -29452 9448 -29388
rect 9384 -29532 9448 -29468
rect 9384 -29612 9448 -29548
rect 9384 -29692 9448 -29628
rect 9384 -29772 9448 -29708
rect 9384 -29852 9448 -29788
rect 9384 -29932 9448 -29868
rect 9384 -30012 9448 -29948
rect 9384 -30092 9448 -30028
rect 9384 -30172 9448 -30108
rect 9384 -30252 9448 -30188
rect 9384 -30332 9448 -30268
rect 9384 -30412 9448 -30348
rect 9384 -30492 9448 -30428
rect 9384 -30572 9448 -30508
rect 9384 -30652 9448 -30588
rect 9384 -30732 9448 -30668
rect 9384 -30812 9448 -30748
rect 9384 -30892 9448 -30828
rect 9384 -30972 9448 -30908
rect 9384 -31052 9448 -30988
rect 9384 -31132 9448 -31068
rect 9384 -31212 9448 -31148
rect 9384 -31292 9448 -31228
rect 9384 -31372 9448 -31308
rect 9384 -31452 9448 -31388
rect 9384 -31532 9448 -31468
rect 9384 -31612 9448 -31548
rect 9384 -31692 9448 -31628
rect 9384 -31772 9448 -31708
rect 9384 -31852 9448 -31788
rect 9384 -31932 9448 -31868
rect 9384 -32012 9448 -31948
rect 9384 -32092 9448 -32028
rect 9384 -32172 9448 -32108
rect 9384 -32252 9448 -32188
rect 9384 -32332 9448 -32268
rect 9384 -32412 9448 -32348
rect 9384 -32492 9448 -32428
rect 9384 -32572 9448 -32508
rect 9384 -32652 9448 -32588
rect 9384 -32732 9448 -32668
rect 9384 -32812 9448 -32748
rect 9384 -32892 9448 -32828
rect 9384 -32972 9448 -32908
rect 9384 -33052 9448 -32988
rect 9384 -33132 9448 -33068
rect 9384 -33212 9448 -33148
rect 9384 -33292 9448 -33228
rect 9384 -33372 9448 -33308
rect 9384 -33452 9448 -33388
rect 9384 -33532 9448 -33468
rect 9384 -33612 9448 -33548
rect 9384 -33692 9448 -33628
rect 9384 -33772 9448 -33708
rect 9384 -33852 9448 -33788
rect 9384 -33932 9448 -33868
rect 9384 -34012 9448 -33948
rect 9384 -34092 9448 -34028
rect 9384 -34172 9448 -34108
rect 9384 -34252 9448 -34188
rect 9384 -34332 9448 -34268
rect 9384 -34412 9448 -34348
rect 9384 -34492 9448 -34428
rect 9384 -34572 9448 -34508
rect 15703 -28492 15767 -28428
rect 15703 -28572 15767 -28508
rect 15703 -28652 15767 -28588
rect 15703 -28732 15767 -28668
rect 15703 -28812 15767 -28748
rect 15703 -28892 15767 -28828
rect 15703 -28972 15767 -28908
rect 15703 -29052 15767 -28988
rect 15703 -29132 15767 -29068
rect 15703 -29212 15767 -29148
rect 15703 -29292 15767 -29228
rect 15703 -29372 15767 -29308
rect 15703 -29452 15767 -29388
rect 15703 -29532 15767 -29468
rect 15703 -29612 15767 -29548
rect 15703 -29692 15767 -29628
rect 15703 -29772 15767 -29708
rect 15703 -29852 15767 -29788
rect 15703 -29932 15767 -29868
rect 15703 -30012 15767 -29948
rect 15703 -30092 15767 -30028
rect 15703 -30172 15767 -30108
rect 15703 -30252 15767 -30188
rect 15703 -30332 15767 -30268
rect 15703 -30412 15767 -30348
rect 15703 -30492 15767 -30428
rect 15703 -30572 15767 -30508
rect 15703 -30652 15767 -30588
rect 15703 -30732 15767 -30668
rect 15703 -30812 15767 -30748
rect 15703 -30892 15767 -30828
rect 15703 -30972 15767 -30908
rect 15703 -31052 15767 -30988
rect 15703 -31132 15767 -31068
rect 15703 -31212 15767 -31148
rect 15703 -31292 15767 -31228
rect 15703 -31372 15767 -31308
rect 15703 -31452 15767 -31388
rect 15703 -31532 15767 -31468
rect 15703 -31612 15767 -31548
rect 15703 -31692 15767 -31628
rect 15703 -31772 15767 -31708
rect 15703 -31852 15767 -31788
rect 15703 -31932 15767 -31868
rect 15703 -32012 15767 -31948
rect 15703 -32092 15767 -32028
rect 15703 -32172 15767 -32108
rect 15703 -32252 15767 -32188
rect 15703 -32332 15767 -32268
rect 15703 -32412 15767 -32348
rect 15703 -32492 15767 -32428
rect 15703 -32572 15767 -32508
rect 15703 -32652 15767 -32588
rect 15703 -32732 15767 -32668
rect 15703 -32812 15767 -32748
rect 15703 -32892 15767 -32828
rect 15703 -32972 15767 -32908
rect 15703 -33052 15767 -32988
rect 15703 -33132 15767 -33068
rect 15703 -33212 15767 -33148
rect 15703 -33292 15767 -33228
rect 15703 -33372 15767 -33308
rect 15703 -33452 15767 -33388
rect 15703 -33532 15767 -33468
rect 15703 -33612 15767 -33548
rect 15703 -33692 15767 -33628
rect 15703 -33772 15767 -33708
rect 15703 -33852 15767 -33788
rect 15703 -33932 15767 -33868
rect 15703 -34012 15767 -33948
rect 15703 -34092 15767 -34028
rect 15703 -34172 15767 -34108
rect 15703 -34252 15767 -34188
rect 15703 -34332 15767 -34268
rect 15703 -34412 15767 -34348
rect 15703 -34492 15767 -34428
rect 15703 -34572 15767 -34508
rect 22022 -28492 22086 -28428
rect 22022 -28572 22086 -28508
rect 22022 -28652 22086 -28588
rect 22022 -28732 22086 -28668
rect 22022 -28812 22086 -28748
rect 22022 -28892 22086 -28828
rect 22022 -28972 22086 -28908
rect 22022 -29052 22086 -28988
rect 22022 -29132 22086 -29068
rect 22022 -29212 22086 -29148
rect 22022 -29292 22086 -29228
rect 22022 -29372 22086 -29308
rect 22022 -29452 22086 -29388
rect 22022 -29532 22086 -29468
rect 22022 -29612 22086 -29548
rect 22022 -29692 22086 -29628
rect 22022 -29772 22086 -29708
rect 22022 -29852 22086 -29788
rect 22022 -29932 22086 -29868
rect 22022 -30012 22086 -29948
rect 22022 -30092 22086 -30028
rect 22022 -30172 22086 -30108
rect 22022 -30252 22086 -30188
rect 22022 -30332 22086 -30268
rect 22022 -30412 22086 -30348
rect 22022 -30492 22086 -30428
rect 22022 -30572 22086 -30508
rect 22022 -30652 22086 -30588
rect 22022 -30732 22086 -30668
rect 22022 -30812 22086 -30748
rect 22022 -30892 22086 -30828
rect 22022 -30972 22086 -30908
rect 22022 -31052 22086 -30988
rect 22022 -31132 22086 -31068
rect 22022 -31212 22086 -31148
rect 22022 -31292 22086 -31228
rect 22022 -31372 22086 -31308
rect 22022 -31452 22086 -31388
rect 22022 -31532 22086 -31468
rect 22022 -31612 22086 -31548
rect 22022 -31692 22086 -31628
rect 22022 -31772 22086 -31708
rect 22022 -31852 22086 -31788
rect 22022 -31932 22086 -31868
rect 22022 -32012 22086 -31948
rect 22022 -32092 22086 -32028
rect 22022 -32172 22086 -32108
rect 22022 -32252 22086 -32188
rect 22022 -32332 22086 -32268
rect 22022 -32412 22086 -32348
rect 22022 -32492 22086 -32428
rect 22022 -32572 22086 -32508
rect 22022 -32652 22086 -32588
rect 22022 -32732 22086 -32668
rect 22022 -32812 22086 -32748
rect 22022 -32892 22086 -32828
rect 22022 -32972 22086 -32908
rect 22022 -33052 22086 -32988
rect 22022 -33132 22086 -33068
rect 22022 -33212 22086 -33148
rect 22022 -33292 22086 -33228
rect 22022 -33372 22086 -33308
rect 22022 -33452 22086 -33388
rect 22022 -33532 22086 -33468
rect 22022 -33612 22086 -33548
rect 22022 -33692 22086 -33628
rect 22022 -33772 22086 -33708
rect 22022 -33852 22086 -33788
rect 22022 -33932 22086 -33868
rect 22022 -34012 22086 -33948
rect 22022 -34092 22086 -34028
rect 22022 -34172 22086 -34108
rect 22022 -34252 22086 -34188
rect 22022 -34332 22086 -34268
rect 22022 -34412 22086 -34348
rect 22022 -34492 22086 -34428
rect 22022 -34572 22086 -34508
rect 28341 -28492 28405 -28428
rect 28341 -28572 28405 -28508
rect 28341 -28652 28405 -28588
rect 28341 -28732 28405 -28668
rect 28341 -28812 28405 -28748
rect 28341 -28892 28405 -28828
rect 28341 -28972 28405 -28908
rect 28341 -29052 28405 -28988
rect 28341 -29132 28405 -29068
rect 28341 -29212 28405 -29148
rect 28341 -29292 28405 -29228
rect 28341 -29372 28405 -29308
rect 28341 -29452 28405 -29388
rect 28341 -29532 28405 -29468
rect 28341 -29612 28405 -29548
rect 28341 -29692 28405 -29628
rect 28341 -29772 28405 -29708
rect 28341 -29852 28405 -29788
rect 28341 -29932 28405 -29868
rect 28341 -30012 28405 -29948
rect 28341 -30092 28405 -30028
rect 28341 -30172 28405 -30108
rect 28341 -30252 28405 -30188
rect 28341 -30332 28405 -30268
rect 28341 -30412 28405 -30348
rect 28341 -30492 28405 -30428
rect 28341 -30572 28405 -30508
rect 28341 -30652 28405 -30588
rect 28341 -30732 28405 -30668
rect 28341 -30812 28405 -30748
rect 28341 -30892 28405 -30828
rect 28341 -30972 28405 -30908
rect 28341 -31052 28405 -30988
rect 28341 -31132 28405 -31068
rect 28341 -31212 28405 -31148
rect 28341 -31292 28405 -31228
rect 28341 -31372 28405 -31308
rect 28341 -31452 28405 -31388
rect 28341 -31532 28405 -31468
rect 28341 -31612 28405 -31548
rect 28341 -31692 28405 -31628
rect 28341 -31772 28405 -31708
rect 28341 -31852 28405 -31788
rect 28341 -31932 28405 -31868
rect 28341 -32012 28405 -31948
rect 28341 -32092 28405 -32028
rect 28341 -32172 28405 -32108
rect 28341 -32252 28405 -32188
rect 28341 -32332 28405 -32268
rect 28341 -32412 28405 -32348
rect 28341 -32492 28405 -32428
rect 28341 -32572 28405 -32508
rect 28341 -32652 28405 -32588
rect 28341 -32732 28405 -32668
rect 28341 -32812 28405 -32748
rect 28341 -32892 28405 -32828
rect 28341 -32972 28405 -32908
rect 28341 -33052 28405 -32988
rect 28341 -33132 28405 -33068
rect 28341 -33212 28405 -33148
rect 28341 -33292 28405 -33228
rect 28341 -33372 28405 -33308
rect 28341 -33452 28405 -33388
rect 28341 -33532 28405 -33468
rect 28341 -33612 28405 -33548
rect 28341 -33692 28405 -33628
rect 28341 -33772 28405 -33708
rect 28341 -33852 28405 -33788
rect 28341 -33932 28405 -33868
rect 28341 -34012 28405 -33948
rect 28341 -34092 28405 -34028
rect 28341 -34172 28405 -34108
rect 28341 -34252 28405 -34188
rect 28341 -34332 28405 -34268
rect 28341 -34412 28405 -34348
rect 28341 -34492 28405 -34428
rect 28341 -34572 28405 -34508
rect 34660 -28492 34724 -28428
rect 34660 -28572 34724 -28508
rect 34660 -28652 34724 -28588
rect 34660 -28732 34724 -28668
rect 34660 -28812 34724 -28748
rect 34660 -28892 34724 -28828
rect 34660 -28972 34724 -28908
rect 34660 -29052 34724 -28988
rect 34660 -29132 34724 -29068
rect 34660 -29212 34724 -29148
rect 34660 -29292 34724 -29228
rect 34660 -29372 34724 -29308
rect 34660 -29452 34724 -29388
rect 34660 -29532 34724 -29468
rect 34660 -29612 34724 -29548
rect 34660 -29692 34724 -29628
rect 34660 -29772 34724 -29708
rect 34660 -29852 34724 -29788
rect 34660 -29932 34724 -29868
rect 34660 -30012 34724 -29948
rect 34660 -30092 34724 -30028
rect 34660 -30172 34724 -30108
rect 34660 -30252 34724 -30188
rect 34660 -30332 34724 -30268
rect 34660 -30412 34724 -30348
rect 34660 -30492 34724 -30428
rect 34660 -30572 34724 -30508
rect 34660 -30652 34724 -30588
rect 34660 -30732 34724 -30668
rect 34660 -30812 34724 -30748
rect 34660 -30892 34724 -30828
rect 34660 -30972 34724 -30908
rect 34660 -31052 34724 -30988
rect 34660 -31132 34724 -31068
rect 34660 -31212 34724 -31148
rect 34660 -31292 34724 -31228
rect 34660 -31372 34724 -31308
rect 34660 -31452 34724 -31388
rect 34660 -31532 34724 -31468
rect 34660 -31612 34724 -31548
rect 34660 -31692 34724 -31628
rect 34660 -31772 34724 -31708
rect 34660 -31852 34724 -31788
rect 34660 -31932 34724 -31868
rect 34660 -32012 34724 -31948
rect 34660 -32092 34724 -32028
rect 34660 -32172 34724 -32108
rect 34660 -32252 34724 -32188
rect 34660 -32332 34724 -32268
rect 34660 -32412 34724 -32348
rect 34660 -32492 34724 -32428
rect 34660 -32572 34724 -32508
rect 34660 -32652 34724 -32588
rect 34660 -32732 34724 -32668
rect 34660 -32812 34724 -32748
rect 34660 -32892 34724 -32828
rect 34660 -32972 34724 -32908
rect 34660 -33052 34724 -32988
rect 34660 -33132 34724 -33068
rect 34660 -33212 34724 -33148
rect 34660 -33292 34724 -33228
rect 34660 -33372 34724 -33308
rect 34660 -33452 34724 -33388
rect 34660 -33532 34724 -33468
rect 34660 -33612 34724 -33548
rect 34660 -33692 34724 -33628
rect 34660 -33772 34724 -33708
rect 34660 -33852 34724 -33788
rect 34660 -33932 34724 -33868
rect 34660 -34012 34724 -33948
rect 34660 -34092 34724 -34028
rect 34660 -34172 34724 -34108
rect 34660 -34252 34724 -34188
rect 34660 -34332 34724 -34268
rect 34660 -34412 34724 -34348
rect 34660 -34492 34724 -34428
rect 34660 -34572 34724 -34508
rect 40979 -28492 41043 -28428
rect 40979 -28572 41043 -28508
rect 40979 -28652 41043 -28588
rect 40979 -28732 41043 -28668
rect 40979 -28812 41043 -28748
rect 40979 -28892 41043 -28828
rect 40979 -28972 41043 -28908
rect 40979 -29052 41043 -28988
rect 40979 -29132 41043 -29068
rect 40979 -29212 41043 -29148
rect 40979 -29292 41043 -29228
rect 40979 -29372 41043 -29308
rect 40979 -29452 41043 -29388
rect 40979 -29532 41043 -29468
rect 40979 -29612 41043 -29548
rect 40979 -29692 41043 -29628
rect 40979 -29772 41043 -29708
rect 40979 -29852 41043 -29788
rect 40979 -29932 41043 -29868
rect 40979 -30012 41043 -29948
rect 40979 -30092 41043 -30028
rect 40979 -30172 41043 -30108
rect 40979 -30252 41043 -30188
rect 40979 -30332 41043 -30268
rect 40979 -30412 41043 -30348
rect 40979 -30492 41043 -30428
rect 40979 -30572 41043 -30508
rect 40979 -30652 41043 -30588
rect 40979 -30732 41043 -30668
rect 40979 -30812 41043 -30748
rect 40979 -30892 41043 -30828
rect 40979 -30972 41043 -30908
rect 40979 -31052 41043 -30988
rect 40979 -31132 41043 -31068
rect 40979 -31212 41043 -31148
rect 40979 -31292 41043 -31228
rect 40979 -31372 41043 -31308
rect 40979 -31452 41043 -31388
rect 40979 -31532 41043 -31468
rect 40979 -31612 41043 -31548
rect 40979 -31692 41043 -31628
rect 40979 -31772 41043 -31708
rect 40979 -31852 41043 -31788
rect 40979 -31932 41043 -31868
rect 40979 -32012 41043 -31948
rect 40979 -32092 41043 -32028
rect 40979 -32172 41043 -32108
rect 40979 -32252 41043 -32188
rect 40979 -32332 41043 -32268
rect 40979 -32412 41043 -32348
rect 40979 -32492 41043 -32428
rect 40979 -32572 41043 -32508
rect 40979 -32652 41043 -32588
rect 40979 -32732 41043 -32668
rect 40979 -32812 41043 -32748
rect 40979 -32892 41043 -32828
rect 40979 -32972 41043 -32908
rect 40979 -33052 41043 -32988
rect 40979 -33132 41043 -33068
rect 40979 -33212 41043 -33148
rect 40979 -33292 41043 -33228
rect 40979 -33372 41043 -33308
rect 40979 -33452 41043 -33388
rect 40979 -33532 41043 -33468
rect 40979 -33612 41043 -33548
rect 40979 -33692 41043 -33628
rect 40979 -33772 41043 -33708
rect 40979 -33852 41043 -33788
rect 40979 -33932 41043 -33868
rect 40979 -34012 41043 -33948
rect 40979 -34092 41043 -34028
rect 40979 -34172 41043 -34108
rect 40979 -34252 41043 -34188
rect 40979 -34332 41043 -34268
rect 40979 -34412 41043 -34348
rect 40979 -34492 41043 -34428
rect 40979 -34572 41043 -34508
rect 47298 -28492 47362 -28428
rect 47298 -28572 47362 -28508
rect 47298 -28652 47362 -28588
rect 47298 -28732 47362 -28668
rect 47298 -28812 47362 -28748
rect 47298 -28892 47362 -28828
rect 47298 -28972 47362 -28908
rect 47298 -29052 47362 -28988
rect 47298 -29132 47362 -29068
rect 47298 -29212 47362 -29148
rect 47298 -29292 47362 -29228
rect 47298 -29372 47362 -29308
rect 47298 -29452 47362 -29388
rect 47298 -29532 47362 -29468
rect 47298 -29612 47362 -29548
rect 47298 -29692 47362 -29628
rect 47298 -29772 47362 -29708
rect 47298 -29852 47362 -29788
rect 47298 -29932 47362 -29868
rect 47298 -30012 47362 -29948
rect 47298 -30092 47362 -30028
rect 47298 -30172 47362 -30108
rect 47298 -30252 47362 -30188
rect 47298 -30332 47362 -30268
rect 47298 -30412 47362 -30348
rect 47298 -30492 47362 -30428
rect 47298 -30572 47362 -30508
rect 47298 -30652 47362 -30588
rect 47298 -30732 47362 -30668
rect 47298 -30812 47362 -30748
rect 47298 -30892 47362 -30828
rect 47298 -30972 47362 -30908
rect 47298 -31052 47362 -30988
rect 47298 -31132 47362 -31068
rect 47298 -31212 47362 -31148
rect 47298 -31292 47362 -31228
rect 47298 -31372 47362 -31308
rect 47298 -31452 47362 -31388
rect 47298 -31532 47362 -31468
rect 47298 -31612 47362 -31548
rect 47298 -31692 47362 -31628
rect 47298 -31772 47362 -31708
rect 47298 -31852 47362 -31788
rect 47298 -31932 47362 -31868
rect 47298 -32012 47362 -31948
rect 47298 -32092 47362 -32028
rect 47298 -32172 47362 -32108
rect 47298 -32252 47362 -32188
rect 47298 -32332 47362 -32268
rect 47298 -32412 47362 -32348
rect 47298 -32492 47362 -32428
rect 47298 -32572 47362 -32508
rect 47298 -32652 47362 -32588
rect 47298 -32732 47362 -32668
rect 47298 -32812 47362 -32748
rect 47298 -32892 47362 -32828
rect 47298 -32972 47362 -32908
rect 47298 -33052 47362 -32988
rect 47298 -33132 47362 -33068
rect 47298 -33212 47362 -33148
rect 47298 -33292 47362 -33228
rect 47298 -33372 47362 -33308
rect 47298 -33452 47362 -33388
rect 47298 -33532 47362 -33468
rect 47298 -33612 47362 -33548
rect 47298 -33692 47362 -33628
rect 47298 -33772 47362 -33708
rect 47298 -33852 47362 -33788
rect 47298 -33932 47362 -33868
rect 47298 -34012 47362 -33948
rect 47298 -34092 47362 -34028
rect 47298 -34172 47362 -34108
rect 47298 -34252 47362 -34188
rect 47298 -34332 47362 -34268
rect 47298 -34412 47362 -34348
rect 47298 -34492 47362 -34428
rect 47298 -34572 47362 -34508
rect -41168 -34792 -41104 -34728
rect -41168 -34872 -41104 -34808
rect -41168 -34952 -41104 -34888
rect -41168 -35032 -41104 -34968
rect -41168 -35112 -41104 -35048
rect -41168 -35192 -41104 -35128
rect -41168 -35272 -41104 -35208
rect -41168 -35352 -41104 -35288
rect -41168 -35432 -41104 -35368
rect -41168 -35512 -41104 -35448
rect -41168 -35592 -41104 -35528
rect -41168 -35672 -41104 -35608
rect -41168 -35752 -41104 -35688
rect -41168 -35832 -41104 -35768
rect -41168 -35912 -41104 -35848
rect -41168 -35992 -41104 -35928
rect -41168 -36072 -41104 -36008
rect -41168 -36152 -41104 -36088
rect -41168 -36232 -41104 -36168
rect -41168 -36312 -41104 -36248
rect -41168 -36392 -41104 -36328
rect -41168 -36472 -41104 -36408
rect -41168 -36552 -41104 -36488
rect -41168 -36632 -41104 -36568
rect -41168 -36712 -41104 -36648
rect -41168 -36792 -41104 -36728
rect -41168 -36872 -41104 -36808
rect -41168 -36952 -41104 -36888
rect -41168 -37032 -41104 -36968
rect -41168 -37112 -41104 -37048
rect -41168 -37192 -41104 -37128
rect -41168 -37272 -41104 -37208
rect -41168 -37352 -41104 -37288
rect -41168 -37432 -41104 -37368
rect -41168 -37512 -41104 -37448
rect -41168 -37592 -41104 -37528
rect -41168 -37672 -41104 -37608
rect -41168 -37752 -41104 -37688
rect -41168 -37832 -41104 -37768
rect -41168 -37912 -41104 -37848
rect -41168 -37992 -41104 -37928
rect -41168 -38072 -41104 -38008
rect -41168 -38152 -41104 -38088
rect -41168 -38232 -41104 -38168
rect -41168 -38312 -41104 -38248
rect -41168 -38392 -41104 -38328
rect -41168 -38472 -41104 -38408
rect -41168 -38552 -41104 -38488
rect -41168 -38632 -41104 -38568
rect -41168 -38712 -41104 -38648
rect -41168 -38792 -41104 -38728
rect -41168 -38872 -41104 -38808
rect -41168 -38952 -41104 -38888
rect -41168 -39032 -41104 -38968
rect -41168 -39112 -41104 -39048
rect -41168 -39192 -41104 -39128
rect -41168 -39272 -41104 -39208
rect -41168 -39352 -41104 -39288
rect -41168 -39432 -41104 -39368
rect -41168 -39512 -41104 -39448
rect -41168 -39592 -41104 -39528
rect -41168 -39672 -41104 -39608
rect -41168 -39752 -41104 -39688
rect -41168 -39832 -41104 -39768
rect -41168 -39912 -41104 -39848
rect -41168 -39992 -41104 -39928
rect -41168 -40072 -41104 -40008
rect -41168 -40152 -41104 -40088
rect -41168 -40232 -41104 -40168
rect -41168 -40312 -41104 -40248
rect -41168 -40392 -41104 -40328
rect -41168 -40472 -41104 -40408
rect -41168 -40552 -41104 -40488
rect -41168 -40632 -41104 -40568
rect -41168 -40712 -41104 -40648
rect -41168 -40792 -41104 -40728
rect -41168 -40872 -41104 -40808
rect -34849 -34792 -34785 -34728
rect -34849 -34872 -34785 -34808
rect -34849 -34952 -34785 -34888
rect -34849 -35032 -34785 -34968
rect -34849 -35112 -34785 -35048
rect -34849 -35192 -34785 -35128
rect -34849 -35272 -34785 -35208
rect -34849 -35352 -34785 -35288
rect -34849 -35432 -34785 -35368
rect -34849 -35512 -34785 -35448
rect -34849 -35592 -34785 -35528
rect -34849 -35672 -34785 -35608
rect -34849 -35752 -34785 -35688
rect -34849 -35832 -34785 -35768
rect -34849 -35912 -34785 -35848
rect -34849 -35992 -34785 -35928
rect -34849 -36072 -34785 -36008
rect -34849 -36152 -34785 -36088
rect -34849 -36232 -34785 -36168
rect -34849 -36312 -34785 -36248
rect -34849 -36392 -34785 -36328
rect -34849 -36472 -34785 -36408
rect -34849 -36552 -34785 -36488
rect -34849 -36632 -34785 -36568
rect -34849 -36712 -34785 -36648
rect -34849 -36792 -34785 -36728
rect -34849 -36872 -34785 -36808
rect -34849 -36952 -34785 -36888
rect -34849 -37032 -34785 -36968
rect -34849 -37112 -34785 -37048
rect -34849 -37192 -34785 -37128
rect -34849 -37272 -34785 -37208
rect -34849 -37352 -34785 -37288
rect -34849 -37432 -34785 -37368
rect -34849 -37512 -34785 -37448
rect -34849 -37592 -34785 -37528
rect -34849 -37672 -34785 -37608
rect -34849 -37752 -34785 -37688
rect -34849 -37832 -34785 -37768
rect -34849 -37912 -34785 -37848
rect -34849 -37992 -34785 -37928
rect -34849 -38072 -34785 -38008
rect -34849 -38152 -34785 -38088
rect -34849 -38232 -34785 -38168
rect -34849 -38312 -34785 -38248
rect -34849 -38392 -34785 -38328
rect -34849 -38472 -34785 -38408
rect -34849 -38552 -34785 -38488
rect -34849 -38632 -34785 -38568
rect -34849 -38712 -34785 -38648
rect -34849 -38792 -34785 -38728
rect -34849 -38872 -34785 -38808
rect -34849 -38952 -34785 -38888
rect -34849 -39032 -34785 -38968
rect -34849 -39112 -34785 -39048
rect -34849 -39192 -34785 -39128
rect -34849 -39272 -34785 -39208
rect -34849 -39352 -34785 -39288
rect -34849 -39432 -34785 -39368
rect -34849 -39512 -34785 -39448
rect -34849 -39592 -34785 -39528
rect -34849 -39672 -34785 -39608
rect -34849 -39752 -34785 -39688
rect -34849 -39832 -34785 -39768
rect -34849 -39912 -34785 -39848
rect -34849 -39992 -34785 -39928
rect -34849 -40072 -34785 -40008
rect -34849 -40152 -34785 -40088
rect -34849 -40232 -34785 -40168
rect -34849 -40312 -34785 -40248
rect -34849 -40392 -34785 -40328
rect -34849 -40472 -34785 -40408
rect -34849 -40552 -34785 -40488
rect -34849 -40632 -34785 -40568
rect -34849 -40712 -34785 -40648
rect -34849 -40792 -34785 -40728
rect -34849 -40872 -34785 -40808
rect -28530 -34792 -28466 -34728
rect -28530 -34872 -28466 -34808
rect -28530 -34952 -28466 -34888
rect -28530 -35032 -28466 -34968
rect -28530 -35112 -28466 -35048
rect -28530 -35192 -28466 -35128
rect -28530 -35272 -28466 -35208
rect -28530 -35352 -28466 -35288
rect -28530 -35432 -28466 -35368
rect -28530 -35512 -28466 -35448
rect -28530 -35592 -28466 -35528
rect -28530 -35672 -28466 -35608
rect -28530 -35752 -28466 -35688
rect -28530 -35832 -28466 -35768
rect -28530 -35912 -28466 -35848
rect -28530 -35992 -28466 -35928
rect -28530 -36072 -28466 -36008
rect -28530 -36152 -28466 -36088
rect -28530 -36232 -28466 -36168
rect -28530 -36312 -28466 -36248
rect -28530 -36392 -28466 -36328
rect -28530 -36472 -28466 -36408
rect -28530 -36552 -28466 -36488
rect -28530 -36632 -28466 -36568
rect -28530 -36712 -28466 -36648
rect -28530 -36792 -28466 -36728
rect -28530 -36872 -28466 -36808
rect -28530 -36952 -28466 -36888
rect -28530 -37032 -28466 -36968
rect -28530 -37112 -28466 -37048
rect -28530 -37192 -28466 -37128
rect -28530 -37272 -28466 -37208
rect -28530 -37352 -28466 -37288
rect -28530 -37432 -28466 -37368
rect -28530 -37512 -28466 -37448
rect -28530 -37592 -28466 -37528
rect -28530 -37672 -28466 -37608
rect -28530 -37752 -28466 -37688
rect -28530 -37832 -28466 -37768
rect -28530 -37912 -28466 -37848
rect -28530 -37992 -28466 -37928
rect -28530 -38072 -28466 -38008
rect -28530 -38152 -28466 -38088
rect -28530 -38232 -28466 -38168
rect -28530 -38312 -28466 -38248
rect -28530 -38392 -28466 -38328
rect -28530 -38472 -28466 -38408
rect -28530 -38552 -28466 -38488
rect -28530 -38632 -28466 -38568
rect -28530 -38712 -28466 -38648
rect -28530 -38792 -28466 -38728
rect -28530 -38872 -28466 -38808
rect -28530 -38952 -28466 -38888
rect -28530 -39032 -28466 -38968
rect -28530 -39112 -28466 -39048
rect -28530 -39192 -28466 -39128
rect -28530 -39272 -28466 -39208
rect -28530 -39352 -28466 -39288
rect -28530 -39432 -28466 -39368
rect -28530 -39512 -28466 -39448
rect -28530 -39592 -28466 -39528
rect -28530 -39672 -28466 -39608
rect -28530 -39752 -28466 -39688
rect -28530 -39832 -28466 -39768
rect -28530 -39912 -28466 -39848
rect -28530 -39992 -28466 -39928
rect -28530 -40072 -28466 -40008
rect -28530 -40152 -28466 -40088
rect -28530 -40232 -28466 -40168
rect -28530 -40312 -28466 -40248
rect -28530 -40392 -28466 -40328
rect -28530 -40472 -28466 -40408
rect -28530 -40552 -28466 -40488
rect -28530 -40632 -28466 -40568
rect -28530 -40712 -28466 -40648
rect -28530 -40792 -28466 -40728
rect -28530 -40872 -28466 -40808
rect -22211 -34792 -22147 -34728
rect -22211 -34872 -22147 -34808
rect -22211 -34952 -22147 -34888
rect -22211 -35032 -22147 -34968
rect -22211 -35112 -22147 -35048
rect -22211 -35192 -22147 -35128
rect -22211 -35272 -22147 -35208
rect -22211 -35352 -22147 -35288
rect -22211 -35432 -22147 -35368
rect -22211 -35512 -22147 -35448
rect -22211 -35592 -22147 -35528
rect -22211 -35672 -22147 -35608
rect -22211 -35752 -22147 -35688
rect -22211 -35832 -22147 -35768
rect -22211 -35912 -22147 -35848
rect -22211 -35992 -22147 -35928
rect -22211 -36072 -22147 -36008
rect -22211 -36152 -22147 -36088
rect -22211 -36232 -22147 -36168
rect -22211 -36312 -22147 -36248
rect -22211 -36392 -22147 -36328
rect -22211 -36472 -22147 -36408
rect -22211 -36552 -22147 -36488
rect -22211 -36632 -22147 -36568
rect -22211 -36712 -22147 -36648
rect -22211 -36792 -22147 -36728
rect -22211 -36872 -22147 -36808
rect -22211 -36952 -22147 -36888
rect -22211 -37032 -22147 -36968
rect -22211 -37112 -22147 -37048
rect -22211 -37192 -22147 -37128
rect -22211 -37272 -22147 -37208
rect -22211 -37352 -22147 -37288
rect -22211 -37432 -22147 -37368
rect -22211 -37512 -22147 -37448
rect -22211 -37592 -22147 -37528
rect -22211 -37672 -22147 -37608
rect -22211 -37752 -22147 -37688
rect -22211 -37832 -22147 -37768
rect -22211 -37912 -22147 -37848
rect -22211 -37992 -22147 -37928
rect -22211 -38072 -22147 -38008
rect -22211 -38152 -22147 -38088
rect -22211 -38232 -22147 -38168
rect -22211 -38312 -22147 -38248
rect -22211 -38392 -22147 -38328
rect -22211 -38472 -22147 -38408
rect -22211 -38552 -22147 -38488
rect -22211 -38632 -22147 -38568
rect -22211 -38712 -22147 -38648
rect -22211 -38792 -22147 -38728
rect -22211 -38872 -22147 -38808
rect -22211 -38952 -22147 -38888
rect -22211 -39032 -22147 -38968
rect -22211 -39112 -22147 -39048
rect -22211 -39192 -22147 -39128
rect -22211 -39272 -22147 -39208
rect -22211 -39352 -22147 -39288
rect -22211 -39432 -22147 -39368
rect -22211 -39512 -22147 -39448
rect -22211 -39592 -22147 -39528
rect -22211 -39672 -22147 -39608
rect -22211 -39752 -22147 -39688
rect -22211 -39832 -22147 -39768
rect -22211 -39912 -22147 -39848
rect -22211 -39992 -22147 -39928
rect -22211 -40072 -22147 -40008
rect -22211 -40152 -22147 -40088
rect -22211 -40232 -22147 -40168
rect -22211 -40312 -22147 -40248
rect -22211 -40392 -22147 -40328
rect -22211 -40472 -22147 -40408
rect -22211 -40552 -22147 -40488
rect -22211 -40632 -22147 -40568
rect -22211 -40712 -22147 -40648
rect -22211 -40792 -22147 -40728
rect -22211 -40872 -22147 -40808
rect -15892 -34792 -15828 -34728
rect -15892 -34872 -15828 -34808
rect -15892 -34952 -15828 -34888
rect -15892 -35032 -15828 -34968
rect -15892 -35112 -15828 -35048
rect -15892 -35192 -15828 -35128
rect -15892 -35272 -15828 -35208
rect -15892 -35352 -15828 -35288
rect -15892 -35432 -15828 -35368
rect -15892 -35512 -15828 -35448
rect -15892 -35592 -15828 -35528
rect -15892 -35672 -15828 -35608
rect -15892 -35752 -15828 -35688
rect -15892 -35832 -15828 -35768
rect -15892 -35912 -15828 -35848
rect -15892 -35992 -15828 -35928
rect -15892 -36072 -15828 -36008
rect -15892 -36152 -15828 -36088
rect -15892 -36232 -15828 -36168
rect -15892 -36312 -15828 -36248
rect -15892 -36392 -15828 -36328
rect -15892 -36472 -15828 -36408
rect -15892 -36552 -15828 -36488
rect -15892 -36632 -15828 -36568
rect -15892 -36712 -15828 -36648
rect -15892 -36792 -15828 -36728
rect -15892 -36872 -15828 -36808
rect -15892 -36952 -15828 -36888
rect -15892 -37032 -15828 -36968
rect -15892 -37112 -15828 -37048
rect -15892 -37192 -15828 -37128
rect -15892 -37272 -15828 -37208
rect -15892 -37352 -15828 -37288
rect -15892 -37432 -15828 -37368
rect -15892 -37512 -15828 -37448
rect -15892 -37592 -15828 -37528
rect -15892 -37672 -15828 -37608
rect -15892 -37752 -15828 -37688
rect -15892 -37832 -15828 -37768
rect -15892 -37912 -15828 -37848
rect -15892 -37992 -15828 -37928
rect -15892 -38072 -15828 -38008
rect -15892 -38152 -15828 -38088
rect -15892 -38232 -15828 -38168
rect -15892 -38312 -15828 -38248
rect -15892 -38392 -15828 -38328
rect -15892 -38472 -15828 -38408
rect -15892 -38552 -15828 -38488
rect -15892 -38632 -15828 -38568
rect -15892 -38712 -15828 -38648
rect -15892 -38792 -15828 -38728
rect -15892 -38872 -15828 -38808
rect -15892 -38952 -15828 -38888
rect -15892 -39032 -15828 -38968
rect -15892 -39112 -15828 -39048
rect -15892 -39192 -15828 -39128
rect -15892 -39272 -15828 -39208
rect -15892 -39352 -15828 -39288
rect -15892 -39432 -15828 -39368
rect -15892 -39512 -15828 -39448
rect -15892 -39592 -15828 -39528
rect -15892 -39672 -15828 -39608
rect -15892 -39752 -15828 -39688
rect -15892 -39832 -15828 -39768
rect -15892 -39912 -15828 -39848
rect -15892 -39992 -15828 -39928
rect -15892 -40072 -15828 -40008
rect -15892 -40152 -15828 -40088
rect -15892 -40232 -15828 -40168
rect -15892 -40312 -15828 -40248
rect -15892 -40392 -15828 -40328
rect -15892 -40472 -15828 -40408
rect -15892 -40552 -15828 -40488
rect -15892 -40632 -15828 -40568
rect -15892 -40712 -15828 -40648
rect -15892 -40792 -15828 -40728
rect -15892 -40872 -15828 -40808
rect -9573 -34792 -9509 -34728
rect -9573 -34872 -9509 -34808
rect -9573 -34952 -9509 -34888
rect -9573 -35032 -9509 -34968
rect -9573 -35112 -9509 -35048
rect -9573 -35192 -9509 -35128
rect -9573 -35272 -9509 -35208
rect -9573 -35352 -9509 -35288
rect -9573 -35432 -9509 -35368
rect -9573 -35512 -9509 -35448
rect -9573 -35592 -9509 -35528
rect -9573 -35672 -9509 -35608
rect -9573 -35752 -9509 -35688
rect -9573 -35832 -9509 -35768
rect -9573 -35912 -9509 -35848
rect -9573 -35992 -9509 -35928
rect -9573 -36072 -9509 -36008
rect -9573 -36152 -9509 -36088
rect -9573 -36232 -9509 -36168
rect -9573 -36312 -9509 -36248
rect -9573 -36392 -9509 -36328
rect -9573 -36472 -9509 -36408
rect -9573 -36552 -9509 -36488
rect -9573 -36632 -9509 -36568
rect -9573 -36712 -9509 -36648
rect -9573 -36792 -9509 -36728
rect -9573 -36872 -9509 -36808
rect -9573 -36952 -9509 -36888
rect -9573 -37032 -9509 -36968
rect -9573 -37112 -9509 -37048
rect -9573 -37192 -9509 -37128
rect -9573 -37272 -9509 -37208
rect -9573 -37352 -9509 -37288
rect -9573 -37432 -9509 -37368
rect -9573 -37512 -9509 -37448
rect -9573 -37592 -9509 -37528
rect -9573 -37672 -9509 -37608
rect -9573 -37752 -9509 -37688
rect -9573 -37832 -9509 -37768
rect -9573 -37912 -9509 -37848
rect -9573 -37992 -9509 -37928
rect -9573 -38072 -9509 -38008
rect -9573 -38152 -9509 -38088
rect -9573 -38232 -9509 -38168
rect -9573 -38312 -9509 -38248
rect -9573 -38392 -9509 -38328
rect -9573 -38472 -9509 -38408
rect -9573 -38552 -9509 -38488
rect -9573 -38632 -9509 -38568
rect -9573 -38712 -9509 -38648
rect -9573 -38792 -9509 -38728
rect -9573 -38872 -9509 -38808
rect -9573 -38952 -9509 -38888
rect -9573 -39032 -9509 -38968
rect -9573 -39112 -9509 -39048
rect -9573 -39192 -9509 -39128
rect -9573 -39272 -9509 -39208
rect -9573 -39352 -9509 -39288
rect -9573 -39432 -9509 -39368
rect -9573 -39512 -9509 -39448
rect -9573 -39592 -9509 -39528
rect -9573 -39672 -9509 -39608
rect -9573 -39752 -9509 -39688
rect -9573 -39832 -9509 -39768
rect -9573 -39912 -9509 -39848
rect -9573 -39992 -9509 -39928
rect -9573 -40072 -9509 -40008
rect -9573 -40152 -9509 -40088
rect -9573 -40232 -9509 -40168
rect -9573 -40312 -9509 -40248
rect -9573 -40392 -9509 -40328
rect -9573 -40472 -9509 -40408
rect -9573 -40552 -9509 -40488
rect -9573 -40632 -9509 -40568
rect -9573 -40712 -9509 -40648
rect -9573 -40792 -9509 -40728
rect -9573 -40872 -9509 -40808
rect -3254 -34792 -3190 -34728
rect -3254 -34872 -3190 -34808
rect -3254 -34952 -3190 -34888
rect -3254 -35032 -3190 -34968
rect -3254 -35112 -3190 -35048
rect -3254 -35192 -3190 -35128
rect -3254 -35272 -3190 -35208
rect -3254 -35352 -3190 -35288
rect -3254 -35432 -3190 -35368
rect -3254 -35512 -3190 -35448
rect -3254 -35592 -3190 -35528
rect -3254 -35672 -3190 -35608
rect -3254 -35752 -3190 -35688
rect -3254 -35832 -3190 -35768
rect -3254 -35912 -3190 -35848
rect -3254 -35992 -3190 -35928
rect -3254 -36072 -3190 -36008
rect -3254 -36152 -3190 -36088
rect -3254 -36232 -3190 -36168
rect -3254 -36312 -3190 -36248
rect -3254 -36392 -3190 -36328
rect -3254 -36472 -3190 -36408
rect -3254 -36552 -3190 -36488
rect -3254 -36632 -3190 -36568
rect -3254 -36712 -3190 -36648
rect -3254 -36792 -3190 -36728
rect -3254 -36872 -3190 -36808
rect -3254 -36952 -3190 -36888
rect -3254 -37032 -3190 -36968
rect -3254 -37112 -3190 -37048
rect -3254 -37192 -3190 -37128
rect -3254 -37272 -3190 -37208
rect -3254 -37352 -3190 -37288
rect -3254 -37432 -3190 -37368
rect -3254 -37512 -3190 -37448
rect -3254 -37592 -3190 -37528
rect -3254 -37672 -3190 -37608
rect -3254 -37752 -3190 -37688
rect -3254 -37832 -3190 -37768
rect -3254 -37912 -3190 -37848
rect -3254 -37992 -3190 -37928
rect -3254 -38072 -3190 -38008
rect -3254 -38152 -3190 -38088
rect -3254 -38232 -3190 -38168
rect -3254 -38312 -3190 -38248
rect -3254 -38392 -3190 -38328
rect -3254 -38472 -3190 -38408
rect -3254 -38552 -3190 -38488
rect -3254 -38632 -3190 -38568
rect -3254 -38712 -3190 -38648
rect -3254 -38792 -3190 -38728
rect -3254 -38872 -3190 -38808
rect -3254 -38952 -3190 -38888
rect -3254 -39032 -3190 -38968
rect -3254 -39112 -3190 -39048
rect -3254 -39192 -3190 -39128
rect -3254 -39272 -3190 -39208
rect -3254 -39352 -3190 -39288
rect -3254 -39432 -3190 -39368
rect -3254 -39512 -3190 -39448
rect -3254 -39592 -3190 -39528
rect -3254 -39672 -3190 -39608
rect -3254 -39752 -3190 -39688
rect -3254 -39832 -3190 -39768
rect -3254 -39912 -3190 -39848
rect -3254 -39992 -3190 -39928
rect -3254 -40072 -3190 -40008
rect -3254 -40152 -3190 -40088
rect -3254 -40232 -3190 -40168
rect -3254 -40312 -3190 -40248
rect -3254 -40392 -3190 -40328
rect -3254 -40472 -3190 -40408
rect -3254 -40552 -3190 -40488
rect -3254 -40632 -3190 -40568
rect -3254 -40712 -3190 -40648
rect -3254 -40792 -3190 -40728
rect -3254 -40872 -3190 -40808
rect 3065 -34792 3129 -34728
rect 3065 -34872 3129 -34808
rect 3065 -34952 3129 -34888
rect 3065 -35032 3129 -34968
rect 3065 -35112 3129 -35048
rect 3065 -35192 3129 -35128
rect 3065 -35272 3129 -35208
rect 3065 -35352 3129 -35288
rect 3065 -35432 3129 -35368
rect 3065 -35512 3129 -35448
rect 3065 -35592 3129 -35528
rect 3065 -35672 3129 -35608
rect 3065 -35752 3129 -35688
rect 3065 -35832 3129 -35768
rect 3065 -35912 3129 -35848
rect 3065 -35992 3129 -35928
rect 3065 -36072 3129 -36008
rect 3065 -36152 3129 -36088
rect 3065 -36232 3129 -36168
rect 3065 -36312 3129 -36248
rect 3065 -36392 3129 -36328
rect 3065 -36472 3129 -36408
rect 3065 -36552 3129 -36488
rect 3065 -36632 3129 -36568
rect 3065 -36712 3129 -36648
rect 3065 -36792 3129 -36728
rect 3065 -36872 3129 -36808
rect 3065 -36952 3129 -36888
rect 3065 -37032 3129 -36968
rect 3065 -37112 3129 -37048
rect 3065 -37192 3129 -37128
rect 3065 -37272 3129 -37208
rect 3065 -37352 3129 -37288
rect 3065 -37432 3129 -37368
rect 3065 -37512 3129 -37448
rect 3065 -37592 3129 -37528
rect 3065 -37672 3129 -37608
rect 3065 -37752 3129 -37688
rect 3065 -37832 3129 -37768
rect 3065 -37912 3129 -37848
rect 3065 -37992 3129 -37928
rect 3065 -38072 3129 -38008
rect 3065 -38152 3129 -38088
rect 3065 -38232 3129 -38168
rect 3065 -38312 3129 -38248
rect 3065 -38392 3129 -38328
rect 3065 -38472 3129 -38408
rect 3065 -38552 3129 -38488
rect 3065 -38632 3129 -38568
rect 3065 -38712 3129 -38648
rect 3065 -38792 3129 -38728
rect 3065 -38872 3129 -38808
rect 3065 -38952 3129 -38888
rect 3065 -39032 3129 -38968
rect 3065 -39112 3129 -39048
rect 3065 -39192 3129 -39128
rect 3065 -39272 3129 -39208
rect 3065 -39352 3129 -39288
rect 3065 -39432 3129 -39368
rect 3065 -39512 3129 -39448
rect 3065 -39592 3129 -39528
rect 3065 -39672 3129 -39608
rect 3065 -39752 3129 -39688
rect 3065 -39832 3129 -39768
rect 3065 -39912 3129 -39848
rect 3065 -39992 3129 -39928
rect 3065 -40072 3129 -40008
rect 3065 -40152 3129 -40088
rect 3065 -40232 3129 -40168
rect 3065 -40312 3129 -40248
rect 3065 -40392 3129 -40328
rect 3065 -40472 3129 -40408
rect 3065 -40552 3129 -40488
rect 3065 -40632 3129 -40568
rect 3065 -40712 3129 -40648
rect 3065 -40792 3129 -40728
rect 3065 -40872 3129 -40808
rect 9384 -34792 9448 -34728
rect 9384 -34872 9448 -34808
rect 9384 -34952 9448 -34888
rect 9384 -35032 9448 -34968
rect 9384 -35112 9448 -35048
rect 9384 -35192 9448 -35128
rect 9384 -35272 9448 -35208
rect 9384 -35352 9448 -35288
rect 9384 -35432 9448 -35368
rect 9384 -35512 9448 -35448
rect 9384 -35592 9448 -35528
rect 9384 -35672 9448 -35608
rect 9384 -35752 9448 -35688
rect 9384 -35832 9448 -35768
rect 9384 -35912 9448 -35848
rect 9384 -35992 9448 -35928
rect 9384 -36072 9448 -36008
rect 9384 -36152 9448 -36088
rect 9384 -36232 9448 -36168
rect 9384 -36312 9448 -36248
rect 9384 -36392 9448 -36328
rect 9384 -36472 9448 -36408
rect 9384 -36552 9448 -36488
rect 9384 -36632 9448 -36568
rect 9384 -36712 9448 -36648
rect 9384 -36792 9448 -36728
rect 9384 -36872 9448 -36808
rect 9384 -36952 9448 -36888
rect 9384 -37032 9448 -36968
rect 9384 -37112 9448 -37048
rect 9384 -37192 9448 -37128
rect 9384 -37272 9448 -37208
rect 9384 -37352 9448 -37288
rect 9384 -37432 9448 -37368
rect 9384 -37512 9448 -37448
rect 9384 -37592 9448 -37528
rect 9384 -37672 9448 -37608
rect 9384 -37752 9448 -37688
rect 9384 -37832 9448 -37768
rect 9384 -37912 9448 -37848
rect 9384 -37992 9448 -37928
rect 9384 -38072 9448 -38008
rect 9384 -38152 9448 -38088
rect 9384 -38232 9448 -38168
rect 9384 -38312 9448 -38248
rect 9384 -38392 9448 -38328
rect 9384 -38472 9448 -38408
rect 9384 -38552 9448 -38488
rect 9384 -38632 9448 -38568
rect 9384 -38712 9448 -38648
rect 9384 -38792 9448 -38728
rect 9384 -38872 9448 -38808
rect 9384 -38952 9448 -38888
rect 9384 -39032 9448 -38968
rect 9384 -39112 9448 -39048
rect 9384 -39192 9448 -39128
rect 9384 -39272 9448 -39208
rect 9384 -39352 9448 -39288
rect 9384 -39432 9448 -39368
rect 9384 -39512 9448 -39448
rect 9384 -39592 9448 -39528
rect 9384 -39672 9448 -39608
rect 9384 -39752 9448 -39688
rect 9384 -39832 9448 -39768
rect 9384 -39912 9448 -39848
rect 9384 -39992 9448 -39928
rect 9384 -40072 9448 -40008
rect 9384 -40152 9448 -40088
rect 9384 -40232 9448 -40168
rect 9384 -40312 9448 -40248
rect 9384 -40392 9448 -40328
rect 9384 -40472 9448 -40408
rect 9384 -40552 9448 -40488
rect 9384 -40632 9448 -40568
rect 9384 -40712 9448 -40648
rect 9384 -40792 9448 -40728
rect 9384 -40872 9448 -40808
rect 15703 -34792 15767 -34728
rect 15703 -34872 15767 -34808
rect 15703 -34952 15767 -34888
rect 15703 -35032 15767 -34968
rect 15703 -35112 15767 -35048
rect 15703 -35192 15767 -35128
rect 15703 -35272 15767 -35208
rect 15703 -35352 15767 -35288
rect 15703 -35432 15767 -35368
rect 15703 -35512 15767 -35448
rect 15703 -35592 15767 -35528
rect 15703 -35672 15767 -35608
rect 15703 -35752 15767 -35688
rect 15703 -35832 15767 -35768
rect 15703 -35912 15767 -35848
rect 15703 -35992 15767 -35928
rect 15703 -36072 15767 -36008
rect 15703 -36152 15767 -36088
rect 15703 -36232 15767 -36168
rect 15703 -36312 15767 -36248
rect 15703 -36392 15767 -36328
rect 15703 -36472 15767 -36408
rect 15703 -36552 15767 -36488
rect 15703 -36632 15767 -36568
rect 15703 -36712 15767 -36648
rect 15703 -36792 15767 -36728
rect 15703 -36872 15767 -36808
rect 15703 -36952 15767 -36888
rect 15703 -37032 15767 -36968
rect 15703 -37112 15767 -37048
rect 15703 -37192 15767 -37128
rect 15703 -37272 15767 -37208
rect 15703 -37352 15767 -37288
rect 15703 -37432 15767 -37368
rect 15703 -37512 15767 -37448
rect 15703 -37592 15767 -37528
rect 15703 -37672 15767 -37608
rect 15703 -37752 15767 -37688
rect 15703 -37832 15767 -37768
rect 15703 -37912 15767 -37848
rect 15703 -37992 15767 -37928
rect 15703 -38072 15767 -38008
rect 15703 -38152 15767 -38088
rect 15703 -38232 15767 -38168
rect 15703 -38312 15767 -38248
rect 15703 -38392 15767 -38328
rect 15703 -38472 15767 -38408
rect 15703 -38552 15767 -38488
rect 15703 -38632 15767 -38568
rect 15703 -38712 15767 -38648
rect 15703 -38792 15767 -38728
rect 15703 -38872 15767 -38808
rect 15703 -38952 15767 -38888
rect 15703 -39032 15767 -38968
rect 15703 -39112 15767 -39048
rect 15703 -39192 15767 -39128
rect 15703 -39272 15767 -39208
rect 15703 -39352 15767 -39288
rect 15703 -39432 15767 -39368
rect 15703 -39512 15767 -39448
rect 15703 -39592 15767 -39528
rect 15703 -39672 15767 -39608
rect 15703 -39752 15767 -39688
rect 15703 -39832 15767 -39768
rect 15703 -39912 15767 -39848
rect 15703 -39992 15767 -39928
rect 15703 -40072 15767 -40008
rect 15703 -40152 15767 -40088
rect 15703 -40232 15767 -40168
rect 15703 -40312 15767 -40248
rect 15703 -40392 15767 -40328
rect 15703 -40472 15767 -40408
rect 15703 -40552 15767 -40488
rect 15703 -40632 15767 -40568
rect 15703 -40712 15767 -40648
rect 15703 -40792 15767 -40728
rect 15703 -40872 15767 -40808
rect 22022 -34792 22086 -34728
rect 22022 -34872 22086 -34808
rect 22022 -34952 22086 -34888
rect 22022 -35032 22086 -34968
rect 22022 -35112 22086 -35048
rect 22022 -35192 22086 -35128
rect 22022 -35272 22086 -35208
rect 22022 -35352 22086 -35288
rect 22022 -35432 22086 -35368
rect 22022 -35512 22086 -35448
rect 22022 -35592 22086 -35528
rect 22022 -35672 22086 -35608
rect 22022 -35752 22086 -35688
rect 22022 -35832 22086 -35768
rect 22022 -35912 22086 -35848
rect 22022 -35992 22086 -35928
rect 22022 -36072 22086 -36008
rect 22022 -36152 22086 -36088
rect 22022 -36232 22086 -36168
rect 22022 -36312 22086 -36248
rect 22022 -36392 22086 -36328
rect 22022 -36472 22086 -36408
rect 22022 -36552 22086 -36488
rect 22022 -36632 22086 -36568
rect 22022 -36712 22086 -36648
rect 22022 -36792 22086 -36728
rect 22022 -36872 22086 -36808
rect 22022 -36952 22086 -36888
rect 22022 -37032 22086 -36968
rect 22022 -37112 22086 -37048
rect 22022 -37192 22086 -37128
rect 22022 -37272 22086 -37208
rect 22022 -37352 22086 -37288
rect 22022 -37432 22086 -37368
rect 22022 -37512 22086 -37448
rect 22022 -37592 22086 -37528
rect 22022 -37672 22086 -37608
rect 22022 -37752 22086 -37688
rect 22022 -37832 22086 -37768
rect 22022 -37912 22086 -37848
rect 22022 -37992 22086 -37928
rect 22022 -38072 22086 -38008
rect 22022 -38152 22086 -38088
rect 22022 -38232 22086 -38168
rect 22022 -38312 22086 -38248
rect 22022 -38392 22086 -38328
rect 22022 -38472 22086 -38408
rect 22022 -38552 22086 -38488
rect 22022 -38632 22086 -38568
rect 22022 -38712 22086 -38648
rect 22022 -38792 22086 -38728
rect 22022 -38872 22086 -38808
rect 22022 -38952 22086 -38888
rect 22022 -39032 22086 -38968
rect 22022 -39112 22086 -39048
rect 22022 -39192 22086 -39128
rect 22022 -39272 22086 -39208
rect 22022 -39352 22086 -39288
rect 22022 -39432 22086 -39368
rect 22022 -39512 22086 -39448
rect 22022 -39592 22086 -39528
rect 22022 -39672 22086 -39608
rect 22022 -39752 22086 -39688
rect 22022 -39832 22086 -39768
rect 22022 -39912 22086 -39848
rect 22022 -39992 22086 -39928
rect 22022 -40072 22086 -40008
rect 22022 -40152 22086 -40088
rect 22022 -40232 22086 -40168
rect 22022 -40312 22086 -40248
rect 22022 -40392 22086 -40328
rect 22022 -40472 22086 -40408
rect 22022 -40552 22086 -40488
rect 22022 -40632 22086 -40568
rect 22022 -40712 22086 -40648
rect 22022 -40792 22086 -40728
rect 22022 -40872 22086 -40808
rect 28341 -34792 28405 -34728
rect 28341 -34872 28405 -34808
rect 28341 -34952 28405 -34888
rect 28341 -35032 28405 -34968
rect 28341 -35112 28405 -35048
rect 28341 -35192 28405 -35128
rect 28341 -35272 28405 -35208
rect 28341 -35352 28405 -35288
rect 28341 -35432 28405 -35368
rect 28341 -35512 28405 -35448
rect 28341 -35592 28405 -35528
rect 28341 -35672 28405 -35608
rect 28341 -35752 28405 -35688
rect 28341 -35832 28405 -35768
rect 28341 -35912 28405 -35848
rect 28341 -35992 28405 -35928
rect 28341 -36072 28405 -36008
rect 28341 -36152 28405 -36088
rect 28341 -36232 28405 -36168
rect 28341 -36312 28405 -36248
rect 28341 -36392 28405 -36328
rect 28341 -36472 28405 -36408
rect 28341 -36552 28405 -36488
rect 28341 -36632 28405 -36568
rect 28341 -36712 28405 -36648
rect 28341 -36792 28405 -36728
rect 28341 -36872 28405 -36808
rect 28341 -36952 28405 -36888
rect 28341 -37032 28405 -36968
rect 28341 -37112 28405 -37048
rect 28341 -37192 28405 -37128
rect 28341 -37272 28405 -37208
rect 28341 -37352 28405 -37288
rect 28341 -37432 28405 -37368
rect 28341 -37512 28405 -37448
rect 28341 -37592 28405 -37528
rect 28341 -37672 28405 -37608
rect 28341 -37752 28405 -37688
rect 28341 -37832 28405 -37768
rect 28341 -37912 28405 -37848
rect 28341 -37992 28405 -37928
rect 28341 -38072 28405 -38008
rect 28341 -38152 28405 -38088
rect 28341 -38232 28405 -38168
rect 28341 -38312 28405 -38248
rect 28341 -38392 28405 -38328
rect 28341 -38472 28405 -38408
rect 28341 -38552 28405 -38488
rect 28341 -38632 28405 -38568
rect 28341 -38712 28405 -38648
rect 28341 -38792 28405 -38728
rect 28341 -38872 28405 -38808
rect 28341 -38952 28405 -38888
rect 28341 -39032 28405 -38968
rect 28341 -39112 28405 -39048
rect 28341 -39192 28405 -39128
rect 28341 -39272 28405 -39208
rect 28341 -39352 28405 -39288
rect 28341 -39432 28405 -39368
rect 28341 -39512 28405 -39448
rect 28341 -39592 28405 -39528
rect 28341 -39672 28405 -39608
rect 28341 -39752 28405 -39688
rect 28341 -39832 28405 -39768
rect 28341 -39912 28405 -39848
rect 28341 -39992 28405 -39928
rect 28341 -40072 28405 -40008
rect 28341 -40152 28405 -40088
rect 28341 -40232 28405 -40168
rect 28341 -40312 28405 -40248
rect 28341 -40392 28405 -40328
rect 28341 -40472 28405 -40408
rect 28341 -40552 28405 -40488
rect 28341 -40632 28405 -40568
rect 28341 -40712 28405 -40648
rect 28341 -40792 28405 -40728
rect 28341 -40872 28405 -40808
rect 34660 -34792 34724 -34728
rect 34660 -34872 34724 -34808
rect 34660 -34952 34724 -34888
rect 34660 -35032 34724 -34968
rect 34660 -35112 34724 -35048
rect 34660 -35192 34724 -35128
rect 34660 -35272 34724 -35208
rect 34660 -35352 34724 -35288
rect 34660 -35432 34724 -35368
rect 34660 -35512 34724 -35448
rect 34660 -35592 34724 -35528
rect 34660 -35672 34724 -35608
rect 34660 -35752 34724 -35688
rect 34660 -35832 34724 -35768
rect 34660 -35912 34724 -35848
rect 34660 -35992 34724 -35928
rect 34660 -36072 34724 -36008
rect 34660 -36152 34724 -36088
rect 34660 -36232 34724 -36168
rect 34660 -36312 34724 -36248
rect 34660 -36392 34724 -36328
rect 34660 -36472 34724 -36408
rect 34660 -36552 34724 -36488
rect 34660 -36632 34724 -36568
rect 34660 -36712 34724 -36648
rect 34660 -36792 34724 -36728
rect 34660 -36872 34724 -36808
rect 34660 -36952 34724 -36888
rect 34660 -37032 34724 -36968
rect 34660 -37112 34724 -37048
rect 34660 -37192 34724 -37128
rect 34660 -37272 34724 -37208
rect 34660 -37352 34724 -37288
rect 34660 -37432 34724 -37368
rect 34660 -37512 34724 -37448
rect 34660 -37592 34724 -37528
rect 34660 -37672 34724 -37608
rect 34660 -37752 34724 -37688
rect 34660 -37832 34724 -37768
rect 34660 -37912 34724 -37848
rect 34660 -37992 34724 -37928
rect 34660 -38072 34724 -38008
rect 34660 -38152 34724 -38088
rect 34660 -38232 34724 -38168
rect 34660 -38312 34724 -38248
rect 34660 -38392 34724 -38328
rect 34660 -38472 34724 -38408
rect 34660 -38552 34724 -38488
rect 34660 -38632 34724 -38568
rect 34660 -38712 34724 -38648
rect 34660 -38792 34724 -38728
rect 34660 -38872 34724 -38808
rect 34660 -38952 34724 -38888
rect 34660 -39032 34724 -38968
rect 34660 -39112 34724 -39048
rect 34660 -39192 34724 -39128
rect 34660 -39272 34724 -39208
rect 34660 -39352 34724 -39288
rect 34660 -39432 34724 -39368
rect 34660 -39512 34724 -39448
rect 34660 -39592 34724 -39528
rect 34660 -39672 34724 -39608
rect 34660 -39752 34724 -39688
rect 34660 -39832 34724 -39768
rect 34660 -39912 34724 -39848
rect 34660 -39992 34724 -39928
rect 34660 -40072 34724 -40008
rect 34660 -40152 34724 -40088
rect 34660 -40232 34724 -40168
rect 34660 -40312 34724 -40248
rect 34660 -40392 34724 -40328
rect 34660 -40472 34724 -40408
rect 34660 -40552 34724 -40488
rect 34660 -40632 34724 -40568
rect 34660 -40712 34724 -40648
rect 34660 -40792 34724 -40728
rect 34660 -40872 34724 -40808
rect 40979 -34792 41043 -34728
rect 40979 -34872 41043 -34808
rect 40979 -34952 41043 -34888
rect 40979 -35032 41043 -34968
rect 40979 -35112 41043 -35048
rect 40979 -35192 41043 -35128
rect 40979 -35272 41043 -35208
rect 40979 -35352 41043 -35288
rect 40979 -35432 41043 -35368
rect 40979 -35512 41043 -35448
rect 40979 -35592 41043 -35528
rect 40979 -35672 41043 -35608
rect 40979 -35752 41043 -35688
rect 40979 -35832 41043 -35768
rect 40979 -35912 41043 -35848
rect 40979 -35992 41043 -35928
rect 40979 -36072 41043 -36008
rect 40979 -36152 41043 -36088
rect 40979 -36232 41043 -36168
rect 40979 -36312 41043 -36248
rect 40979 -36392 41043 -36328
rect 40979 -36472 41043 -36408
rect 40979 -36552 41043 -36488
rect 40979 -36632 41043 -36568
rect 40979 -36712 41043 -36648
rect 40979 -36792 41043 -36728
rect 40979 -36872 41043 -36808
rect 40979 -36952 41043 -36888
rect 40979 -37032 41043 -36968
rect 40979 -37112 41043 -37048
rect 40979 -37192 41043 -37128
rect 40979 -37272 41043 -37208
rect 40979 -37352 41043 -37288
rect 40979 -37432 41043 -37368
rect 40979 -37512 41043 -37448
rect 40979 -37592 41043 -37528
rect 40979 -37672 41043 -37608
rect 40979 -37752 41043 -37688
rect 40979 -37832 41043 -37768
rect 40979 -37912 41043 -37848
rect 40979 -37992 41043 -37928
rect 40979 -38072 41043 -38008
rect 40979 -38152 41043 -38088
rect 40979 -38232 41043 -38168
rect 40979 -38312 41043 -38248
rect 40979 -38392 41043 -38328
rect 40979 -38472 41043 -38408
rect 40979 -38552 41043 -38488
rect 40979 -38632 41043 -38568
rect 40979 -38712 41043 -38648
rect 40979 -38792 41043 -38728
rect 40979 -38872 41043 -38808
rect 40979 -38952 41043 -38888
rect 40979 -39032 41043 -38968
rect 40979 -39112 41043 -39048
rect 40979 -39192 41043 -39128
rect 40979 -39272 41043 -39208
rect 40979 -39352 41043 -39288
rect 40979 -39432 41043 -39368
rect 40979 -39512 41043 -39448
rect 40979 -39592 41043 -39528
rect 40979 -39672 41043 -39608
rect 40979 -39752 41043 -39688
rect 40979 -39832 41043 -39768
rect 40979 -39912 41043 -39848
rect 40979 -39992 41043 -39928
rect 40979 -40072 41043 -40008
rect 40979 -40152 41043 -40088
rect 40979 -40232 41043 -40168
rect 40979 -40312 41043 -40248
rect 40979 -40392 41043 -40328
rect 40979 -40472 41043 -40408
rect 40979 -40552 41043 -40488
rect 40979 -40632 41043 -40568
rect 40979 -40712 41043 -40648
rect 40979 -40792 41043 -40728
rect 40979 -40872 41043 -40808
rect 47298 -34792 47362 -34728
rect 47298 -34872 47362 -34808
rect 47298 -34952 47362 -34888
rect 47298 -35032 47362 -34968
rect 47298 -35112 47362 -35048
rect 47298 -35192 47362 -35128
rect 47298 -35272 47362 -35208
rect 47298 -35352 47362 -35288
rect 47298 -35432 47362 -35368
rect 47298 -35512 47362 -35448
rect 47298 -35592 47362 -35528
rect 47298 -35672 47362 -35608
rect 47298 -35752 47362 -35688
rect 47298 -35832 47362 -35768
rect 47298 -35912 47362 -35848
rect 47298 -35992 47362 -35928
rect 47298 -36072 47362 -36008
rect 47298 -36152 47362 -36088
rect 47298 -36232 47362 -36168
rect 47298 -36312 47362 -36248
rect 47298 -36392 47362 -36328
rect 47298 -36472 47362 -36408
rect 47298 -36552 47362 -36488
rect 47298 -36632 47362 -36568
rect 47298 -36712 47362 -36648
rect 47298 -36792 47362 -36728
rect 47298 -36872 47362 -36808
rect 47298 -36952 47362 -36888
rect 47298 -37032 47362 -36968
rect 47298 -37112 47362 -37048
rect 47298 -37192 47362 -37128
rect 47298 -37272 47362 -37208
rect 47298 -37352 47362 -37288
rect 47298 -37432 47362 -37368
rect 47298 -37512 47362 -37448
rect 47298 -37592 47362 -37528
rect 47298 -37672 47362 -37608
rect 47298 -37752 47362 -37688
rect 47298 -37832 47362 -37768
rect 47298 -37912 47362 -37848
rect 47298 -37992 47362 -37928
rect 47298 -38072 47362 -38008
rect 47298 -38152 47362 -38088
rect 47298 -38232 47362 -38168
rect 47298 -38312 47362 -38248
rect 47298 -38392 47362 -38328
rect 47298 -38472 47362 -38408
rect 47298 -38552 47362 -38488
rect 47298 -38632 47362 -38568
rect 47298 -38712 47362 -38648
rect 47298 -38792 47362 -38728
rect 47298 -38872 47362 -38808
rect 47298 -38952 47362 -38888
rect 47298 -39032 47362 -38968
rect 47298 -39112 47362 -39048
rect 47298 -39192 47362 -39128
rect 47298 -39272 47362 -39208
rect 47298 -39352 47362 -39288
rect 47298 -39432 47362 -39368
rect 47298 -39512 47362 -39448
rect 47298 -39592 47362 -39528
rect 47298 -39672 47362 -39608
rect 47298 -39752 47362 -39688
rect 47298 -39832 47362 -39768
rect 47298 -39912 47362 -39848
rect 47298 -39992 47362 -39928
rect 47298 -40072 47362 -40008
rect 47298 -40152 47362 -40088
rect 47298 -40232 47362 -40168
rect 47298 -40312 47362 -40248
rect 47298 -40392 47362 -40328
rect 47298 -40472 47362 -40408
rect 47298 -40552 47362 -40488
rect 47298 -40632 47362 -40568
rect 47298 -40712 47362 -40648
rect 47298 -40792 47362 -40728
rect 47298 -40872 47362 -40808
rect -41168 -41092 -41104 -41028
rect -41168 -41172 -41104 -41108
rect -41168 -41252 -41104 -41188
rect -41168 -41332 -41104 -41268
rect -41168 -41412 -41104 -41348
rect -41168 -41492 -41104 -41428
rect -41168 -41572 -41104 -41508
rect -41168 -41652 -41104 -41588
rect -41168 -41732 -41104 -41668
rect -41168 -41812 -41104 -41748
rect -41168 -41892 -41104 -41828
rect -41168 -41972 -41104 -41908
rect -41168 -42052 -41104 -41988
rect -41168 -42132 -41104 -42068
rect -41168 -42212 -41104 -42148
rect -41168 -42292 -41104 -42228
rect -41168 -42372 -41104 -42308
rect -41168 -42452 -41104 -42388
rect -41168 -42532 -41104 -42468
rect -41168 -42612 -41104 -42548
rect -41168 -42692 -41104 -42628
rect -41168 -42772 -41104 -42708
rect -41168 -42852 -41104 -42788
rect -41168 -42932 -41104 -42868
rect -41168 -43012 -41104 -42948
rect -41168 -43092 -41104 -43028
rect -41168 -43172 -41104 -43108
rect -41168 -43252 -41104 -43188
rect -41168 -43332 -41104 -43268
rect -41168 -43412 -41104 -43348
rect -41168 -43492 -41104 -43428
rect -41168 -43572 -41104 -43508
rect -41168 -43652 -41104 -43588
rect -41168 -43732 -41104 -43668
rect -41168 -43812 -41104 -43748
rect -41168 -43892 -41104 -43828
rect -41168 -43972 -41104 -43908
rect -41168 -44052 -41104 -43988
rect -41168 -44132 -41104 -44068
rect -41168 -44212 -41104 -44148
rect -41168 -44292 -41104 -44228
rect -41168 -44372 -41104 -44308
rect -41168 -44452 -41104 -44388
rect -41168 -44532 -41104 -44468
rect -41168 -44612 -41104 -44548
rect -41168 -44692 -41104 -44628
rect -41168 -44772 -41104 -44708
rect -41168 -44852 -41104 -44788
rect -41168 -44932 -41104 -44868
rect -41168 -45012 -41104 -44948
rect -41168 -45092 -41104 -45028
rect -41168 -45172 -41104 -45108
rect -41168 -45252 -41104 -45188
rect -41168 -45332 -41104 -45268
rect -41168 -45412 -41104 -45348
rect -41168 -45492 -41104 -45428
rect -41168 -45572 -41104 -45508
rect -41168 -45652 -41104 -45588
rect -41168 -45732 -41104 -45668
rect -41168 -45812 -41104 -45748
rect -41168 -45892 -41104 -45828
rect -41168 -45972 -41104 -45908
rect -41168 -46052 -41104 -45988
rect -41168 -46132 -41104 -46068
rect -41168 -46212 -41104 -46148
rect -41168 -46292 -41104 -46228
rect -41168 -46372 -41104 -46308
rect -41168 -46452 -41104 -46388
rect -41168 -46532 -41104 -46468
rect -41168 -46612 -41104 -46548
rect -41168 -46692 -41104 -46628
rect -41168 -46772 -41104 -46708
rect -41168 -46852 -41104 -46788
rect -41168 -46932 -41104 -46868
rect -41168 -47012 -41104 -46948
rect -41168 -47092 -41104 -47028
rect -41168 -47172 -41104 -47108
rect -34849 -41092 -34785 -41028
rect -34849 -41172 -34785 -41108
rect -34849 -41252 -34785 -41188
rect -34849 -41332 -34785 -41268
rect -34849 -41412 -34785 -41348
rect -34849 -41492 -34785 -41428
rect -34849 -41572 -34785 -41508
rect -34849 -41652 -34785 -41588
rect -34849 -41732 -34785 -41668
rect -34849 -41812 -34785 -41748
rect -34849 -41892 -34785 -41828
rect -34849 -41972 -34785 -41908
rect -34849 -42052 -34785 -41988
rect -34849 -42132 -34785 -42068
rect -34849 -42212 -34785 -42148
rect -34849 -42292 -34785 -42228
rect -34849 -42372 -34785 -42308
rect -34849 -42452 -34785 -42388
rect -34849 -42532 -34785 -42468
rect -34849 -42612 -34785 -42548
rect -34849 -42692 -34785 -42628
rect -34849 -42772 -34785 -42708
rect -34849 -42852 -34785 -42788
rect -34849 -42932 -34785 -42868
rect -34849 -43012 -34785 -42948
rect -34849 -43092 -34785 -43028
rect -34849 -43172 -34785 -43108
rect -34849 -43252 -34785 -43188
rect -34849 -43332 -34785 -43268
rect -34849 -43412 -34785 -43348
rect -34849 -43492 -34785 -43428
rect -34849 -43572 -34785 -43508
rect -34849 -43652 -34785 -43588
rect -34849 -43732 -34785 -43668
rect -34849 -43812 -34785 -43748
rect -34849 -43892 -34785 -43828
rect -34849 -43972 -34785 -43908
rect -34849 -44052 -34785 -43988
rect -34849 -44132 -34785 -44068
rect -34849 -44212 -34785 -44148
rect -34849 -44292 -34785 -44228
rect -34849 -44372 -34785 -44308
rect -34849 -44452 -34785 -44388
rect -34849 -44532 -34785 -44468
rect -34849 -44612 -34785 -44548
rect -34849 -44692 -34785 -44628
rect -34849 -44772 -34785 -44708
rect -34849 -44852 -34785 -44788
rect -34849 -44932 -34785 -44868
rect -34849 -45012 -34785 -44948
rect -34849 -45092 -34785 -45028
rect -34849 -45172 -34785 -45108
rect -34849 -45252 -34785 -45188
rect -34849 -45332 -34785 -45268
rect -34849 -45412 -34785 -45348
rect -34849 -45492 -34785 -45428
rect -34849 -45572 -34785 -45508
rect -34849 -45652 -34785 -45588
rect -34849 -45732 -34785 -45668
rect -34849 -45812 -34785 -45748
rect -34849 -45892 -34785 -45828
rect -34849 -45972 -34785 -45908
rect -34849 -46052 -34785 -45988
rect -34849 -46132 -34785 -46068
rect -34849 -46212 -34785 -46148
rect -34849 -46292 -34785 -46228
rect -34849 -46372 -34785 -46308
rect -34849 -46452 -34785 -46388
rect -34849 -46532 -34785 -46468
rect -34849 -46612 -34785 -46548
rect -34849 -46692 -34785 -46628
rect -34849 -46772 -34785 -46708
rect -34849 -46852 -34785 -46788
rect -34849 -46932 -34785 -46868
rect -34849 -47012 -34785 -46948
rect -34849 -47092 -34785 -47028
rect -34849 -47172 -34785 -47108
rect -28530 -41092 -28466 -41028
rect -28530 -41172 -28466 -41108
rect -28530 -41252 -28466 -41188
rect -28530 -41332 -28466 -41268
rect -28530 -41412 -28466 -41348
rect -28530 -41492 -28466 -41428
rect -28530 -41572 -28466 -41508
rect -28530 -41652 -28466 -41588
rect -28530 -41732 -28466 -41668
rect -28530 -41812 -28466 -41748
rect -28530 -41892 -28466 -41828
rect -28530 -41972 -28466 -41908
rect -28530 -42052 -28466 -41988
rect -28530 -42132 -28466 -42068
rect -28530 -42212 -28466 -42148
rect -28530 -42292 -28466 -42228
rect -28530 -42372 -28466 -42308
rect -28530 -42452 -28466 -42388
rect -28530 -42532 -28466 -42468
rect -28530 -42612 -28466 -42548
rect -28530 -42692 -28466 -42628
rect -28530 -42772 -28466 -42708
rect -28530 -42852 -28466 -42788
rect -28530 -42932 -28466 -42868
rect -28530 -43012 -28466 -42948
rect -28530 -43092 -28466 -43028
rect -28530 -43172 -28466 -43108
rect -28530 -43252 -28466 -43188
rect -28530 -43332 -28466 -43268
rect -28530 -43412 -28466 -43348
rect -28530 -43492 -28466 -43428
rect -28530 -43572 -28466 -43508
rect -28530 -43652 -28466 -43588
rect -28530 -43732 -28466 -43668
rect -28530 -43812 -28466 -43748
rect -28530 -43892 -28466 -43828
rect -28530 -43972 -28466 -43908
rect -28530 -44052 -28466 -43988
rect -28530 -44132 -28466 -44068
rect -28530 -44212 -28466 -44148
rect -28530 -44292 -28466 -44228
rect -28530 -44372 -28466 -44308
rect -28530 -44452 -28466 -44388
rect -28530 -44532 -28466 -44468
rect -28530 -44612 -28466 -44548
rect -28530 -44692 -28466 -44628
rect -28530 -44772 -28466 -44708
rect -28530 -44852 -28466 -44788
rect -28530 -44932 -28466 -44868
rect -28530 -45012 -28466 -44948
rect -28530 -45092 -28466 -45028
rect -28530 -45172 -28466 -45108
rect -28530 -45252 -28466 -45188
rect -28530 -45332 -28466 -45268
rect -28530 -45412 -28466 -45348
rect -28530 -45492 -28466 -45428
rect -28530 -45572 -28466 -45508
rect -28530 -45652 -28466 -45588
rect -28530 -45732 -28466 -45668
rect -28530 -45812 -28466 -45748
rect -28530 -45892 -28466 -45828
rect -28530 -45972 -28466 -45908
rect -28530 -46052 -28466 -45988
rect -28530 -46132 -28466 -46068
rect -28530 -46212 -28466 -46148
rect -28530 -46292 -28466 -46228
rect -28530 -46372 -28466 -46308
rect -28530 -46452 -28466 -46388
rect -28530 -46532 -28466 -46468
rect -28530 -46612 -28466 -46548
rect -28530 -46692 -28466 -46628
rect -28530 -46772 -28466 -46708
rect -28530 -46852 -28466 -46788
rect -28530 -46932 -28466 -46868
rect -28530 -47012 -28466 -46948
rect -28530 -47092 -28466 -47028
rect -28530 -47172 -28466 -47108
rect -22211 -41092 -22147 -41028
rect -22211 -41172 -22147 -41108
rect -22211 -41252 -22147 -41188
rect -22211 -41332 -22147 -41268
rect -22211 -41412 -22147 -41348
rect -22211 -41492 -22147 -41428
rect -22211 -41572 -22147 -41508
rect -22211 -41652 -22147 -41588
rect -22211 -41732 -22147 -41668
rect -22211 -41812 -22147 -41748
rect -22211 -41892 -22147 -41828
rect -22211 -41972 -22147 -41908
rect -22211 -42052 -22147 -41988
rect -22211 -42132 -22147 -42068
rect -22211 -42212 -22147 -42148
rect -22211 -42292 -22147 -42228
rect -22211 -42372 -22147 -42308
rect -22211 -42452 -22147 -42388
rect -22211 -42532 -22147 -42468
rect -22211 -42612 -22147 -42548
rect -22211 -42692 -22147 -42628
rect -22211 -42772 -22147 -42708
rect -22211 -42852 -22147 -42788
rect -22211 -42932 -22147 -42868
rect -22211 -43012 -22147 -42948
rect -22211 -43092 -22147 -43028
rect -22211 -43172 -22147 -43108
rect -22211 -43252 -22147 -43188
rect -22211 -43332 -22147 -43268
rect -22211 -43412 -22147 -43348
rect -22211 -43492 -22147 -43428
rect -22211 -43572 -22147 -43508
rect -22211 -43652 -22147 -43588
rect -22211 -43732 -22147 -43668
rect -22211 -43812 -22147 -43748
rect -22211 -43892 -22147 -43828
rect -22211 -43972 -22147 -43908
rect -22211 -44052 -22147 -43988
rect -22211 -44132 -22147 -44068
rect -22211 -44212 -22147 -44148
rect -22211 -44292 -22147 -44228
rect -22211 -44372 -22147 -44308
rect -22211 -44452 -22147 -44388
rect -22211 -44532 -22147 -44468
rect -22211 -44612 -22147 -44548
rect -22211 -44692 -22147 -44628
rect -22211 -44772 -22147 -44708
rect -22211 -44852 -22147 -44788
rect -22211 -44932 -22147 -44868
rect -22211 -45012 -22147 -44948
rect -22211 -45092 -22147 -45028
rect -22211 -45172 -22147 -45108
rect -22211 -45252 -22147 -45188
rect -22211 -45332 -22147 -45268
rect -22211 -45412 -22147 -45348
rect -22211 -45492 -22147 -45428
rect -22211 -45572 -22147 -45508
rect -22211 -45652 -22147 -45588
rect -22211 -45732 -22147 -45668
rect -22211 -45812 -22147 -45748
rect -22211 -45892 -22147 -45828
rect -22211 -45972 -22147 -45908
rect -22211 -46052 -22147 -45988
rect -22211 -46132 -22147 -46068
rect -22211 -46212 -22147 -46148
rect -22211 -46292 -22147 -46228
rect -22211 -46372 -22147 -46308
rect -22211 -46452 -22147 -46388
rect -22211 -46532 -22147 -46468
rect -22211 -46612 -22147 -46548
rect -22211 -46692 -22147 -46628
rect -22211 -46772 -22147 -46708
rect -22211 -46852 -22147 -46788
rect -22211 -46932 -22147 -46868
rect -22211 -47012 -22147 -46948
rect -22211 -47092 -22147 -47028
rect -22211 -47172 -22147 -47108
rect -15892 -41092 -15828 -41028
rect -15892 -41172 -15828 -41108
rect -15892 -41252 -15828 -41188
rect -15892 -41332 -15828 -41268
rect -15892 -41412 -15828 -41348
rect -15892 -41492 -15828 -41428
rect -15892 -41572 -15828 -41508
rect -15892 -41652 -15828 -41588
rect -15892 -41732 -15828 -41668
rect -15892 -41812 -15828 -41748
rect -15892 -41892 -15828 -41828
rect -15892 -41972 -15828 -41908
rect -15892 -42052 -15828 -41988
rect -15892 -42132 -15828 -42068
rect -15892 -42212 -15828 -42148
rect -15892 -42292 -15828 -42228
rect -15892 -42372 -15828 -42308
rect -15892 -42452 -15828 -42388
rect -15892 -42532 -15828 -42468
rect -15892 -42612 -15828 -42548
rect -15892 -42692 -15828 -42628
rect -15892 -42772 -15828 -42708
rect -15892 -42852 -15828 -42788
rect -15892 -42932 -15828 -42868
rect -15892 -43012 -15828 -42948
rect -15892 -43092 -15828 -43028
rect -15892 -43172 -15828 -43108
rect -15892 -43252 -15828 -43188
rect -15892 -43332 -15828 -43268
rect -15892 -43412 -15828 -43348
rect -15892 -43492 -15828 -43428
rect -15892 -43572 -15828 -43508
rect -15892 -43652 -15828 -43588
rect -15892 -43732 -15828 -43668
rect -15892 -43812 -15828 -43748
rect -15892 -43892 -15828 -43828
rect -15892 -43972 -15828 -43908
rect -15892 -44052 -15828 -43988
rect -15892 -44132 -15828 -44068
rect -15892 -44212 -15828 -44148
rect -15892 -44292 -15828 -44228
rect -15892 -44372 -15828 -44308
rect -15892 -44452 -15828 -44388
rect -15892 -44532 -15828 -44468
rect -15892 -44612 -15828 -44548
rect -15892 -44692 -15828 -44628
rect -15892 -44772 -15828 -44708
rect -15892 -44852 -15828 -44788
rect -15892 -44932 -15828 -44868
rect -15892 -45012 -15828 -44948
rect -15892 -45092 -15828 -45028
rect -15892 -45172 -15828 -45108
rect -15892 -45252 -15828 -45188
rect -15892 -45332 -15828 -45268
rect -15892 -45412 -15828 -45348
rect -15892 -45492 -15828 -45428
rect -15892 -45572 -15828 -45508
rect -15892 -45652 -15828 -45588
rect -15892 -45732 -15828 -45668
rect -15892 -45812 -15828 -45748
rect -15892 -45892 -15828 -45828
rect -15892 -45972 -15828 -45908
rect -15892 -46052 -15828 -45988
rect -15892 -46132 -15828 -46068
rect -15892 -46212 -15828 -46148
rect -15892 -46292 -15828 -46228
rect -15892 -46372 -15828 -46308
rect -15892 -46452 -15828 -46388
rect -15892 -46532 -15828 -46468
rect -15892 -46612 -15828 -46548
rect -15892 -46692 -15828 -46628
rect -15892 -46772 -15828 -46708
rect -15892 -46852 -15828 -46788
rect -15892 -46932 -15828 -46868
rect -15892 -47012 -15828 -46948
rect -15892 -47092 -15828 -47028
rect -15892 -47172 -15828 -47108
rect -9573 -41092 -9509 -41028
rect -9573 -41172 -9509 -41108
rect -9573 -41252 -9509 -41188
rect -9573 -41332 -9509 -41268
rect -9573 -41412 -9509 -41348
rect -9573 -41492 -9509 -41428
rect -9573 -41572 -9509 -41508
rect -9573 -41652 -9509 -41588
rect -9573 -41732 -9509 -41668
rect -9573 -41812 -9509 -41748
rect -9573 -41892 -9509 -41828
rect -9573 -41972 -9509 -41908
rect -9573 -42052 -9509 -41988
rect -9573 -42132 -9509 -42068
rect -9573 -42212 -9509 -42148
rect -9573 -42292 -9509 -42228
rect -9573 -42372 -9509 -42308
rect -9573 -42452 -9509 -42388
rect -9573 -42532 -9509 -42468
rect -9573 -42612 -9509 -42548
rect -9573 -42692 -9509 -42628
rect -9573 -42772 -9509 -42708
rect -9573 -42852 -9509 -42788
rect -9573 -42932 -9509 -42868
rect -9573 -43012 -9509 -42948
rect -9573 -43092 -9509 -43028
rect -9573 -43172 -9509 -43108
rect -9573 -43252 -9509 -43188
rect -9573 -43332 -9509 -43268
rect -9573 -43412 -9509 -43348
rect -9573 -43492 -9509 -43428
rect -9573 -43572 -9509 -43508
rect -9573 -43652 -9509 -43588
rect -9573 -43732 -9509 -43668
rect -9573 -43812 -9509 -43748
rect -9573 -43892 -9509 -43828
rect -9573 -43972 -9509 -43908
rect -9573 -44052 -9509 -43988
rect -9573 -44132 -9509 -44068
rect -9573 -44212 -9509 -44148
rect -9573 -44292 -9509 -44228
rect -9573 -44372 -9509 -44308
rect -9573 -44452 -9509 -44388
rect -9573 -44532 -9509 -44468
rect -9573 -44612 -9509 -44548
rect -9573 -44692 -9509 -44628
rect -9573 -44772 -9509 -44708
rect -9573 -44852 -9509 -44788
rect -9573 -44932 -9509 -44868
rect -9573 -45012 -9509 -44948
rect -9573 -45092 -9509 -45028
rect -9573 -45172 -9509 -45108
rect -9573 -45252 -9509 -45188
rect -9573 -45332 -9509 -45268
rect -9573 -45412 -9509 -45348
rect -9573 -45492 -9509 -45428
rect -9573 -45572 -9509 -45508
rect -9573 -45652 -9509 -45588
rect -9573 -45732 -9509 -45668
rect -9573 -45812 -9509 -45748
rect -9573 -45892 -9509 -45828
rect -9573 -45972 -9509 -45908
rect -9573 -46052 -9509 -45988
rect -9573 -46132 -9509 -46068
rect -9573 -46212 -9509 -46148
rect -9573 -46292 -9509 -46228
rect -9573 -46372 -9509 -46308
rect -9573 -46452 -9509 -46388
rect -9573 -46532 -9509 -46468
rect -9573 -46612 -9509 -46548
rect -9573 -46692 -9509 -46628
rect -9573 -46772 -9509 -46708
rect -9573 -46852 -9509 -46788
rect -9573 -46932 -9509 -46868
rect -9573 -47012 -9509 -46948
rect -9573 -47092 -9509 -47028
rect -9573 -47172 -9509 -47108
rect -3254 -41092 -3190 -41028
rect -3254 -41172 -3190 -41108
rect -3254 -41252 -3190 -41188
rect -3254 -41332 -3190 -41268
rect -3254 -41412 -3190 -41348
rect -3254 -41492 -3190 -41428
rect -3254 -41572 -3190 -41508
rect -3254 -41652 -3190 -41588
rect -3254 -41732 -3190 -41668
rect -3254 -41812 -3190 -41748
rect -3254 -41892 -3190 -41828
rect -3254 -41972 -3190 -41908
rect -3254 -42052 -3190 -41988
rect -3254 -42132 -3190 -42068
rect -3254 -42212 -3190 -42148
rect -3254 -42292 -3190 -42228
rect -3254 -42372 -3190 -42308
rect -3254 -42452 -3190 -42388
rect -3254 -42532 -3190 -42468
rect -3254 -42612 -3190 -42548
rect -3254 -42692 -3190 -42628
rect -3254 -42772 -3190 -42708
rect -3254 -42852 -3190 -42788
rect -3254 -42932 -3190 -42868
rect -3254 -43012 -3190 -42948
rect -3254 -43092 -3190 -43028
rect -3254 -43172 -3190 -43108
rect -3254 -43252 -3190 -43188
rect -3254 -43332 -3190 -43268
rect -3254 -43412 -3190 -43348
rect -3254 -43492 -3190 -43428
rect -3254 -43572 -3190 -43508
rect -3254 -43652 -3190 -43588
rect -3254 -43732 -3190 -43668
rect -3254 -43812 -3190 -43748
rect -3254 -43892 -3190 -43828
rect -3254 -43972 -3190 -43908
rect -3254 -44052 -3190 -43988
rect -3254 -44132 -3190 -44068
rect -3254 -44212 -3190 -44148
rect -3254 -44292 -3190 -44228
rect -3254 -44372 -3190 -44308
rect -3254 -44452 -3190 -44388
rect -3254 -44532 -3190 -44468
rect -3254 -44612 -3190 -44548
rect -3254 -44692 -3190 -44628
rect -3254 -44772 -3190 -44708
rect -3254 -44852 -3190 -44788
rect -3254 -44932 -3190 -44868
rect -3254 -45012 -3190 -44948
rect -3254 -45092 -3190 -45028
rect -3254 -45172 -3190 -45108
rect -3254 -45252 -3190 -45188
rect -3254 -45332 -3190 -45268
rect -3254 -45412 -3190 -45348
rect -3254 -45492 -3190 -45428
rect -3254 -45572 -3190 -45508
rect -3254 -45652 -3190 -45588
rect -3254 -45732 -3190 -45668
rect -3254 -45812 -3190 -45748
rect -3254 -45892 -3190 -45828
rect -3254 -45972 -3190 -45908
rect -3254 -46052 -3190 -45988
rect -3254 -46132 -3190 -46068
rect -3254 -46212 -3190 -46148
rect -3254 -46292 -3190 -46228
rect -3254 -46372 -3190 -46308
rect -3254 -46452 -3190 -46388
rect -3254 -46532 -3190 -46468
rect -3254 -46612 -3190 -46548
rect -3254 -46692 -3190 -46628
rect -3254 -46772 -3190 -46708
rect -3254 -46852 -3190 -46788
rect -3254 -46932 -3190 -46868
rect -3254 -47012 -3190 -46948
rect -3254 -47092 -3190 -47028
rect -3254 -47172 -3190 -47108
rect 3065 -41092 3129 -41028
rect 3065 -41172 3129 -41108
rect 3065 -41252 3129 -41188
rect 3065 -41332 3129 -41268
rect 3065 -41412 3129 -41348
rect 3065 -41492 3129 -41428
rect 3065 -41572 3129 -41508
rect 3065 -41652 3129 -41588
rect 3065 -41732 3129 -41668
rect 3065 -41812 3129 -41748
rect 3065 -41892 3129 -41828
rect 3065 -41972 3129 -41908
rect 3065 -42052 3129 -41988
rect 3065 -42132 3129 -42068
rect 3065 -42212 3129 -42148
rect 3065 -42292 3129 -42228
rect 3065 -42372 3129 -42308
rect 3065 -42452 3129 -42388
rect 3065 -42532 3129 -42468
rect 3065 -42612 3129 -42548
rect 3065 -42692 3129 -42628
rect 3065 -42772 3129 -42708
rect 3065 -42852 3129 -42788
rect 3065 -42932 3129 -42868
rect 3065 -43012 3129 -42948
rect 3065 -43092 3129 -43028
rect 3065 -43172 3129 -43108
rect 3065 -43252 3129 -43188
rect 3065 -43332 3129 -43268
rect 3065 -43412 3129 -43348
rect 3065 -43492 3129 -43428
rect 3065 -43572 3129 -43508
rect 3065 -43652 3129 -43588
rect 3065 -43732 3129 -43668
rect 3065 -43812 3129 -43748
rect 3065 -43892 3129 -43828
rect 3065 -43972 3129 -43908
rect 3065 -44052 3129 -43988
rect 3065 -44132 3129 -44068
rect 3065 -44212 3129 -44148
rect 3065 -44292 3129 -44228
rect 3065 -44372 3129 -44308
rect 3065 -44452 3129 -44388
rect 3065 -44532 3129 -44468
rect 3065 -44612 3129 -44548
rect 3065 -44692 3129 -44628
rect 3065 -44772 3129 -44708
rect 3065 -44852 3129 -44788
rect 3065 -44932 3129 -44868
rect 3065 -45012 3129 -44948
rect 3065 -45092 3129 -45028
rect 3065 -45172 3129 -45108
rect 3065 -45252 3129 -45188
rect 3065 -45332 3129 -45268
rect 3065 -45412 3129 -45348
rect 3065 -45492 3129 -45428
rect 3065 -45572 3129 -45508
rect 3065 -45652 3129 -45588
rect 3065 -45732 3129 -45668
rect 3065 -45812 3129 -45748
rect 3065 -45892 3129 -45828
rect 3065 -45972 3129 -45908
rect 3065 -46052 3129 -45988
rect 3065 -46132 3129 -46068
rect 3065 -46212 3129 -46148
rect 3065 -46292 3129 -46228
rect 3065 -46372 3129 -46308
rect 3065 -46452 3129 -46388
rect 3065 -46532 3129 -46468
rect 3065 -46612 3129 -46548
rect 3065 -46692 3129 -46628
rect 3065 -46772 3129 -46708
rect 3065 -46852 3129 -46788
rect 3065 -46932 3129 -46868
rect 3065 -47012 3129 -46948
rect 3065 -47092 3129 -47028
rect 3065 -47172 3129 -47108
rect 9384 -41092 9448 -41028
rect 9384 -41172 9448 -41108
rect 9384 -41252 9448 -41188
rect 9384 -41332 9448 -41268
rect 9384 -41412 9448 -41348
rect 9384 -41492 9448 -41428
rect 9384 -41572 9448 -41508
rect 9384 -41652 9448 -41588
rect 9384 -41732 9448 -41668
rect 9384 -41812 9448 -41748
rect 9384 -41892 9448 -41828
rect 9384 -41972 9448 -41908
rect 9384 -42052 9448 -41988
rect 9384 -42132 9448 -42068
rect 9384 -42212 9448 -42148
rect 9384 -42292 9448 -42228
rect 9384 -42372 9448 -42308
rect 9384 -42452 9448 -42388
rect 9384 -42532 9448 -42468
rect 9384 -42612 9448 -42548
rect 9384 -42692 9448 -42628
rect 9384 -42772 9448 -42708
rect 9384 -42852 9448 -42788
rect 9384 -42932 9448 -42868
rect 9384 -43012 9448 -42948
rect 9384 -43092 9448 -43028
rect 9384 -43172 9448 -43108
rect 9384 -43252 9448 -43188
rect 9384 -43332 9448 -43268
rect 9384 -43412 9448 -43348
rect 9384 -43492 9448 -43428
rect 9384 -43572 9448 -43508
rect 9384 -43652 9448 -43588
rect 9384 -43732 9448 -43668
rect 9384 -43812 9448 -43748
rect 9384 -43892 9448 -43828
rect 9384 -43972 9448 -43908
rect 9384 -44052 9448 -43988
rect 9384 -44132 9448 -44068
rect 9384 -44212 9448 -44148
rect 9384 -44292 9448 -44228
rect 9384 -44372 9448 -44308
rect 9384 -44452 9448 -44388
rect 9384 -44532 9448 -44468
rect 9384 -44612 9448 -44548
rect 9384 -44692 9448 -44628
rect 9384 -44772 9448 -44708
rect 9384 -44852 9448 -44788
rect 9384 -44932 9448 -44868
rect 9384 -45012 9448 -44948
rect 9384 -45092 9448 -45028
rect 9384 -45172 9448 -45108
rect 9384 -45252 9448 -45188
rect 9384 -45332 9448 -45268
rect 9384 -45412 9448 -45348
rect 9384 -45492 9448 -45428
rect 9384 -45572 9448 -45508
rect 9384 -45652 9448 -45588
rect 9384 -45732 9448 -45668
rect 9384 -45812 9448 -45748
rect 9384 -45892 9448 -45828
rect 9384 -45972 9448 -45908
rect 9384 -46052 9448 -45988
rect 9384 -46132 9448 -46068
rect 9384 -46212 9448 -46148
rect 9384 -46292 9448 -46228
rect 9384 -46372 9448 -46308
rect 9384 -46452 9448 -46388
rect 9384 -46532 9448 -46468
rect 9384 -46612 9448 -46548
rect 9384 -46692 9448 -46628
rect 9384 -46772 9448 -46708
rect 9384 -46852 9448 -46788
rect 9384 -46932 9448 -46868
rect 9384 -47012 9448 -46948
rect 9384 -47092 9448 -47028
rect 9384 -47172 9448 -47108
rect 15703 -41092 15767 -41028
rect 15703 -41172 15767 -41108
rect 15703 -41252 15767 -41188
rect 15703 -41332 15767 -41268
rect 15703 -41412 15767 -41348
rect 15703 -41492 15767 -41428
rect 15703 -41572 15767 -41508
rect 15703 -41652 15767 -41588
rect 15703 -41732 15767 -41668
rect 15703 -41812 15767 -41748
rect 15703 -41892 15767 -41828
rect 15703 -41972 15767 -41908
rect 15703 -42052 15767 -41988
rect 15703 -42132 15767 -42068
rect 15703 -42212 15767 -42148
rect 15703 -42292 15767 -42228
rect 15703 -42372 15767 -42308
rect 15703 -42452 15767 -42388
rect 15703 -42532 15767 -42468
rect 15703 -42612 15767 -42548
rect 15703 -42692 15767 -42628
rect 15703 -42772 15767 -42708
rect 15703 -42852 15767 -42788
rect 15703 -42932 15767 -42868
rect 15703 -43012 15767 -42948
rect 15703 -43092 15767 -43028
rect 15703 -43172 15767 -43108
rect 15703 -43252 15767 -43188
rect 15703 -43332 15767 -43268
rect 15703 -43412 15767 -43348
rect 15703 -43492 15767 -43428
rect 15703 -43572 15767 -43508
rect 15703 -43652 15767 -43588
rect 15703 -43732 15767 -43668
rect 15703 -43812 15767 -43748
rect 15703 -43892 15767 -43828
rect 15703 -43972 15767 -43908
rect 15703 -44052 15767 -43988
rect 15703 -44132 15767 -44068
rect 15703 -44212 15767 -44148
rect 15703 -44292 15767 -44228
rect 15703 -44372 15767 -44308
rect 15703 -44452 15767 -44388
rect 15703 -44532 15767 -44468
rect 15703 -44612 15767 -44548
rect 15703 -44692 15767 -44628
rect 15703 -44772 15767 -44708
rect 15703 -44852 15767 -44788
rect 15703 -44932 15767 -44868
rect 15703 -45012 15767 -44948
rect 15703 -45092 15767 -45028
rect 15703 -45172 15767 -45108
rect 15703 -45252 15767 -45188
rect 15703 -45332 15767 -45268
rect 15703 -45412 15767 -45348
rect 15703 -45492 15767 -45428
rect 15703 -45572 15767 -45508
rect 15703 -45652 15767 -45588
rect 15703 -45732 15767 -45668
rect 15703 -45812 15767 -45748
rect 15703 -45892 15767 -45828
rect 15703 -45972 15767 -45908
rect 15703 -46052 15767 -45988
rect 15703 -46132 15767 -46068
rect 15703 -46212 15767 -46148
rect 15703 -46292 15767 -46228
rect 15703 -46372 15767 -46308
rect 15703 -46452 15767 -46388
rect 15703 -46532 15767 -46468
rect 15703 -46612 15767 -46548
rect 15703 -46692 15767 -46628
rect 15703 -46772 15767 -46708
rect 15703 -46852 15767 -46788
rect 15703 -46932 15767 -46868
rect 15703 -47012 15767 -46948
rect 15703 -47092 15767 -47028
rect 15703 -47172 15767 -47108
rect 22022 -41092 22086 -41028
rect 22022 -41172 22086 -41108
rect 22022 -41252 22086 -41188
rect 22022 -41332 22086 -41268
rect 22022 -41412 22086 -41348
rect 22022 -41492 22086 -41428
rect 22022 -41572 22086 -41508
rect 22022 -41652 22086 -41588
rect 22022 -41732 22086 -41668
rect 22022 -41812 22086 -41748
rect 22022 -41892 22086 -41828
rect 22022 -41972 22086 -41908
rect 22022 -42052 22086 -41988
rect 22022 -42132 22086 -42068
rect 22022 -42212 22086 -42148
rect 22022 -42292 22086 -42228
rect 22022 -42372 22086 -42308
rect 22022 -42452 22086 -42388
rect 22022 -42532 22086 -42468
rect 22022 -42612 22086 -42548
rect 22022 -42692 22086 -42628
rect 22022 -42772 22086 -42708
rect 22022 -42852 22086 -42788
rect 22022 -42932 22086 -42868
rect 22022 -43012 22086 -42948
rect 22022 -43092 22086 -43028
rect 22022 -43172 22086 -43108
rect 22022 -43252 22086 -43188
rect 22022 -43332 22086 -43268
rect 22022 -43412 22086 -43348
rect 22022 -43492 22086 -43428
rect 22022 -43572 22086 -43508
rect 22022 -43652 22086 -43588
rect 22022 -43732 22086 -43668
rect 22022 -43812 22086 -43748
rect 22022 -43892 22086 -43828
rect 22022 -43972 22086 -43908
rect 22022 -44052 22086 -43988
rect 22022 -44132 22086 -44068
rect 22022 -44212 22086 -44148
rect 22022 -44292 22086 -44228
rect 22022 -44372 22086 -44308
rect 22022 -44452 22086 -44388
rect 22022 -44532 22086 -44468
rect 22022 -44612 22086 -44548
rect 22022 -44692 22086 -44628
rect 22022 -44772 22086 -44708
rect 22022 -44852 22086 -44788
rect 22022 -44932 22086 -44868
rect 22022 -45012 22086 -44948
rect 22022 -45092 22086 -45028
rect 22022 -45172 22086 -45108
rect 22022 -45252 22086 -45188
rect 22022 -45332 22086 -45268
rect 22022 -45412 22086 -45348
rect 22022 -45492 22086 -45428
rect 22022 -45572 22086 -45508
rect 22022 -45652 22086 -45588
rect 22022 -45732 22086 -45668
rect 22022 -45812 22086 -45748
rect 22022 -45892 22086 -45828
rect 22022 -45972 22086 -45908
rect 22022 -46052 22086 -45988
rect 22022 -46132 22086 -46068
rect 22022 -46212 22086 -46148
rect 22022 -46292 22086 -46228
rect 22022 -46372 22086 -46308
rect 22022 -46452 22086 -46388
rect 22022 -46532 22086 -46468
rect 22022 -46612 22086 -46548
rect 22022 -46692 22086 -46628
rect 22022 -46772 22086 -46708
rect 22022 -46852 22086 -46788
rect 22022 -46932 22086 -46868
rect 22022 -47012 22086 -46948
rect 22022 -47092 22086 -47028
rect 22022 -47172 22086 -47108
rect 28341 -41092 28405 -41028
rect 28341 -41172 28405 -41108
rect 28341 -41252 28405 -41188
rect 28341 -41332 28405 -41268
rect 28341 -41412 28405 -41348
rect 28341 -41492 28405 -41428
rect 28341 -41572 28405 -41508
rect 28341 -41652 28405 -41588
rect 28341 -41732 28405 -41668
rect 28341 -41812 28405 -41748
rect 28341 -41892 28405 -41828
rect 28341 -41972 28405 -41908
rect 28341 -42052 28405 -41988
rect 28341 -42132 28405 -42068
rect 28341 -42212 28405 -42148
rect 28341 -42292 28405 -42228
rect 28341 -42372 28405 -42308
rect 28341 -42452 28405 -42388
rect 28341 -42532 28405 -42468
rect 28341 -42612 28405 -42548
rect 28341 -42692 28405 -42628
rect 28341 -42772 28405 -42708
rect 28341 -42852 28405 -42788
rect 28341 -42932 28405 -42868
rect 28341 -43012 28405 -42948
rect 28341 -43092 28405 -43028
rect 28341 -43172 28405 -43108
rect 28341 -43252 28405 -43188
rect 28341 -43332 28405 -43268
rect 28341 -43412 28405 -43348
rect 28341 -43492 28405 -43428
rect 28341 -43572 28405 -43508
rect 28341 -43652 28405 -43588
rect 28341 -43732 28405 -43668
rect 28341 -43812 28405 -43748
rect 28341 -43892 28405 -43828
rect 28341 -43972 28405 -43908
rect 28341 -44052 28405 -43988
rect 28341 -44132 28405 -44068
rect 28341 -44212 28405 -44148
rect 28341 -44292 28405 -44228
rect 28341 -44372 28405 -44308
rect 28341 -44452 28405 -44388
rect 28341 -44532 28405 -44468
rect 28341 -44612 28405 -44548
rect 28341 -44692 28405 -44628
rect 28341 -44772 28405 -44708
rect 28341 -44852 28405 -44788
rect 28341 -44932 28405 -44868
rect 28341 -45012 28405 -44948
rect 28341 -45092 28405 -45028
rect 28341 -45172 28405 -45108
rect 28341 -45252 28405 -45188
rect 28341 -45332 28405 -45268
rect 28341 -45412 28405 -45348
rect 28341 -45492 28405 -45428
rect 28341 -45572 28405 -45508
rect 28341 -45652 28405 -45588
rect 28341 -45732 28405 -45668
rect 28341 -45812 28405 -45748
rect 28341 -45892 28405 -45828
rect 28341 -45972 28405 -45908
rect 28341 -46052 28405 -45988
rect 28341 -46132 28405 -46068
rect 28341 -46212 28405 -46148
rect 28341 -46292 28405 -46228
rect 28341 -46372 28405 -46308
rect 28341 -46452 28405 -46388
rect 28341 -46532 28405 -46468
rect 28341 -46612 28405 -46548
rect 28341 -46692 28405 -46628
rect 28341 -46772 28405 -46708
rect 28341 -46852 28405 -46788
rect 28341 -46932 28405 -46868
rect 28341 -47012 28405 -46948
rect 28341 -47092 28405 -47028
rect 28341 -47172 28405 -47108
rect 34660 -41092 34724 -41028
rect 34660 -41172 34724 -41108
rect 34660 -41252 34724 -41188
rect 34660 -41332 34724 -41268
rect 34660 -41412 34724 -41348
rect 34660 -41492 34724 -41428
rect 34660 -41572 34724 -41508
rect 34660 -41652 34724 -41588
rect 34660 -41732 34724 -41668
rect 34660 -41812 34724 -41748
rect 34660 -41892 34724 -41828
rect 34660 -41972 34724 -41908
rect 34660 -42052 34724 -41988
rect 34660 -42132 34724 -42068
rect 34660 -42212 34724 -42148
rect 34660 -42292 34724 -42228
rect 34660 -42372 34724 -42308
rect 34660 -42452 34724 -42388
rect 34660 -42532 34724 -42468
rect 34660 -42612 34724 -42548
rect 34660 -42692 34724 -42628
rect 34660 -42772 34724 -42708
rect 34660 -42852 34724 -42788
rect 34660 -42932 34724 -42868
rect 34660 -43012 34724 -42948
rect 34660 -43092 34724 -43028
rect 34660 -43172 34724 -43108
rect 34660 -43252 34724 -43188
rect 34660 -43332 34724 -43268
rect 34660 -43412 34724 -43348
rect 34660 -43492 34724 -43428
rect 34660 -43572 34724 -43508
rect 34660 -43652 34724 -43588
rect 34660 -43732 34724 -43668
rect 34660 -43812 34724 -43748
rect 34660 -43892 34724 -43828
rect 34660 -43972 34724 -43908
rect 34660 -44052 34724 -43988
rect 34660 -44132 34724 -44068
rect 34660 -44212 34724 -44148
rect 34660 -44292 34724 -44228
rect 34660 -44372 34724 -44308
rect 34660 -44452 34724 -44388
rect 34660 -44532 34724 -44468
rect 34660 -44612 34724 -44548
rect 34660 -44692 34724 -44628
rect 34660 -44772 34724 -44708
rect 34660 -44852 34724 -44788
rect 34660 -44932 34724 -44868
rect 34660 -45012 34724 -44948
rect 34660 -45092 34724 -45028
rect 34660 -45172 34724 -45108
rect 34660 -45252 34724 -45188
rect 34660 -45332 34724 -45268
rect 34660 -45412 34724 -45348
rect 34660 -45492 34724 -45428
rect 34660 -45572 34724 -45508
rect 34660 -45652 34724 -45588
rect 34660 -45732 34724 -45668
rect 34660 -45812 34724 -45748
rect 34660 -45892 34724 -45828
rect 34660 -45972 34724 -45908
rect 34660 -46052 34724 -45988
rect 34660 -46132 34724 -46068
rect 34660 -46212 34724 -46148
rect 34660 -46292 34724 -46228
rect 34660 -46372 34724 -46308
rect 34660 -46452 34724 -46388
rect 34660 -46532 34724 -46468
rect 34660 -46612 34724 -46548
rect 34660 -46692 34724 -46628
rect 34660 -46772 34724 -46708
rect 34660 -46852 34724 -46788
rect 34660 -46932 34724 -46868
rect 34660 -47012 34724 -46948
rect 34660 -47092 34724 -47028
rect 34660 -47172 34724 -47108
rect 40979 -41092 41043 -41028
rect 40979 -41172 41043 -41108
rect 40979 -41252 41043 -41188
rect 40979 -41332 41043 -41268
rect 40979 -41412 41043 -41348
rect 40979 -41492 41043 -41428
rect 40979 -41572 41043 -41508
rect 40979 -41652 41043 -41588
rect 40979 -41732 41043 -41668
rect 40979 -41812 41043 -41748
rect 40979 -41892 41043 -41828
rect 40979 -41972 41043 -41908
rect 40979 -42052 41043 -41988
rect 40979 -42132 41043 -42068
rect 40979 -42212 41043 -42148
rect 40979 -42292 41043 -42228
rect 40979 -42372 41043 -42308
rect 40979 -42452 41043 -42388
rect 40979 -42532 41043 -42468
rect 40979 -42612 41043 -42548
rect 40979 -42692 41043 -42628
rect 40979 -42772 41043 -42708
rect 40979 -42852 41043 -42788
rect 40979 -42932 41043 -42868
rect 40979 -43012 41043 -42948
rect 40979 -43092 41043 -43028
rect 40979 -43172 41043 -43108
rect 40979 -43252 41043 -43188
rect 40979 -43332 41043 -43268
rect 40979 -43412 41043 -43348
rect 40979 -43492 41043 -43428
rect 40979 -43572 41043 -43508
rect 40979 -43652 41043 -43588
rect 40979 -43732 41043 -43668
rect 40979 -43812 41043 -43748
rect 40979 -43892 41043 -43828
rect 40979 -43972 41043 -43908
rect 40979 -44052 41043 -43988
rect 40979 -44132 41043 -44068
rect 40979 -44212 41043 -44148
rect 40979 -44292 41043 -44228
rect 40979 -44372 41043 -44308
rect 40979 -44452 41043 -44388
rect 40979 -44532 41043 -44468
rect 40979 -44612 41043 -44548
rect 40979 -44692 41043 -44628
rect 40979 -44772 41043 -44708
rect 40979 -44852 41043 -44788
rect 40979 -44932 41043 -44868
rect 40979 -45012 41043 -44948
rect 40979 -45092 41043 -45028
rect 40979 -45172 41043 -45108
rect 40979 -45252 41043 -45188
rect 40979 -45332 41043 -45268
rect 40979 -45412 41043 -45348
rect 40979 -45492 41043 -45428
rect 40979 -45572 41043 -45508
rect 40979 -45652 41043 -45588
rect 40979 -45732 41043 -45668
rect 40979 -45812 41043 -45748
rect 40979 -45892 41043 -45828
rect 40979 -45972 41043 -45908
rect 40979 -46052 41043 -45988
rect 40979 -46132 41043 -46068
rect 40979 -46212 41043 -46148
rect 40979 -46292 41043 -46228
rect 40979 -46372 41043 -46308
rect 40979 -46452 41043 -46388
rect 40979 -46532 41043 -46468
rect 40979 -46612 41043 -46548
rect 40979 -46692 41043 -46628
rect 40979 -46772 41043 -46708
rect 40979 -46852 41043 -46788
rect 40979 -46932 41043 -46868
rect 40979 -47012 41043 -46948
rect 40979 -47092 41043 -47028
rect 40979 -47172 41043 -47108
rect 47298 -41092 47362 -41028
rect 47298 -41172 47362 -41108
rect 47298 -41252 47362 -41188
rect 47298 -41332 47362 -41268
rect 47298 -41412 47362 -41348
rect 47298 -41492 47362 -41428
rect 47298 -41572 47362 -41508
rect 47298 -41652 47362 -41588
rect 47298 -41732 47362 -41668
rect 47298 -41812 47362 -41748
rect 47298 -41892 47362 -41828
rect 47298 -41972 47362 -41908
rect 47298 -42052 47362 -41988
rect 47298 -42132 47362 -42068
rect 47298 -42212 47362 -42148
rect 47298 -42292 47362 -42228
rect 47298 -42372 47362 -42308
rect 47298 -42452 47362 -42388
rect 47298 -42532 47362 -42468
rect 47298 -42612 47362 -42548
rect 47298 -42692 47362 -42628
rect 47298 -42772 47362 -42708
rect 47298 -42852 47362 -42788
rect 47298 -42932 47362 -42868
rect 47298 -43012 47362 -42948
rect 47298 -43092 47362 -43028
rect 47298 -43172 47362 -43108
rect 47298 -43252 47362 -43188
rect 47298 -43332 47362 -43268
rect 47298 -43412 47362 -43348
rect 47298 -43492 47362 -43428
rect 47298 -43572 47362 -43508
rect 47298 -43652 47362 -43588
rect 47298 -43732 47362 -43668
rect 47298 -43812 47362 -43748
rect 47298 -43892 47362 -43828
rect 47298 -43972 47362 -43908
rect 47298 -44052 47362 -43988
rect 47298 -44132 47362 -44068
rect 47298 -44212 47362 -44148
rect 47298 -44292 47362 -44228
rect 47298 -44372 47362 -44308
rect 47298 -44452 47362 -44388
rect 47298 -44532 47362 -44468
rect 47298 -44612 47362 -44548
rect 47298 -44692 47362 -44628
rect 47298 -44772 47362 -44708
rect 47298 -44852 47362 -44788
rect 47298 -44932 47362 -44868
rect 47298 -45012 47362 -44948
rect 47298 -45092 47362 -45028
rect 47298 -45172 47362 -45108
rect 47298 -45252 47362 -45188
rect 47298 -45332 47362 -45268
rect 47298 -45412 47362 -45348
rect 47298 -45492 47362 -45428
rect 47298 -45572 47362 -45508
rect 47298 -45652 47362 -45588
rect 47298 -45732 47362 -45668
rect 47298 -45812 47362 -45748
rect 47298 -45892 47362 -45828
rect 47298 -45972 47362 -45908
rect 47298 -46052 47362 -45988
rect 47298 -46132 47362 -46068
rect 47298 -46212 47362 -46148
rect 47298 -46292 47362 -46228
rect 47298 -46372 47362 -46308
rect 47298 -46452 47362 -46388
rect 47298 -46532 47362 -46468
rect 47298 -46612 47362 -46548
rect 47298 -46692 47362 -46628
rect 47298 -46772 47362 -46708
rect 47298 -46852 47362 -46788
rect 47298 -46932 47362 -46868
rect 47298 -47012 47362 -46948
rect 47298 -47092 47362 -47028
rect 47298 -47172 47362 -47108
<< mimcap >>
rect -47283 47052 -41283 47100
rect -47283 41148 -47235 47052
rect -41331 41148 -41283 47052
rect -47283 41100 -41283 41148
rect -40964 47052 -34964 47100
rect -40964 41148 -40916 47052
rect -35012 41148 -34964 47052
rect -40964 41100 -34964 41148
rect -34645 47052 -28645 47100
rect -34645 41148 -34597 47052
rect -28693 41148 -28645 47052
rect -34645 41100 -28645 41148
rect -28326 47052 -22326 47100
rect -28326 41148 -28278 47052
rect -22374 41148 -22326 47052
rect -28326 41100 -22326 41148
rect -22007 47052 -16007 47100
rect -22007 41148 -21959 47052
rect -16055 41148 -16007 47052
rect -22007 41100 -16007 41148
rect -15688 47052 -9688 47100
rect -15688 41148 -15640 47052
rect -9736 41148 -9688 47052
rect -15688 41100 -9688 41148
rect -9369 47052 -3369 47100
rect -9369 41148 -9321 47052
rect -3417 41148 -3369 47052
rect -9369 41100 -3369 41148
rect -3050 47052 2950 47100
rect -3050 41148 -3002 47052
rect 2902 41148 2950 47052
rect -3050 41100 2950 41148
rect 3269 47052 9269 47100
rect 3269 41148 3317 47052
rect 9221 41148 9269 47052
rect 3269 41100 9269 41148
rect 9588 47052 15588 47100
rect 9588 41148 9636 47052
rect 15540 41148 15588 47052
rect 9588 41100 15588 41148
rect 15907 47052 21907 47100
rect 15907 41148 15955 47052
rect 21859 41148 21907 47052
rect 15907 41100 21907 41148
rect 22226 47052 28226 47100
rect 22226 41148 22274 47052
rect 28178 41148 28226 47052
rect 22226 41100 28226 41148
rect 28545 47052 34545 47100
rect 28545 41148 28593 47052
rect 34497 41148 34545 47052
rect 28545 41100 34545 41148
rect 34864 47052 40864 47100
rect 34864 41148 34912 47052
rect 40816 41148 40864 47052
rect 34864 41100 40864 41148
rect 41183 47052 47183 47100
rect 41183 41148 41231 47052
rect 47135 41148 47183 47052
rect 41183 41100 47183 41148
rect -47283 40752 -41283 40800
rect -47283 34848 -47235 40752
rect -41331 34848 -41283 40752
rect -47283 34800 -41283 34848
rect -40964 40752 -34964 40800
rect -40964 34848 -40916 40752
rect -35012 34848 -34964 40752
rect -40964 34800 -34964 34848
rect -34645 40752 -28645 40800
rect -34645 34848 -34597 40752
rect -28693 34848 -28645 40752
rect -34645 34800 -28645 34848
rect -28326 40752 -22326 40800
rect -28326 34848 -28278 40752
rect -22374 34848 -22326 40752
rect -28326 34800 -22326 34848
rect -22007 40752 -16007 40800
rect -22007 34848 -21959 40752
rect -16055 34848 -16007 40752
rect -22007 34800 -16007 34848
rect -15688 40752 -9688 40800
rect -15688 34848 -15640 40752
rect -9736 34848 -9688 40752
rect -15688 34800 -9688 34848
rect -9369 40752 -3369 40800
rect -9369 34848 -9321 40752
rect -3417 34848 -3369 40752
rect -9369 34800 -3369 34848
rect -3050 40752 2950 40800
rect -3050 34848 -3002 40752
rect 2902 34848 2950 40752
rect -3050 34800 2950 34848
rect 3269 40752 9269 40800
rect 3269 34848 3317 40752
rect 9221 34848 9269 40752
rect 3269 34800 9269 34848
rect 9588 40752 15588 40800
rect 9588 34848 9636 40752
rect 15540 34848 15588 40752
rect 9588 34800 15588 34848
rect 15907 40752 21907 40800
rect 15907 34848 15955 40752
rect 21859 34848 21907 40752
rect 15907 34800 21907 34848
rect 22226 40752 28226 40800
rect 22226 34848 22274 40752
rect 28178 34848 28226 40752
rect 22226 34800 28226 34848
rect 28545 40752 34545 40800
rect 28545 34848 28593 40752
rect 34497 34848 34545 40752
rect 28545 34800 34545 34848
rect 34864 40752 40864 40800
rect 34864 34848 34912 40752
rect 40816 34848 40864 40752
rect 34864 34800 40864 34848
rect 41183 40752 47183 40800
rect 41183 34848 41231 40752
rect 47135 34848 47183 40752
rect 41183 34800 47183 34848
rect -47283 34452 -41283 34500
rect -47283 28548 -47235 34452
rect -41331 28548 -41283 34452
rect -47283 28500 -41283 28548
rect -40964 34452 -34964 34500
rect -40964 28548 -40916 34452
rect -35012 28548 -34964 34452
rect -40964 28500 -34964 28548
rect -34645 34452 -28645 34500
rect -34645 28548 -34597 34452
rect -28693 28548 -28645 34452
rect -34645 28500 -28645 28548
rect -28326 34452 -22326 34500
rect -28326 28548 -28278 34452
rect -22374 28548 -22326 34452
rect -28326 28500 -22326 28548
rect -22007 34452 -16007 34500
rect -22007 28548 -21959 34452
rect -16055 28548 -16007 34452
rect -22007 28500 -16007 28548
rect -15688 34452 -9688 34500
rect -15688 28548 -15640 34452
rect -9736 28548 -9688 34452
rect -15688 28500 -9688 28548
rect -9369 34452 -3369 34500
rect -9369 28548 -9321 34452
rect -3417 28548 -3369 34452
rect -9369 28500 -3369 28548
rect -3050 34452 2950 34500
rect -3050 28548 -3002 34452
rect 2902 28548 2950 34452
rect -3050 28500 2950 28548
rect 3269 34452 9269 34500
rect 3269 28548 3317 34452
rect 9221 28548 9269 34452
rect 3269 28500 9269 28548
rect 9588 34452 15588 34500
rect 9588 28548 9636 34452
rect 15540 28548 15588 34452
rect 9588 28500 15588 28548
rect 15907 34452 21907 34500
rect 15907 28548 15955 34452
rect 21859 28548 21907 34452
rect 15907 28500 21907 28548
rect 22226 34452 28226 34500
rect 22226 28548 22274 34452
rect 28178 28548 28226 34452
rect 22226 28500 28226 28548
rect 28545 34452 34545 34500
rect 28545 28548 28593 34452
rect 34497 28548 34545 34452
rect 28545 28500 34545 28548
rect 34864 34452 40864 34500
rect 34864 28548 34912 34452
rect 40816 28548 40864 34452
rect 34864 28500 40864 28548
rect 41183 34452 47183 34500
rect 41183 28548 41231 34452
rect 47135 28548 47183 34452
rect 41183 28500 47183 28548
rect -47283 28152 -41283 28200
rect -47283 22248 -47235 28152
rect -41331 22248 -41283 28152
rect -47283 22200 -41283 22248
rect -40964 28152 -34964 28200
rect -40964 22248 -40916 28152
rect -35012 22248 -34964 28152
rect -40964 22200 -34964 22248
rect -34645 28152 -28645 28200
rect -34645 22248 -34597 28152
rect -28693 22248 -28645 28152
rect -34645 22200 -28645 22248
rect -28326 28152 -22326 28200
rect -28326 22248 -28278 28152
rect -22374 22248 -22326 28152
rect -28326 22200 -22326 22248
rect -22007 28152 -16007 28200
rect -22007 22248 -21959 28152
rect -16055 22248 -16007 28152
rect -22007 22200 -16007 22248
rect -15688 28152 -9688 28200
rect -15688 22248 -15640 28152
rect -9736 22248 -9688 28152
rect -15688 22200 -9688 22248
rect -9369 28152 -3369 28200
rect -9369 22248 -9321 28152
rect -3417 22248 -3369 28152
rect -9369 22200 -3369 22248
rect -3050 28152 2950 28200
rect -3050 22248 -3002 28152
rect 2902 22248 2950 28152
rect -3050 22200 2950 22248
rect 3269 28152 9269 28200
rect 3269 22248 3317 28152
rect 9221 22248 9269 28152
rect 3269 22200 9269 22248
rect 9588 28152 15588 28200
rect 9588 22248 9636 28152
rect 15540 22248 15588 28152
rect 9588 22200 15588 22248
rect 15907 28152 21907 28200
rect 15907 22248 15955 28152
rect 21859 22248 21907 28152
rect 15907 22200 21907 22248
rect 22226 28152 28226 28200
rect 22226 22248 22274 28152
rect 28178 22248 28226 28152
rect 22226 22200 28226 22248
rect 28545 28152 34545 28200
rect 28545 22248 28593 28152
rect 34497 22248 34545 28152
rect 28545 22200 34545 22248
rect 34864 28152 40864 28200
rect 34864 22248 34912 28152
rect 40816 22248 40864 28152
rect 34864 22200 40864 22248
rect 41183 28152 47183 28200
rect 41183 22248 41231 28152
rect 47135 22248 47183 28152
rect 41183 22200 47183 22248
rect -47283 21852 -41283 21900
rect -47283 15948 -47235 21852
rect -41331 15948 -41283 21852
rect -47283 15900 -41283 15948
rect -40964 21852 -34964 21900
rect -40964 15948 -40916 21852
rect -35012 15948 -34964 21852
rect -40964 15900 -34964 15948
rect -34645 21852 -28645 21900
rect -34645 15948 -34597 21852
rect -28693 15948 -28645 21852
rect -34645 15900 -28645 15948
rect -28326 21852 -22326 21900
rect -28326 15948 -28278 21852
rect -22374 15948 -22326 21852
rect -28326 15900 -22326 15948
rect -22007 21852 -16007 21900
rect -22007 15948 -21959 21852
rect -16055 15948 -16007 21852
rect -22007 15900 -16007 15948
rect -15688 21852 -9688 21900
rect -15688 15948 -15640 21852
rect -9736 15948 -9688 21852
rect -15688 15900 -9688 15948
rect -9369 21852 -3369 21900
rect -9369 15948 -9321 21852
rect -3417 15948 -3369 21852
rect -9369 15900 -3369 15948
rect -3050 21852 2950 21900
rect -3050 15948 -3002 21852
rect 2902 15948 2950 21852
rect -3050 15900 2950 15948
rect 3269 21852 9269 21900
rect 3269 15948 3317 21852
rect 9221 15948 9269 21852
rect 3269 15900 9269 15948
rect 9588 21852 15588 21900
rect 9588 15948 9636 21852
rect 15540 15948 15588 21852
rect 9588 15900 15588 15948
rect 15907 21852 21907 21900
rect 15907 15948 15955 21852
rect 21859 15948 21907 21852
rect 15907 15900 21907 15948
rect 22226 21852 28226 21900
rect 22226 15948 22274 21852
rect 28178 15948 28226 21852
rect 22226 15900 28226 15948
rect 28545 21852 34545 21900
rect 28545 15948 28593 21852
rect 34497 15948 34545 21852
rect 28545 15900 34545 15948
rect 34864 21852 40864 21900
rect 34864 15948 34912 21852
rect 40816 15948 40864 21852
rect 34864 15900 40864 15948
rect 41183 21852 47183 21900
rect 41183 15948 41231 21852
rect 47135 15948 47183 21852
rect 41183 15900 47183 15948
rect -47283 15552 -41283 15600
rect -47283 9648 -47235 15552
rect -41331 9648 -41283 15552
rect -47283 9600 -41283 9648
rect -40964 15552 -34964 15600
rect -40964 9648 -40916 15552
rect -35012 9648 -34964 15552
rect -40964 9600 -34964 9648
rect -34645 15552 -28645 15600
rect -34645 9648 -34597 15552
rect -28693 9648 -28645 15552
rect -34645 9600 -28645 9648
rect -28326 15552 -22326 15600
rect -28326 9648 -28278 15552
rect -22374 9648 -22326 15552
rect -28326 9600 -22326 9648
rect -22007 15552 -16007 15600
rect -22007 9648 -21959 15552
rect -16055 9648 -16007 15552
rect -22007 9600 -16007 9648
rect -15688 15552 -9688 15600
rect -15688 9648 -15640 15552
rect -9736 9648 -9688 15552
rect -15688 9600 -9688 9648
rect -9369 15552 -3369 15600
rect -9369 9648 -9321 15552
rect -3417 9648 -3369 15552
rect -9369 9600 -3369 9648
rect -3050 15552 2950 15600
rect -3050 9648 -3002 15552
rect 2902 9648 2950 15552
rect -3050 9600 2950 9648
rect 3269 15552 9269 15600
rect 3269 9648 3317 15552
rect 9221 9648 9269 15552
rect 3269 9600 9269 9648
rect 9588 15552 15588 15600
rect 9588 9648 9636 15552
rect 15540 9648 15588 15552
rect 9588 9600 15588 9648
rect 15907 15552 21907 15600
rect 15907 9648 15955 15552
rect 21859 9648 21907 15552
rect 15907 9600 21907 9648
rect 22226 15552 28226 15600
rect 22226 9648 22274 15552
rect 28178 9648 28226 15552
rect 22226 9600 28226 9648
rect 28545 15552 34545 15600
rect 28545 9648 28593 15552
rect 34497 9648 34545 15552
rect 28545 9600 34545 9648
rect 34864 15552 40864 15600
rect 34864 9648 34912 15552
rect 40816 9648 40864 15552
rect 34864 9600 40864 9648
rect 41183 15552 47183 15600
rect 41183 9648 41231 15552
rect 47135 9648 47183 15552
rect 41183 9600 47183 9648
rect -47283 9252 -41283 9300
rect -47283 3348 -47235 9252
rect -41331 3348 -41283 9252
rect -47283 3300 -41283 3348
rect -40964 9252 -34964 9300
rect -40964 3348 -40916 9252
rect -35012 3348 -34964 9252
rect -40964 3300 -34964 3348
rect -34645 9252 -28645 9300
rect -34645 3348 -34597 9252
rect -28693 3348 -28645 9252
rect -34645 3300 -28645 3348
rect -28326 9252 -22326 9300
rect -28326 3348 -28278 9252
rect -22374 3348 -22326 9252
rect -28326 3300 -22326 3348
rect -22007 9252 -16007 9300
rect -22007 3348 -21959 9252
rect -16055 3348 -16007 9252
rect -22007 3300 -16007 3348
rect -15688 9252 -9688 9300
rect -15688 3348 -15640 9252
rect -9736 3348 -9688 9252
rect -15688 3300 -9688 3348
rect -9369 9252 -3369 9300
rect -9369 3348 -9321 9252
rect -3417 3348 -3369 9252
rect -9369 3300 -3369 3348
rect -3050 9252 2950 9300
rect -3050 3348 -3002 9252
rect 2902 3348 2950 9252
rect -3050 3300 2950 3348
rect 3269 9252 9269 9300
rect 3269 3348 3317 9252
rect 9221 3348 9269 9252
rect 3269 3300 9269 3348
rect 9588 9252 15588 9300
rect 9588 3348 9636 9252
rect 15540 3348 15588 9252
rect 9588 3300 15588 3348
rect 15907 9252 21907 9300
rect 15907 3348 15955 9252
rect 21859 3348 21907 9252
rect 15907 3300 21907 3348
rect 22226 9252 28226 9300
rect 22226 3348 22274 9252
rect 28178 3348 28226 9252
rect 22226 3300 28226 3348
rect 28545 9252 34545 9300
rect 28545 3348 28593 9252
rect 34497 3348 34545 9252
rect 28545 3300 34545 3348
rect 34864 9252 40864 9300
rect 34864 3348 34912 9252
rect 40816 3348 40864 9252
rect 34864 3300 40864 3348
rect 41183 9252 47183 9300
rect 41183 3348 41231 9252
rect 47135 3348 47183 9252
rect 41183 3300 47183 3348
rect -47283 2952 -41283 3000
rect -47283 -2952 -47235 2952
rect -41331 -2952 -41283 2952
rect -47283 -3000 -41283 -2952
rect -40964 2952 -34964 3000
rect -40964 -2952 -40916 2952
rect -35012 -2952 -34964 2952
rect -40964 -3000 -34964 -2952
rect -34645 2952 -28645 3000
rect -34645 -2952 -34597 2952
rect -28693 -2952 -28645 2952
rect -34645 -3000 -28645 -2952
rect -28326 2952 -22326 3000
rect -28326 -2952 -28278 2952
rect -22374 -2952 -22326 2952
rect -28326 -3000 -22326 -2952
rect -22007 2952 -16007 3000
rect -22007 -2952 -21959 2952
rect -16055 -2952 -16007 2952
rect -22007 -3000 -16007 -2952
rect -15688 2952 -9688 3000
rect -15688 -2952 -15640 2952
rect -9736 -2952 -9688 2952
rect -15688 -3000 -9688 -2952
rect -9369 2952 -3369 3000
rect -9369 -2952 -9321 2952
rect -3417 -2952 -3369 2952
rect -9369 -3000 -3369 -2952
rect -3050 2952 2950 3000
rect -3050 -2952 -3002 2952
rect 2902 -2952 2950 2952
rect -3050 -3000 2950 -2952
rect 3269 2952 9269 3000
rect 3269 -2952 3317 2952
rect 9221 -2952 9269 2952
rect 3269 -3000 9269 -2952
rect 9588 2952 15588 3000
rect 9588 -2952 9636 2952
rect 15540 -2952 15588 2952
rect 9588 -3000 15588 -2952
rect 15907 2952 21907 3000
rect 15907 -2952 15955 2952
rect 21859 -2952 21907 2952
rect 15907 -3000 21907 -2952
rect 22226 2952 28226 3000
rect 22226 -2952 22274 2952
rect 28178 -2952 28226 2952
rect 22226 -3000 28226 -2952
rect 28545 2952 34545 3000
rect 28545 -2952 28593 2952
rect 34497 -2952 34545 2952
rect 28545 -3000 34545 -2952
rect 34864 2952 40864 3000
rect 34864 -2952 34912 2952
rect 40816 -2952 40864 2952
rect 34864 -3000 40864 -2952
rect 41183 2952 47183 3000
rect 41183 -2952 41231 2952
rect 47135 -2952 47183 2952
rect 41183 -3000 47183 -2952
rect -47283 -3348 -41283 -3300
rect -47283 -9252 -47235 -3348
rect -41331 -9252 -41283 -3348
rect -47283 -9300 -41283 -9252
rect -40964 -3348 -34964 -3300
rect -40964 -9252 -40916 -3348
rect -35012 -9252 -34964 -3348
rect -40964 -9300 -34964 -9252
rect -34645 -3348 -28645 -3300
rect -34645 -9252 -34597 -3348
rect -28693 -9252 -28645 -3348
rect -34645 -9300 -28645 -9252
rect -28326 -3348 -22326 -3300
rect -28326 -9252 -28278 -3348
rect -22374 -9252 -22326 -3348
rect -28326 -9300 -22326 -9252
rect -22007 -3348 -16007 -3300
rect -22007 -9252 -21959 -3348
rect -16055 -9252 -16007 -3348
rect -22007 -9300 -16007 -9252
rect -15688 -3348 -9688 -3300
rect -15688 -9252 -15640 -3348
rect -9736 -9252 -9688 -3348
rect -15688 -9300 -9688 -9252
rect -9369 -3348 -3369 -3300
rect -9369 -9252 -9321 -3348
rect -3417 -9252 -3369 -3348
rect -9369 -9300 -3369 -9252
rect -3050 -3348 2950 -3300
rect -3050 -9252 -3002 -3348
rect 2902 -9252 2950 -3348
rect -3050 -9300 2950 -9252
rect 3269 -3348 9269 -3300
rect 3269 -9252 3317 -3348
rect 9221 -9252 9269 -3348
rect 3269 -9300 9269 -9252
rect 9588 -3348 15588 -3300
rect 9588 -9252 9636 -3348
rect 15540 -9252 15588 -3348
rect 9588 -9300 15588 -9252
rect 15907 -3348 21907 -3300
rect 15907 -9252 15955 -3348
rect 21859 -9252 21907 -3348
rect 15907 -9300 21907 -9252
rect 22226 -3348 28226 -3300
rect 22226 -9252 22274 -3348
rect 28178 -9252 28226 -3348
rect 22226 -9300 28226 -9252
rect 28545 -3348 34545 -3300
rect 28545 -9252 28593 -3348
rect 34497 -9252 34545 -3348
rect 28545 -9300 34545 -9252
rect 34864 -3348 40864 -3300
rect 34864 -9252 34912 -3348
rect 40816 -9252 40864 -3348
rect 34864 -9300 40864 -9252
rect 41183 -3348 47183 -3300
rect 41183 -9252 41231 -3348
rect 47135 -9252 47183 -3348
rect 41183 -9300 47183 -9252
rect -47283 -9648 -41283 -9600
rect -47283 -15552 -47235 -9648
rect -41331 -15552 -41283 -9648
rect -47283 -15600 -41283 -15552
rect -40964 -9648 -34964 -9600
rect -40964 -15552 -40916 -9648
rect -35012 -15552 -34964 -9648
rect -40964 -15600 -34964 -15552
rect -34645 -9648 -28645 -9600
rect -34645 -15552 -34597 -9648
rect -28693 -15552 -28645 -9648
rect -34645 -15600 -28645 -15552
rect -28326 -9648 -22326 -9600
rect -28326 -15552 -28278 -9648
rect -22374 -15552 -22326 -9648
rect -28326 -15600 -22326 -15552
rect -22007 -9648 -16007 -9600
rect -22007 -15552 -21959 -9648
rect -16055 -15552 -16007 -9648
rect -22007 -15600 -16007 -15552
rect -15688 -9648 -9688 -9600
rect -15688 -15552 -15640 -9648
rect -9736 -15552 -9688 -9648
rect -15688 -15600 -9688 -15552
rect -9369 -9648 -3369 -9600
rect -9369 -15552 -9321 -9648
rect -3417 -15552 -3369 -9648
rect -9369 -15600 -3369 -15552
rect -3050 -9648 2950 -9600
rect -3050 -15552 -3002 -9648
rect 2902 -15552 2950 -9648
rect -3050 -15600 2950 -15552
rect 3269 -9648 9269 -9600
rect 3269 -15552 3317 -9648
rect 9221 -15552 9269 -9648
rect 3269 -15600 9269 -15552
rect 9588 -9648 15588 -9600
rect 9588 -15552 9636 -9648
rect 15540 -15552 15588 -9648
rect 9588 -15600 15588 -15552
rect 15907 -9648 21907 -9600
rect 15907 -15552 15955 -9648
rect 21859 -15552 21907 -9648
rect 15907 -15600 21907 -15552
rect 22226 -9648 28226 -9600
rect 22226 -15552 22274 -9648
rect 28178 -15552 28226 -9648
rect 22226 -15600 28226 -15552
rect 28545 -9648 34545 -9600
rect 28545 -15552 28593 -9648
rect 34497 -15552 34545 -9648
rect 28545 -15600 34545 -15552
rect 34864 -9648 40864 -9600
rect 34864 -15552 34912 -9648
rect 40816 -15552 40864 -9648
rect 34864 -15600 40864 -15552
rect 41183 -9648 47183 -9600
rect 41183 -15552 41231 -9648
rect 47135 -15552 47183 -9648
rect 41183 -15600 47183 -15552
rect -47283 -15948 -41283 -15900
rect -47283 -21852 -47235 -15948
rect -41331 -21852 -41283 -15948
rect -47283 -21900 -41283 -21852
rect -40964 -15948 -34964 -15900
rect -40964 -21852 -40916 -15948
rect -35012 -21852 -34964 -15948
rect -40964 -21900 -34964 -21852
rect -34645 -15948 -28645 -15900
rect -34645 -21852 -34597 -15948
rect -28693 -21852 -28645 -15948
rect -34645 -21900 -28645 -21852
rect -28326 -15948 -22326 -15900
rect -28326 -21852 -28278 -15948
rect -22374 -21852 -22326 -15948
rect -28326 -21900 -22326 -21852
rect -22007 -15948 -16007 -15900
rect -22007 -21852 -21959 -15948
rect -16055 -21852 -16007 -15948
rect -22007 -21900 -16007 -21852
rect -15688 -15948 -9688 -15900
rect -15688 -21852 -15640 -15948
rect -9736 -21852 -9688 -15948
rect -15688 -21900 -9688 -21852
rect -9369 -15948 -3369 -15900
rect -9369 -21852 -9321 -15948
rect -3417 -21852 -3369 -15948
rect -9369 -21900 -3369 -21852
rect -3050 -15948 2950 -15900
rect -3050 -21852 -3002 -15948
rect 2902 -21852 2950 -15948
rect -3050 -21900 2950 -21852
rect 3269 -15948 9269 -15900
rect 3269 -21852 3317 -15948
rect 9221 -21852 9269 -15948
rect 3269 -21900 9269 -21852
rect 9588 -15948 15588 -15900
rect 9588 -21852 9636 -15948
rect 15540 -21852 15588 -15948
rect 9588 -21900 15588 -21852
rect 15907 -15948 21907 -15900
rect 15907 -21852 15955 -15948
rect 21859 -21852 21907 -15948
rect 15907 -21900 21907 -21852
rect 22226 -15948 28226 -15900
rect 22226 -21852 22274 -15948
rect 28178 -21852 28226 -15948
rect 22226 -21900 28226 -21852
rect 28545 -15948 34545 -15900
rect 28545 -21852 28593 -15948
rect 34497 -21852 34545 -15948
rect 28545 -21900 34545 -21852
rect 34864 -15948 40864 -15900
rect 34864 -21852 34912 -15948
rect 40816 -21852 40864 -15948
rect 34864 -21900 40864 -21852
rect 41183 -15948 47183 -15900
rect 41183 -21852 41231 -15948
rect 47135 -21852 47183 -15948
rect 41183 -21900 47183 -21852
rect -47283 -22248 -41283 -22200
rect -47283 -28152 -47235 -22248
rect -41331 -28152 -41283 -22248
rect -47283 -28200 -41283 -28152
rect -40964 -22248 -34964 -22200
rect -40964 -28152 -40916 -22248
rect -35012 -28152 -34964 -22248
rect -40964 -28200 -34964 -28152
rect -34645 -22248 -28645 -22200
rect -34645 -28152 -34597 -22248
rect -28693 -28152 -28645 -22248
rect -34645 -28200 -28645 -28152
rect -28326 -22248 -22326 -22200
rect -28326 -28152 -28278 -22248
rect -22374 -28152 -22326 -22248
rect -28326 -28200 -22326 -28152
rect -22007 -22248 -16007 -22200
rect -22007 -28152 -21959 -22248
rect -16055 -28152 -16007 -22248
rect -22007 -28200 -16007 -28152
rect -15688 -22248 -9688 -22200
rect -15688 -28152 -15640 -22248
rect -9736 -28152 -9688 -22248
rect -15688 -28200 -9688 -28152
rect -9369 -22248 -3369 -22200
rect -9369 -28152 -9321 -22248
rect -3417 -28152 -3369 -22248
rect -9369 -28200 -3369 -28152
rect -3050 -22248 2950 -22200
rect -3050 -28152 -3002 -22248
rect 2902 -28152 2950 -22248
rect -3050 -28200 2950 -28152
rect 3269 -22248 9269 -22200
rect 3269 -28152 3317 -22248
rect 9221 -28152 9269 -22248
rect 3269 -28200 9269 -28152
rect 9588 -22248 15588 -22200
rect 9588 -28152 9636 -22248
rect 15540 -28152 15588 -22248
rect 9588 -28200 15588 -28152
rect 15907 -22248 21907 -22200
rect 15907 -28152 15955 -22248
rect 21859 -28152 21907 -22248
rect 15907 -28200 21907 -28152
rect 22226 -22248 28226 -22200
rect 22226 -28152 22274 -22248
rect 28178 -28152 28226 -22248
rect 22226 -28200 28226 -28152
rect 28545 -22248 34545 -22200
rect 28545 -28152 28593 -22248
rect 34497 -28152 34545 -22248
rect 28545 -28200 34545 -28152
rect 34864 -22248 40864 -22200
rect 34864 -28152 34912 -22248
rect 40816 -28152 40864 -22248
rect 34864 -28200 40864 -28152
rect 41183 -22248 47183 -22200
rect 41183 -28152 41231 -22248
rect 47135 -28152 47183 -22248
rect 41183 -28200 47183 -28152
rect -47283 -28548 -41283 -28500
rect -47283 -34452 -47235 -28548
rect -41331 -34452 -41283 -28548
rect -47283 -34500 -41283 -34452
rect -40964 -28548 -34964 -28500
rect -40964 -34452 -40916 -28548
rect -35012 -34452 -34964 -28548
rect -40964 -34500 -34964 -34452
rect -34645 -28548 -28645 -28500
rect -34645 -34452 -34597 -28548
rect -28693 -34452 -28645 -28548
rect -34645 -34500 -28645 -34452
rect -28326 -28548 -22326 -28500
rect -28326 -34452 -28278 -28548
rect -22374 -34452 -22326 -28548
rect -28326 -34500 -22326 -34452
rect -22007 -28548 -16007 -28500
rect -22007 -34452 -21959 -28548
rect -16055 -34452 -16007 -28548
rect -22007 -34500 -16007 -34452
rect -15688 -28548 -9688 -28500
rect -15688 -34452 -15640 -28548
rect -9736 -34452 -9688 -28548
rect -15688 -34500 -9688 -34452
rect -9369 -28548 -3369 -28500
rect -9369 -34452 -9321 -28548
rect -3417 -34452 -3369 -28548
rect -9369 -34500 -3369 -34452
rect -3050 -28548 2950 -28500
rect -3050 -34452 -3002 -28548
rect 2902 -34452 2950 -28548
rect -3050 -34500 2950 -34452
rect 3269 -28548 9269 -28500
rect 3269 -34452 3317 -28548
rect 9221 -34452 9269 -28548
rect 3269 -34500 9269 -34452
rect 9588 -28548 15588 -28500
rect 9588 -34452 9636 -28548
rect 15540 -34452 15588 -28548
rect 9588 -34500 15588 -34452
rect 15907 -28548 21907 -28500
rect 15907 -34452 15955 -28548
rect 21859 -34452 21907 -28548
rect 15907 -34500 21907 -34452
rect 22226 -28548 28226 -28500
rect 22226 -34452 22274 -28548
rect 28178 -34452 28226 -28548
rect 22226 -34500 28226 -34452
rect 28545 -28548 34545 -28500
rect 28545 -34452 28593 -28548
rect 34497 -34452 34545 -28548
rect 28545 -34500 34545 -34452
rect 34864 -28548 40864 -28500
rect 34864 -34452 34912 -28548
rect 40816 -34452 40864 -28548
rect 34864 -34500 40864 -34452
rect 41183 -28548 47183 -28500
rect 41183 -34452 41231 -28548
rect 47135 -34452 47183 -28548
rect 41183 -34500 47183 -34452
rect -47283 -34848 -41283 -34800
rect -47283 -40752 -47235 -34848
rect -41331 -40752 -41283 -34848
rect -47283 -40800 -41283 -40752
rect -40964 -34848 -34964 -34800
rect -40964 -40752 -40916 -34848
rect -35012 -40752 -34964 -34848
rect -40964 -40800 -34964 -40752
rect -34645 -34848 -28645 -34800
rect -34645 -40752 -34597 -34848
rect -28693 -40752 -28645 -34848
rect -34645 -40800 -28645 -40752
rect -28326 -34848 -22326 -34800
rect -28326 -40752 -28278 -34848
rect -22374 -40752 -22326 -34848
rect -28326 -40800 -22326 -40752
rect -22007 -34848 -16007 -34800
rect -22007 -40752 -21959 -34848
rect -16055 -40752 -16007 -34848
rect -22007 -40800 -16007 -40752
rect -15688 -34848 -9688 -34800
rect -15688 -40752 -15640 -34848
rect -9736 -40752 -9688 -34848
rect -15688 -40800 -9688 -40752
rect -9369 -34848 -3369 -34800
rect -9369 -40752 -9321 -34848
rect -3417 -40752 -3369 -34848
rect -9369 -40800 -3369 -40752
rect -3050 -34848 2950 -34800
rect -3050 -40752 -3002 -34848
rect 2902 -40752 2950 -34848
rect -3050 -40800 2950 -40752
rect 3269 -34848 9269 -34800
rect 3269 -40752 3317 -34848
rect 9221 -40752 9269 -34848
rect 3269 -40800 9269 -40752
rect 9588 -34848 15588 -34800
rect 9588 -40752 9636 -34848
rect 15540 -40752 15588 -34848
rect 9588 -40800 15588 -40752
rect 15907 -34848 21907 -34800
rect 15907 -40752 15955 -34848
rect 21859 -40752 21907 -34848
rect 15907 -40800 21907 -40752
rect 22226 -34848 28226 -34800
rect 22226 -40752 22274 -34848
rect 28178 -40752 28226 -34848
rect 22226 -40800 28226 -40752
rect 28545 -34848 34545 -34800
rect 28545 -40752 28593 -34848
rect 34497 -40752 34545 -34848
rect 28545 -40800 34545 -40752
rect 34864 -34848 40864 -34800
rect 34864 -40752 34912 -34848
rect 40816 -40752 40864 -34848
rect 34864 -40800 40864 -40752
rect 41183 -34848 47183 -34800
rect 41183 -40752 41231 -34848
rect 47135 -40752 47183 -34848
rect 41183 -40800 47183 -40752
rect -47283 -41148 -41283 -41100
rect -47283 -47052 -47235 -41148
rect -41331 -47052 -41283 -41148
rect -47283 -47100 -41283 -47052
rect -40964 -41148 -34964 -41100
rect -40964 -47052 -40916 -41148
rect -35012 -47052 -34964 -41148
rect -40964 -47100 -34964 -47052
rect -34645 -41148 -28645 -41100
rect -34645 -47052 -34597 -41148
rect -28693 -47052 -28645 -41148
rect -34645 -47100 -28645 -47052
rect -28326 -41148 -22326 -41100
rect -28326 -47052 -28278 -41148
rect -22374 -47052 -22326 -41148
rect -28326 -47100 -22326 -47052
rect -22007 -41148 -16007 -41100
rect -22007 -47052 -21959 -41148
rect -16055 -47052 -16007 -41148
rect -22007 -47100 -16007 -47052
rect -15688 -41148 -9688 -41100
rect -15688 -47052 -15640 -41148
rect -9736 -47052 -9688 -41148
rect -15688 -47100 -9688 -47052
rect -9369 -41148 -3369 -41100
rect -9369 -47052 -9321 -41148
rect -3417 -47052 -3369 -41148
rect -9369 -47100 -3369 -47052
rect -3050 -41148 2950 -41100
rect -3050 -47052 -3002 -41148
rect 2902 -47052 2950 -41148
rect -3050 -47100 2950 -47052
rect 3269 -41148 9269 -41100
rect 3269 -47052 3317 -41148
rect 9221 -47052 9269 -41148
rect 3269 -47100 9269 -47052
rect 9588 -41148 15588 -41100
rect 9588 -47052 9636 -41148
rect 15540 -47052 15588 -41148
rect 9588 -47100 15588 -47052
rect 15907 -41148 21907 -41100
rect 15907 -47052 15955 -41148
rect 21859 -47052 21907 -41148
rect 15907 -47100 21907 -47052
rect 22226 -41148 28226 -41100
rect 22226 -47052 22274 -41148
rect 28178 -47052 28226 -41148
rect 22226 -47100 28226 -47052
rect 28545 -41148 34545 -41100
rect 28545 -47052 28593 -41148
rect 34497 -47052 34545 -41148
rect 28545 -47100 34545 -47052
rect 34864 -41148 40864 -41100
rect 34864 -47052 34912 -41148
rect 40816 -47052 40864 -41148
rect 34864 -47100 40864 -47052
rect 41183 -41148 47183 -41100
rect 41183 -47052 41231 -41148
rect 47135 -47052 47183 -41148
rect 41183 -47100 47183 -47052
<< mimcapcontact >>
rect -47235 41148 -41331 47052
rect -40916 41148 -35012 47052
rect -34597 41148 -28693 47052
rect -28278 41148 -22374 47052
rect -21959 41148 -16055 47052
rect -15640 41148 -9736 47052
rect -9321 41148 -3417 47052
rect -3002 41148 2902 47052
rect 3317 41148 9221 47052
rect 9636 41148 15540 47052
rect 15955 41148 21859 47052
rect 22274 41148 28178 47052
rect 28593 41148 34497 47052
rect 34912 41148 40816 47052
rect 41231 41148 47135 47052
rect -47235 34848 -41331 40752
rect -40916 34848 -35012 40752
rect -34597 34848 -28693 40752
rect -28278 34848 -22374 40752
rect -21959 34848 -16055 40752
rect -15640 34848 -9736 40752
rect -9321 34848 -3417 40752
rect -3002 34848 2902 40752
rect 3317 34848 9221 40752
rect 9636 34848 15540 40752
rect 15955 34848 21859 40752
rect 22274 34848 28178 40752
rect 28593 34848 34497 40752
rect 34912 34848 40816 40752
rect 41231 34848 47135 40752
rect -47235 28548 -41331 34452
rect -40916 28548 -35012 34452
rect -34597 28548 -28693 34452
rect -28278 28548 -22374 34452
rect -21959 28548 -16055 34452
rect -15640 28548 -9736 34452
rect -9321 28548 -3417 34452
rect -3002 28548 2902 34452
rect 3317 28548 9221 34452
rect 9636 28548 15540 34452
rect 15955 28548 21859 34452
rect 22274 28548 28178 34452
rect 28593 28548 34497 34452
rect 34912 28548 40816 34452
rect 41231 28548 47135 34452
rect -47235 22248 -41331 28152
rect -40916 22248 -35012 28152
rect -34597 22248 -28693 28152
rect -28278 22248 -22374 28152
rect -21959 22248 -16055 28152
rect -15640 22248 -9736 28152
rect -9321 22248 -3417 28152
rect -3002 22248 2902 28152
rect 3317 22248 9221 28152
rect 9636 22248 15540 28152
rect 15955 22248 21859 28152
rect 22274 22248 28178 28152
rect 28593 22248 34497 28152
rect 34912 22248 40816 28152
rect 41231 22248 47135 28152
rect -47235 15948 -41331 21852
rect -40916 15948 -35012 21852
rect -34597 15948 -28693 21852
rect -28278 15948 -22374 21852
rect -21959 15948 -16055 21852
rect -15640 15948 -9736 21852
rect -9321 15948 -3417 21852
rect -3002 15948 2902 21852
rect 3317 15948 9221 21852
rect 9636 15948 15540 21852
rect 15955 15948 21859 21852
rect 22274 15948 28178 21852
rect 28593 15948 34497 21852
rect 34912 15948 40816 21852
rect 41231 15948 47135 21852
rect -47235 9648 -41331 15552
rect -40916 9648 -35012 15552
rect -34597 9648 -28693 15552
rect -28278 9648 -22374 15552
rect -21959 9648 -16055 15552
rect -15640 9648 -9736 15552
rect -9321 9648 -3417 15552
rect -3002 9648 2902 15552
rect 3317 9648 9221 15552
rect 9636 9648 15540 15552
rect 15955 9648 21859 15552
rect 22274 9648 28178 15552
rect 28593 9648 34497 15552
rect 34912 9648 40816 15552
rect 41231 9648 47135 15552
rect -47235 3348 -41331 9252
rect -40916 3348 -35012 9252
rect -34597 3348 -28693 9252
rect -28278 3348 -22374 9252
rect -21959 3348 -16055 9252
rect -15640 3348 -9736 9252
rect -9321 3348 -3417 9252
rect -3002 3348 2902 9252
rect 3317 3348 9221 9252
rect 9636 3348 15540 9252
rect 15955 3348 21859 9252
rect 22274 3348 28178 9252
rect 28593 3348 34497 9252
rect 34912 3348 40816 9252
rect 41231 3348 47135 9252
rect -47235 -2952 -41331 2952
rect -40916 -2952 -35012 2952
rect -34597 -2952 -28693 2952
rect -28278 -2952 -22374 2952
rect -21959 -2952 -16055 2952
rect -15640 -2952 -9736 2952
rect -9321 -2952 -3417 2952
rect -3002 -2952 2902 2952
rect 3317 -2952 9221 2952
rect 9636 -2952 15540 2952
rect 15955 -2952 21859 2952
rect 22274 -2952 28178 2952
rect 28593 -2952 34497 2952
rect 34912 -2952 40816 2952
rect 41231 -2952 47135 2952
rect -47235 -9252 -41331 -3348
rect -40916 -9252 -35012 -3348
rect -34597 -9252 -28693 -3348
rect -28278 -9252 -22374 -3348
rect -21959 -9252 -16055 -3348
rect -15640 -9252 -9736 -3348
rect -9321 -9252 -3417 -3348
rect -3002 -9252 2902 -3348
rect 3317 -9252 9221 -3348
rect 9636 -9252 15540 -3348
rect 15955 -9252 21859 -3348
rect 22274 -9252 28178 -3348
rect 28593 -9252 34497 -3348
rect 34912 -9252 40816 -3348
rect 41231 -9252 47135 -3348
rect -47235 -15552 -41331 -9648
rect -40916 -15552 -35012 -9648
rect -34597 -15552 -28693 -9648
rect -28278 -15552 -22374 -9648
rect -21959 -15552 -16055 -9648
rect -15640 -15552 -9736 -9648
rect -9321 -15552 -3417 -9648
rect -3002 -15552 2902 -9648
rect 3317 -15552 9221 -9648
rect 9636 -15552 15540 -9648
rect 15955 -15552 21859 -9648
rect 22274 -15552 28178 -9648
rect 28593 -15552 34497 -9648
rect 34912 -15552 40816 -9648
rect 41231 -15552 47135 -9648
rect -47235 -21852 -41331 -15948
rect -40916 -21852 -35012 -15948
rect -34597 -21852 -28693 -15948
rect -28278 -21852 -22374 -15948
rect -21959 -21852 -16055 -15948
rect -15640 -21852 -9736 -15948
rect -9321 -21852 -3417 -15948
rect -3002 -21852 2902 -15948
rect 3317 -21852 9221 -15948
rect 9636 -21852 15540 -15948
rect 15955 -21852 21859 -15948
rect 22274 -21852 28178 -15948
rect 28593 -21852 34497 -15948
rect 34912 -21852 40816 -15948
rect 41231 -21852 47135 -15948
rect -47235 -28152 -41331 -22248
rect -40916 -28152 -35012 -22248
rect -34597 -28152 -28693 -22248
rect -28278 -28152 -22374 -22248
rect -21959 -28152 -16055 -22248
rect -15640 -28152 -9736 -22248
rect -9321 -28152 -3417 -22248
rect -3002 -28152 2902 -22248
rect 3317 -28152 9221 -22248
rect 9636 -28152 15540 -22248
rect 15955 -28152 21859 -22248
rect 22274 -28152 28178 -22248
rect 28593 -28152 34497 -22248
rect 34912 -28152 40816 -22248
rect 41231 -28152 47135 -22248
rect -47235 -34452 -41331 -28548
rect -40916 -34452 -35012 -28548
rect -34597 -34452 -28693 -28548
rect -28278 -34452 -22374 -28548
rect -21959 -34452 -16055 -28548
rect -15640 -34452 -9736 -28548
rect -9321 -34452 -3417 -28548
rect -3002 -34452 2902 -28548
rect 3317 -34452 9221 -28548
rect 9636 -34452 15540 -28548
rect 15955 -34452 21859 -28548
rect 22274 -34452 28178 -28548
rect 28593 -34452 34497 -28548
rect 34912 -34452 40816 -28548
rect 41231 -34452 47135 -28548
rect -47235 -40752 -41331 -34848
rect -40916 -40752 -35012 -34848
rect -34597 -40752 -28693 -34848
rect -28278 -40752 -22374 -34848
rect -21959 -40752 -16055 -34848
rect -15640 -40752 -9736 -34848
rect -9321 -40752 -3417 -34848
rect -3002 -40752 2902 -34848
rect 3317 -40752 9221 -34848
rect 9636 -40752 15540 -34848
rect 15955 -40752 21859 -34848
rect 22274 -40752 28178 -34848
rect 28593 -40752 34497 -34848
rect 34912 -40752 40816 -34848
rect 41231 -40752 47135 -34848
rect -47235 -47052 -41331 -41148
rect -40916 -47052 -35012 -41148
rect -34597 -47052 -28693 -41148
rect -28278 -47052 -22374 -41148
rect -21959 -47052 -16055 -41148
rect -15640 -47052 -9736 -41148
rect -9321 -47052 -3417 -41148
rect -3002 -47052 2902 -41148
rect 3317 -47052 9221 -41148
rect 9636 -47052 15540 -41148
rect 15955 -47052 21859 -41148
rect 22274 -47052 28178 -41148
rect 28593 -47052 34497 -41148
rect 34912 -47052 40816 -41148
rect 41231 -47052 47135 -41148
<< metal4 >>
rect -44335 47061 -44231 47250
rect -41215 47188 -41111 47250
rect -41215 47172 -41088 47188
rect -41215 47108 -41168 47172
rect -41104 47108 -41088 47172
rect -41215 47092 -41088 47108
rect -47244 47052 -41322 47061
rect -47244 41148 -47235 47052
rect -41331 41148 -41322 47052
rect -47244 41139 -41322 41148
rect -41215 47028 -41168 47092
rect -41104 47028 -41088 47092
rect -38016 47061 -37912 47250
rect -34896 47188 -34792 47250
rect -34896 47172 -34769 47188
rect -34896 47108 -34849 47172
rect -34785 47108 -34769 47172
rect -34896 47092 -34769 47108
rect -41215 47012 -41088 47028
rect -41215 46948 -41168 47012
rect -41104 46948 -41088 47012
rect -41215 46932 -41088 46948
rect -41215 46868 -41168 46932
rect -41104 46868 -41088 46932
rect -41215 46852 -41088 46868
rect -41215 46788 -41168 46852
rect -41104 46788 -41088 46852
rect -41215 46772 -41088 46788
rect -41215 46708 -41168 46772
rect -41104 46708 -41088 46772
rect -41215 46692 -41088 46708
rect -41215 46628 -41168 46692
rect -41104 46628 -41088 46692
rect -41215 46612 -41088 46628
rect -41215 46548 -41168 46612
rect -41104 46548 -41088 46612
rect -41215 46532 -41088 46548
rect -41215 46468 -41168 46532
rect -41104 46468 -41088 46532
rect -41215 46452 -41088 46468
rect -41215 46388 -41168 46452
rect -41104 46388 -41088 46452
rect -41215 46372 -41088 46388
rect -41215 46308 -41168 46372
rect -41104 46308 -41088 46372
rect -41215 46292 -41088 46308
rect -41215 46228 -41168 46292
rect -41104 46228 -41088 46292
rect -41215 46212 -41088 46228
rect -41215 46148 -41168 46212
rect -41104 46148 -41088 46212
rect -41215 46132 -41088 46148
rect -41215 46068 -41168 46132
rect -41104 46068 -41088 46132
rect -41215 46052 -41088 46068
rect -41215 45988 -41168 46052
rect -41104 45988 -41088 46052
rect -41215 45972 -41088 45988
rect -41215 45908 -41168 45972
rect -41104 45908 -41088 45972
rect -41215 45892 -41088 45908
rect -41215 45828 -41168 45892
rect -41104 45828 -41088 45892
rect -41215 45812 -41088 45828
rect -41215 45748 -41168 45812
rect -41104 45748 -41088 45812
rect -41215 45732 -41088 45748
rect -41215 45668 -41168 45732
rect -41104 45668 -41088 45732
rect -41215 45652 -41088 45668
rect -41215 45588 -41168 45652
rect -41104 45588 -41088 45652
rect -41215 45572 -41088 45588
rect -41215 45508 -41168 45572
rect -41104 45508 -41088 45572
rect -41215 45492 -41088 45508
rect -41215 45428 -41168 45492
rect -41104 45428 -41088 45492
rect -41215 45412 -41088 45428
rect -41215 45348 -41168 45412
rect -41104 45348 -41088 45412
rect -41215 45332 -41088 45348
rect -41215 45268 -41168 45332
rect -41104 45268 -41088 45332
rect -41215 45252 -41088 45268
rect -41215 45188 -41168 45252
rect -41104 45188 -41088 45252
rect -41215 45172 -41088 45188
rect -41215 45108 -41168 45172
rect -41104 45108 -41088 45172
rect -41215 45092 -41088 45108
rect -41215 45028 -41168 45092
rect -41104 45028 -41088 45092
rect -41215 45012 -41088 45028
rect -41215 44948 -41168 45012
rect -41104 44948 -41088 45012
rect -41215 44932 -41088 44948
rect -41215 44868 -41168 44932
rect -41104 44868 -41088 44932
rect -41215 44852 -41088 44868
rect -41215 44788 -41168 44852
rect -41104 44788 -41088 44852
rect -41215 44772 -41088 44788
rect -41215 44708 -41168 44772
rect -41104 44708 -41088 44772
rect -41215 44692 -41088 44708
rect -41215 44628 -41168 44692
rect -41104 44628 -41088 44692
rect -41215 44612 -41088 44628
rect -41215 44548 -41168 44612
rect -41104 44548 -41088 44612
rect -41215 44532 -41088 44548
rect -41215 44468 -41168 44532
rect -41104 44468 -41088 44532
rect -41215 44452 -41088 44468
rect -41215 44388 -41168 44452
rect -41104 44388 -41088 44452
rect -41215 44372 -41088 44388
rect -41215 44308 -41168 44372
rect -41104 44308 -41088 44372
rect -41215 44292 -41088 44308
rect -41215 44228 -41168 44292
rect -41104 44228 -41088 44292
rect -41215 44212 -41088 44228
rect -41215 44148 -41168 44212
rect -41104 44148 -41088 44212
rect -41215 44132 -41088 44148
rect -41215 44068 -41168 44132
rect -41104 44068 -41088 44132
rect -41215 44052 -41088 44068
rect -41215 43988 -41168 44052
rect -41104 43988 -41088 44052
rect -41215 43972 -41088 43988
rect -41215 43908 -41168 43972
rect -41104 43908 -41088 43972
rect -41215 43892 -41088 43908
rect -41215 43828 -41168 43892
rect -41104 43828 -41088 43892
rect -41215 43812 -41088 43828
rect -41215 43748 -41168 43812
rect -41104 43748 -41088 43812
rect -41215 43732 -41088 43748
rect -41215 43668 -41168 43732
rect -41104 43668 -41088 43732
rect -41215 43652 -41088 43668
rect -41215 43588 -41168 43652
rect -41104 43588 -41088 43652
rect -41215 43572 -41088 43588
rect -41215 43508 -41168 43572
rect -41104 43508 -41088 43572
rect -41215 43492 -41088 43508
rect -41215 43428 -41168 43492
rect -41104 43428 -41088 43492
rect -41215 43412 -41088 43428
rect -41215 43348 -41168 43412
rect -41104 43348 -41088 43412
rect -41215 43332 -41088 43348
rect -41215 43268 -41168 43332
rect -41104 43268 -41088 43332
rect -41215 43252 -41088 43268
rect -41215 43188 -41168 43252
rect -41104 43188 -41088 43252
rect -41215 43172 -41088 43188
rect -41215 43108 -41168 43172
rect -41104 43108 -41088 43172
rect -41215 43092 -41088 43108
rect -41215 43028 -41168 43092
rect -41104 43028 -41088 43092
rect -41215 43012 -41088 43028
rect -41215 42948 -41168 43012
rect -41104 42948 -41088 43012
rect -41215 42932 -41088 42948
rect -41215 42868 -41168 42932
rect -41104 42868 -41088 42932
rect -41215 42852 -41088 42868
rect -41215 42788 -41168 42852
rect -41104 42788 -41088 42852
rect -41215 42772 -41088 42788
rect -41215 42708 -41168 42772
rect -41104 42708 -41088 42772
rect -41215 42692 -41088 42708
rect -41215 42628 -41168 42692
rect -41104 42628 -41088 42692
rect -41215 42612 -41088 42628
rect -41215 42548 -41168 42612
rect -41104 42548 -41088 42612
rect -41215 42532 -41088 42548
rect -41215 42468 -41168 42532
rect -41104 42468 -41088 42532
rect -41215 42452 -41088 42468
rect -41215 42388 -41168 42452
rect -41104 42388 -41088 42452
rect -41215 42372 -41088 42388
rect -41215 42308 -41168 42372
rect -41104 42308 -41088 42372
rect -41215 42292 -41088 42308
rect -41215 42228 -41168 42292
rect -41104 42228 -41088 42292
rect -41215 42212 -41088 42228
rect -41215 42148 -41168 42212
rect -41104 42148 -41088 42212
rect -41215 42132 -41088 42148
rect -41215 42068 -41168 42132
rect -41104 42068 -41088 42132
rect -41215 42052 -41088 42068
rect -41215 41988 -41168 42052
rect -41104 41988 -41088 42052
rect -41215 41972 -41088 41988
rect -41215 41908 -41168 41972
rect -41104 41908 -41088 41972
rect -41215 41892 -41088 41908
rect -41215 41828 -41168 41892
rect -41104 41828 -41088 41892
rect -41215 41812 -41088 41828
rect -41215 41748 -41168 41812
rect -41104 41748 -41088 41812
rect -41215 41732 -41088 41748
rect -41215 41668 -41168 41732
rect -41104 41668 -41088 41732
rect -41215 41652 -41088 41668
rect -41215 41588 -41168 41652
rect -41104 41588 -41088 41652
rect -41215 41572 -41088 41588
rect -41215 41508 -41168 41572
rect -41104 41508 -41088 41572
rect -41215 41492 -41088 41508
rect -41215 41428 -41168 41492
rect -41104 41428 -41088 41492
rect -41215 41412 -41088 41428
rect -41215 41348 -41168 41412
rect -41104 41348 -41088 41412
rect -41215 41332 -41088 41348
rect -41215 41268 -41168 41332
rect -41104 41268 -41088 41332
rect -41215 41252 -41088 41268
rect -41215 41188 -41168 41252
rect -41104 41188 -41088 41252
rect -41215 41172 -41088 41188
rect -44335 40761 -44231 41139
rect -41215 41108 -41168 41172
rect -41104 41108 -41088 41172
rect -40925 47052 -35003 47061
rect -40925 41148 -40916 47052
rect -35012 41148 -35003 47052
rect -40925 41139 -35003 41148
rect -34896 47028 -34849 47092
rect -34785 47028 -34769 47092
rect -31697 47061 -31593 47250
rect -28577 47188 -28473 47250
rect -28577 47172 -28450 47188
rect -28577 47108 -28530 47172
rect -28466 47108 -28450 47172
rect -28577 47092 -28450 47108
rect -34896 47012 -34769 47028
rect -34896 46948 -34849 47012
rect -34785 46948 -34769 47012
rect -34896 46932 -34769 46948
rect -34896 46868 -34849 46932
rect -34785 46868 -34769 46932
rect -34896 46852 -34769 46868
rect -34896 46788 -34849 46852
rect -34785 46788 -34769 46852
rect -34896 46772 -34769 46788
rect -34896 46708 -34849 46772
rect -34785 46708 -34769 46772
rect -34896 46692 -34769 46708
rect -34896 46628 -34849 46692
rect -34785 46628 -34769 46692
rect -34896 46612 -34769 46628
rect -34896 46548 -34849 46612
rect -34785 46548 -34769 46612
rect -34896 46532 -34769 46548
rect -34896 46468 -34849 46532
rect -34785 46468 -34769 46532
rect -34896 46452 -34769 46468
rect -34896 46388 -34849 46452
rect -34785 46388 -34769 46452
rect -34896 46372 -34769 46388
rect -34896 46308 -34849 46372
rect -34785 46308 -34769 46372
rect -34896 46292 -34769 46308
rect -34896 46228 -34849 46292
rect -34785 46228 -34769 46292
rect -34896 46212 -34769 46228
rect -34896 46148 -34849 46212
rect -34785 46148 -34769 46212
rect -34896 46132 -34769 46148
rect -34896 46068 -34849 46132
rect -34785 46068 -34769 46132
rect -34896 46052 -34769 46068
rect -34896 45988 -34849 46052
rect -34785 45988 -34769 46052
rect -34896 45972 -34769 45988
rect -34896 45908 -34849 45972
rect -34785 45908 -34769 45972
rect -34896 45892 -34769 45908
rect -34896 45828 -34849 45892
rect -34785 45828 -34769 45892
rect -34896 45812 -34769 45828
rect -34896 45748 -34849 45812
rect -34785 45748 -34769 45812
rect -34896 45732 -34769 45748
rect -34896 45668 -34849 45732
rect -34785 45668 -34769 45732
rect -34896 45652 -34769 45668
rect -34896 45588 -34849 45652
rect -34785 45588 -34769 45652
rect -34896 45572 -34769 45588
rect -34896 45508 -34849 45572
rect -34785 45508 -34769 45572
rect -34896 45492 -34769 45508
rect -34896 45428 -34849 45492
rect -34785 45428 -34769 45492
rect -34896 45412 -34769 45428
rect -34896 45348 -34849 45412
rect -34785 45348 -34769 45412
rect -34896 45332 -34769 45348
rect -34896 45268 -34849 45332
rect -34785 45268 -34769 45332
rect -34896 45252 -34769 45268
rect -34896 45188 -34849 45252
rect -34785 45188 -34769 45252
rect -34896 45172 -34769 45188
rect -34896 45108 -34849 45172
rect -34785 45108 -34769 45172
rect -34896 45092 -34769 45108
rect -34896 45028 -34849 45092
rect -34785 45028 -34769 45092
rect -34896 45012 -34769 45028
rect -34896 44948 -34849 45012
rect -34785 44948 -34769 45012
rect -34896 44932 -34769 44948
rect -34896 44868 -34849 44932
rect -34785 44868 -34769 44932
rect -34896 44852 -34769 44868
rect -34896 44788 -34849 44852
rect -34785 44788 -34769 44852
rect -34896 44772 -34769 44788
rect -34896 44708 -34849 44772
rect -34785 44708 -34769 44772
rect -34896 44692 -34769 44708
rect -34896 44628 -34849 44692
rect -34785 44628 -34769 44692
rect -34896 44612 -34769 44628
rect -34896 44548 -34849 44612
rect -34785 44548 -34769 44612
rect -34896 44532 -34769 44548
rect -34896 44468 -34849 44532
rect -34785 44468 -34769 44532
rect -34896 44452 -34769 44468
rect -34896 44388 -34849 44452
rect -34785 44388 -34769 44452
rect -34896 44372 -34769 44388
rect -34896 44308 -34849 44372
rect -34785 44308 -34769 44372
rect -34896 44292 -34769 44308
rect -34896 44228 -34849 44292
rect -34785 44228 -34769 44292
rect -34896 44212 -34769 44228
rect -34896 44148 -34849 44212
rect -34785 44148 -34769 44212
rect -34896 44132 -34769 44148
rect -34896 44068 -34849 44132
rect -34785 44068 -34769 44132
rect -34896 44052 -34769 44068
rect -34896 43988 -34849 44052
rect -34785 43988 -34769 44052
rect -34896 43972 -34769 43988
rect -34896 43908 -34849 43972
rect -34785 43908 -34769 43972
rect -34896 43892 -34769 43908
rect -34896 43828 -34849 43892
rect -34785 43828 -34769 43892
rect -34896 43812 -34769 43828
rect -34896 43748 -34849 43812
rect -34785 43748 -34769 43812
rect -34896 43732 -34769 43748
rect -34896 43668 -34849 43732
rect -34785 43668 -34769 43732
rect -34896 43652 -34769 43668
rect -34896 43588 -34849 43652
rect -34785 43588 -34769 43652
rect -34896 43572 -34769 43588
rect -34896 43508 -34849 43572
rect -34785 43508 -34769 43572
rect -34896 43492 -34769 43508
rect -34896 43428 -34849 43492
rect -34785 43428 -34769 43492
rect -34896 43412 -34769 43428
rect -34896 43348 -34849 43412
rect -34785 43348 -34769 43412
rect -34896 43332 -34769 43348
rect -34896 43268 -34849 43332
rect -34785 43268 -34769 43332
rect -34896 43252 -34769 43268
rect -34896 43188 -34849 43252
rect -34785 43188 -34769 43252
rect -34896 43172 -34769 43188
rect -34896 43108 -34849 43172
rect -34785 43108 -34769 43172
rect -34896 43092 -34769 43108
rect -34896 43028 -34849 43092
rect -34785 43028 -34769 43092
rect -34896 43012 -34769 43028
rect -34896 42948 -34849 43012
rect -34785 42948 -34769 43012
rect -34896 42932 -34769 42948
rect -34896 42868 -34849 42932
rect -34785 42868 -34769 42932
rect -34896 42852 -34769 42868
rect -34896 42788 -34849 42852
rect -34785 42788 -34769 42852
rect -34896 42772 -34769 42788
rect -34896 42708 -34849 42772
rect -34785 42708 -34769 42772
rect -34896 42692 -34769 42708
rect -34896 42628 -34849 42692
rect -34785 42628 -34769 42692
rect -34896 42612 -34769 42628
rect -34896 42548 -34849 42612
rect -34785 42548 -34769 42612
rect -34896 42532 -34769 42548
rect -34896 42468 -34849 42532
rect -34785 42468 -34769 42532
rect -34896 42452 -34769 42468
rect -34896 42388 -34849 42452
rect -34785 42388 -34769 42452
rect -34896 42372 -34769 42388
rect -34896 42308 -34849 42372
rect -34785 42308 -34769 42372
rect -34896 42292 -34769 42308
rect -34896 42228 -34849 42292
rect -34785 42228 -34769 42292
rect -34896 42212 -34769 42228
rect -34896 42148 -34849 42212
rect -34785 42148 -34769 42212
rect -34896 42132 -34769 42148
rect -34896 42068 -34849 42132
rect -34785 42068 -34769 42132
rect -34896 42052 -34769 42068
rect -34896 41988 -34849 42052
rect -34785 41988 -34769 42052
rect -34896 41972 -34769 41988
rect -34896 41908 -34849 41972
rect -34785 41908 -34769 41972
rect -34896 41892 -34769 41908
rect -34896 41828 -34849 41892
rect -34785 41828 -34769 41892
rect -34896 41812 -34769 41828
rect -34896 41748 -34849 41812
rect -34785 41748 -34769 41812
rect -34896 41732 -34769 41748
rect -34896 41668 -34849 41732
rect -34785 41668 -34769 41732
rect -34896 41652 -34769 41668
rect -34896 41588 -34849 41652
rect -34785 41588 -34769 41652
rect -34896 41572 -34769 41588
rect -34896 41508 -34849 41572
rect -34785 41508 -34769 41572
rect -34896 41492 -34769 41508
rect -34896 41428 -34849 41492
rect -34785 41428 -34769 41492
rect -34896 41412 -34769 41428
rect -34896 41348 -34849 41412
rect -34785 41348 -34769 41412
rect -34896 41332 -34769 41348
rect -34896 41268 -34849 41332
rect -34785 41268 -34769 41332
rect -34896 41252 -34769 41268
rect -34896 41188 -34849 41252
rect -34785 41188 -34769 41252
rect -34896 41172 -34769 41188
rect -41215 41092 -41088 41108
rect -41215 41028 -41168 41092
rect -41104 41028 -41088 41092
rect -41215 41012 -41088 41028
rect -41215 40888 -41111 41012
rect -41215 40872 -41088 40888
rect -41215 40808 -41168 40872
rect -41104 40808 -41088 40872
rect -41215 40792 -41088 40808
rect -47244 40752 -41322 40761
rect -47244 34848 -47235 40752
rect -41331 34848 -41322 40752
rect -47244 34839 -41322 34848
rect -41215 40728 -41168 40792
rect -41104 40728 -41088 40792
rect -38016 40761 -37912 41139
rect -34896 41108 -34849 41172
rect -34785 41108 -34769 41172
rect -34606 47052 -28684 47061
rect -34606 41148 -34597 47052
rect -28693 41148 -28684 47052
rect -34606 41139 -28684 41148
rect -28577 47028 -28530 47092
rect -28466 47028 -28450 47092
rect -25378 47061 -25274 47250
rect -22258 47188 -22154 47250
rect -22258 47172 -22131 47188
rect -22258 47108 -22211 47172
rect -22147 47108 -22131 47172
rect -22258 47092 -22131 47108
rect -28577 47012 -28450 47028
rect -28577 46948 -28530 47012
rect -28466 46948 -28450 47012
rect -28577 46932 -28450 46948
rect -28577 46868 -28530 46932
rect -28466 46868 -28450 46932
rect -28577 46852 -28450 46868
rect -28577 46788 -28530 46852
rect -28466 46788 -28450 46852
rect -28577 46772 -28450 46788
rect -28577 46708 -28530 46772
rect -28466 46708 -28450 46772
rect -28577 46692 -28450 46708
rect -28577 46628 -28530 46692
rect -28466 46628 -28450 46692
rect -28577 46612 -28450 46628
rect -28577 46548 -28530 46612
rect -28466 46548 -28450 46612
rect -28577 46532 -28450 46548
rect -28577 46468 -28530 46532
rect -28466 46468 -28450 46532
rect -28577 46452 -28450 46468
rect -28577 46388 -28530 46452
rect -28466 46388 -28450 46452
rect -28577 46372 -28450 46388
rect -28577 46308 -28530 46372
rect -28466 46308 -28450 46372
rect -28577 46292 -28450 46308
rect -28577 46228 -28530 46292
rect -28466 46228 -28450 46292
rect -28577 46212 -28450 46228
rect -28577 46148 -28530 46212
rect -28466 46148 -28450 46212
rect -28577 46132 -28450 46148
rect -28577 46068 -28530 46132
rect -28466 46068 -28450 46132
rect -28577 46052 -28450 46068
rect -28577 45988 -28530 46052
rect -28466 45988 -28450 46052
rect -28577 45972 -28450 45988
rect -28577 45908 -28530 45972
rect -28466 45908 -28450 45972
rect -28577 45892 -28450 45908
rect -28577 45828 -28530 45892
rect -28466 45828 -28450 45892
rect -28577 45812 -28450 45828
rect -28577 45748 -28530 45812
rect -28466 45748 -28450 45812
rect -28577 45732 -28450 45748
rect -28577 45668 -28530 45732
rect -28466 45668 -28450 45732
rect -28577 45652 -28450 45668
rect -28577 45588 -28530 45652
rect -28466 45588 -28450 45652
rect -28577 45572 -28450 45588
rect -28577 45508 -28530 45572
rect -28466 45508 -28450 45572
rect -28577 45492 -28450 45508
rect -28577 45428 -28530 45492
rect -28466 45428 -28450 45492
rect -28577 45412 -28450 45428
rect -28577 45348 -28530 45412
rect -28466 45348 -28450 45412
rect -28577 45332 -28450 45348
rect -28577 45268 -28530 45332
rect -28466 45268 -28450 45332
rect -28577 45252 -28450 45268
rect -28577 45188 -28530 45252
rect -28466 45188 -28450 45252
rect -28577 45172 -28450 45188
rect -28577 45108 -28530 45172
rect -28466 45108 -28450 45172
rect -28577 45092 -28450 45108
rect -28577 45028 -28530 45092
rect -28466 45028 -28450 45092
rect -28577 45012 -28450 45028
rect -28577 44948 -28530 45012
rect -28466 44948 -28450 45012
rect -28577 44932 -28450 44948
rect -28577 44868 -28530 44932
rect -28466 44868 -28450 44932
rect -28577 44852 -28450 44868
rect -28577 44788 -28530 44852
rect -28466 44788 -28450 44852
rect -28577 44772 -28450 44788
rect -28577 44708 -28530 44772
rect -28466 44708 -28450 44772
rect -28577 44692 -28450 44708
rect -28577 44628 -28530 44692
rect -28466 44628 -28450 44692
rect -28577 44612 -28450 44628
rect -28577 44548 -28530 44612
rect -28466 44548 -28450 44612
rect -28577 44532 -28450 44548
rect -28577 44468 -28530 44532
rect -28466 44468 -28450 44532
rect -28577 44452 -28450 44468
rect -28577 44388 -28530 44452
rect -28466 44388 -28450 44452
rect -28577 44372 -28450 44388
rect -28577 44308 -28530 44372
rect -28466 44308 -28450 44372
rect -28577 44292 -28450 44308
rect -28577 44228 -28530 44292
rect -28466 44228 -28450 44292
rect -28577 44212 -28450 44228
rect -28577 44148 -28530 44212
rect -28466 44148 -28450 44212
rect -28577 44132 -28450 44148
rect -28577 44068 -28530 44132
rect -28466 44068 -28450 44132
rect -28577 44052 -28450 44068
rect -28577 43988 -28530 44052
rect -28466 43988 -28450 44052
rect -28577 43972 -28450 43988
rect -28577 43908 -28530 43972
rect -28466 43908 -28450 43972
rect -28577 43892 -28450 43908
rect -28577 43828 -28530 43892
rect -28466 43828 -28450 43892
rect -28577 43812 -28450 43828
rect -28577 43748 -28530 43812
rect -28466 43748 -28450 43812
rect -28577 43732 -28450 43748
rect -28577 43668 -28530 43732
rect -28466 43668 -28450 43732
rect -28577 43652 -28450 43668
rect -28577 43588 -28530 43652
rect -28466 43588 -28450 43652
rect -28577 43572 -28450 43588
rect -28577 43508 -28530 43572
rect -28466 43508 -28450 43572
rect -28577 43492 -28450 43508
rect -28577 43428 -28530 43492
rect -28466 43428 -28450 43492
rect -28577 43412 -28450 43428
rect -28577 43348 -28530 43412
rect -28466 43348 -28450 43412
rect -28577 43332 -28450 43348
rect -28577 43268 -28530 43332
rect -28466 43268 -28450 43332
rect -28577 43252 -28450 43268
rect -28577 43188 -28530 43252
rect -28466 43188 -28450 43252
rect -28577 43172 -28450 43188
rect -28577 43108 -28530 43172
rect -28466 43108 -28450 43172
rect -28577 43092 -28450 43108
rect -28577 43028 -28530 43092
rect -28466 43028 -28450 43092
rect -28577 43012 -28450 43028
rect -28577 42948 -28530 43012
rect -28466 42948 -28450 43012
rect -28577 42932 -28450 42948
rect -28577 42868 -28530 42932
rect -28466 42868 -28450 42932
rect -28577 42852 -28450 42868
rect -28577 42788 -28530 42852
rect -28466 42788 -28450 42852
rect -28577 42772 -28450 42788
rect -28577 42708 -28530 42772
rect -28466 42708 -28450 42772
rect -28577 42692 -28450 42708
rect -28577 42628 -28530 42692
rect -28466 42628 -28450 42692
rect -28577 42612 -28450 42628
rect -28577 42548 -28530 42612
rect -28466 42548 -28450 42612
rect -28577 42532 -28450 42548
rect -28577 42468 -28530 42532
rect -28466 42468 -28450 42532
rect -28577 42452 -28450 42468
rect -28577 42388 -28530 42452
rect -28466 42388 -28450 42452
rect -28577 42372 -28450 42388
rect -28577 42308 -28530 42372
rect -28466 42308 -28450 42372
rect -28577 42292 -28450 42308
rect -28577 42228 -28530 42292
rect -28466 42228 -28450 42292
rect -28577 42212 -28450 42228
rect -28577 42148 -28530 42212
rect -28466 42148 -28450 42212
rect -28577 42132 -28450 42148
rect -28577 42068 -28530 42132
rect -28466 42068 -28450 42132
rect -28577 42052 -28450 42068
rect -28577 41988 -28530 42052
rect -28466 41988 -28450 42052
rect -28577 41972 -28450 41988
rect -28577 41908 -28530 41972
rect -28466 41908 -28450 41972
rect -28577 41892 -28450 41908
rect -28577 41828 -28530 41892
rect -28466 41828 -28450 41892
rect -28577 41812 -28450 41828
rect -28577 41748 -28530 41812
rect -28466 41748 -28450 41812
rect -28577 41732 -28450 41748
rect -28577 41668 -28530 41732
rect -28466 41668 -28450 41732
rect -28577 41652 -28450 41668
rect -28577 41588 -28530 41652
rect -28466 41588 -28450 41652
rect -28577 41572 -28450 41588
rect -28577 41508 -28530 41572
rect -28466 41508 -28450 41572
rect -28577 41492 -28450 41508
rect -28577 41428 -28530 41492
rect -28466 41428 -28450 41492
rect -28577 41412 -28450 41428
rect -28577 41348 -28530 41412
rect -28466 41348 -28450 41412
rect -28577 41332 -28450 41348
rect -28577 41268 -28530 41332
rect -28466 41268 -28450 41332
rect -28577 41252 -28450 41268
rect -28577 41188 -28530 41252
rect -28466 41188 -28450 41252
rect -28577 41172 -28450 41188
rect -34896 41092 -34769 41108
rect -34896 41028 -34849 41092
rect -34785 41028 -34769 41092
rect -34896 41012 -34769 41028
rect -34896 40888 -34792 41012
rect -34896 40872 -34769 40888
rect -34896 40808 -34849 40872
rect -34785 40808 -34769 40872
rect -34896 40792 -34769 40808
rect -41215 40712 -41088 40728
rect -41215 40648 -41168 40712
rect -41104 40648 -41088 40712
rect -41215 40632 -41088 40648
rect -41215 40568 -41168 40632
rect -41104 40568 -41088 40632
rect -41215 40552 -41088 40568
rect -41215 40488 -41168 40552
rect -41104 40488 -41088 40552
rect -41215 40472 -41088 40488
rect -41215 40408 -41168 40472
rect -41104 40408 -41088 40472
rect -41215 40392 -41088 40408
rect -41215 40328 -41168 40392
rect -41104 40328 -41088 40392
rect -41215 40312 -41088 40328
rect -41215 40248 -41168 40312
rect -41104 40248 -41088 40312
rect -41215 40232 -41088 40248
rect -41215 40168 -41168 40232
rect -41104 40168 -41088 40232
rect -41215 40152 -41088 40168
rect -41215 40088 -41168 40152
rect -41104 40088 -41088 40152
rect -41215 40072 -41088 40088
rect -41215 40008 -41168 40072
rect -41104 40008 -41088 40072
rect -41215 39992 -41088 40008
rect -41215 39928 -41168 39992
rect -41104 39928 -41088 39992
rect -41215 39912 -41088 39928
rect -41215 39848 -41168 39912
rect -41104 39848 -41088 39912
rect -41215 39832 -41088 39848
rect -41215 39768 -41168 39832
rect -41104 39768 -41088 39832
rect -41215 39752 -41088 39768
rect -41215 39688 -41168 39752
rect -41104 39688 -41088 39752
rect -41215 39672 -41088 39688
rect -41215 39608 -41168 39672
rect -41104 39608 -41088 39672
rect -41215 39592 -41088 39608
rect -41215 39528 -41168 39592
rect -41104 39528 -41088 39592
rect -41215 39512 -41088 39528
rect -41215 39448 -41168 39512
rect -41104 39448 -41088 39512
rect -41215 39432 -41088 39448
rect -41215 39368 -41168 39432
rect -41104 39368 -41088 39432
rect -41215 39352 -41088 39368
rect -41215 39288 -41168 39352
rect -41104 39288 -41088 39352
rect -41215 39272 -41088 39288
rect -41215 39208 -41168 39272
rect -41104 39208 -41088 39272
rect -41215 39192 -41088 39208
rect -41215 39128 -41168 39192
rect -41104 39128 -41088 39192
rect -41215 39112 -41088 39128
rect -41215 39048 -41168 39112
rect -41104 39048 -41088 39112
rect -41215 39032 -41088 39048
rect -41215 38968 -41168 39032
rect -41104 38968 -41088 39032
rect -41215 38952 -41088 38968
rect -41215 38888 -41168 38952
rect -41104 38888 -41088 38952
rect -41215 38872 -41088 38888
rect -41215 38808 -41168 38872
rect -41104 38808 -41088 38872
rect -41215 38792 -41088 38808
rect -41215 38728 -41168 38792
rect -41104 38728 -41088 38792
rect -41215 38712 -41088 38728
rect -41215 38648 -41168 38712
rect -41104 38648 -41088 38712
rect -41215 38632 -41088 38648
rect -41215 38568 -41168 38632
rect -41104 38568 -41088 38632
rect -41215 38552 -41088 38568
rect -41215 38488 -41168 38552
rect -41104 38488 -41088 38552
rect -41215 38472 -41088 38488
rect -41215 38408 -41168 38472
rect -41104 38408 -41088 38472
rect -41215 38392 -41088 38408
rect -41215 38328 -41168 38392
rect -41104 38328 -41088 38392
rect -41215 38312 -41088 38328
rect -41215 38248 -41168 38312
rect -41104 38248 -41088 38312
rect -41215 38232 -41088 38248
rect -41215 38168 -41168 38232
rect -41104 38168 -41088 38232
rect -41215 38152 -41088 38168
rect -41215 38088 -41168 38152
rect -41104 38088 -41088 38152
rect -41215 38072 -41088 38088
rect -41215 38008 -41168 38072
rect -41104 38008 -41088 38072
rect -41215 37992 -41088 38008
rect -41215 37928 -41168 37992
rect -41104 37928 -41088 37992
rect -41215 37912 -41088 37928
rect -41215 37848 -41168 37912
rect -41104 37848 -41088 37912
rect -41215 37832 -41088 37848
rect -41215 37768 -41168 37832
rect -41104 37768 -41088 37832
rect -41215 37752 -41088 37768
rect -41215 37688 -41168 37752
rect -41104 37688 -41088 37752
rect -41215 37672 -41088 37688
rect -41215 37608 -41168 37672
rect -41104 37608 -41088 37672
rect -41215 37592 -41088 37608
rect -41215 37528 -41168 37592
rect -41104 37528 -41088 37592
rect -41215 37512 -41088 37528
rect -41215 37448 -41168 37512
rect -41104 37448 -41088 37512
rect -41215 37432 -41088 37448
rect -41215 37368 -41168 37432
rect -41104 37368 -41088 37432
rect -41215 37352 -41088 37368
rect -41215 37288 -41168 37352
rect -41104 37288 -41088 37352
rect -41215 37272 -41088 37288
rect -41215 37208 -41168 37272
rect -41104 37208 -41088 37272
rect -41215 37192 -41088 37208
rect -41215 37128 -41168 37192
rect -41104 37128 -41088 37192
rect -41215 37112 -41088 37128
rect -41215 37048 -41168 37112
rect -41104 37048 -41088 37112
rect -41215 37032 -41088 37048
rect -41215 36968 -41168 37032
rect -41104 36968 -41088 37032
rect -41215 36952 -41088 36968
rect -41215 36888 -41168 36952
rect -41104 36888 -41088 36952
rect -41215 36872 -41088 36888
rect -41215 36808 -41168 36872
rect -41104 36808 -41088 36872
rect -41215 36792 -41088 36808
rect -41215 36728 -41168 36792
rect -41104 36728 -41088 36792
rect -41215 36712 -41088 36728
rect -41215 36648 -41168 36712
rect -41104 36648 -41088 36712
rect -41215 36632 -41088 36648
rect -41215 36568 -41168 36632
rect -41104 36568 -41088 36632
rect -41215 36552 -41088 36568
rect -41215 36488 -41168 36552
rect -41104 36488 -41088 36552
rect -41215 36472 -41088 36488
rect -41215 36408 -41168 36472
rect -41104 36408 -41088 36472
rect -41215 36392 -41088 36408
rect -41215 36328 -41168 36392
rect -41104 36328 -41088 36392
rect -41215 36312 -41088 36328
rect -41215 36248 -41168 36312
rect -41104 36248 -41088 36312
rect -41215 36232 -41088 36248
rect -41215 36168 -41168 36232
rect -41104 36168 -41088 36232
rect -41215 36152 -41088 36168
rect -41215 36088 -41168 36152
rect -41104 36088 -41088 36152
rect -41215 36072 -41088 36088
rect -41215 36008 -41168 36072
rect -41104 36008 -41088 36072
rect -41215 35992 -41088 36008
rect -41215 35928 -41168 35992
rect -41104 35928 -41088 35992
rect -41215 35912 -41088 35928
rect -41215 35848 -41168 35912
rect -41104 35848 -41088 35912
rect -41215 35832 -41088 35848
rect -41215 35768 -41168 35832
rect -41104 35768 -41088 35832
rect -41215 35752 -41088 35768
rect -41215 35688 -41168 35752
rect -41104 35688 -41088 35752
rect -41215 35672 -41088 35688
rect -41215 35608 -41168 35672
rect -41104 35608 -41088 35672
rect -41215 35592 -41088 35608
rect -41215 35528 -41168 35592
rect -41104 35528 -41088 35592
rect -41215 35512 -41088 35528
rect -41215 35448 -41168 35512
rect -41104 35448 -41088 35512
rect -41215 35432 -41088 35448
rect -41215 35368 -41168 35432
rect -41104 35368 -41088 35432
rect -41215 35352 -41088 35368
rect -41215 35288 -41168 35352
rect -41104 35288 -41088 35352
rect -41215 35272 -41088 35288
rect -41215 35208 -41168 35272
rect -41104 35208 -41088 35272
rect -41215 35192 -41088 35208
rect -41215 35128 -41168 35192
rect -41104 35128 -41088 35192
rect -41215 35112 -41088 35128
rect -41215 35048 -41168 35112
rect -41104 35048 -41088 35112
rect -41215 35032 -41088 35048
rect -41215 34968 -41168 35032
rect -41104 34968 -41088 35032
rect -41215 34952 -41088 34968
rect -41215 34888 -41168 34952
rect -41104 34888 -41088 34952
rect -41215 34872 -41088 34888
rect -44335 34461 -44231 34839
rect -41215 34808 -41168 34872
rect -41104 34808 -41088 34872
rect -40925 40752 -35003 40761
rect -40925 34848 -40916 40752
rect -35012 34848 -35003 40752
rect -40925 34839 -35003 34848
rect -34896 40728 -34849 40792
rect -34785 40728 -34769 40792
rect -31697 40761 -31593 41139
rect -28577 41108 -28530 41172
rect -28466 41108 -28450 41172
rect -28287 47052 -22365 47061
rect -28287 41148 -28278 47052
rect -22374 41148 -22365 47052
rect -28287 41139 -22365 41148
rect -22258 47028 -22211 47092
rect -22147 47028 -22131 47092
rect -19059 47061 -18955 47250
rect -15939 47188 -15835 47250
rect -15939 47172 -15812 47188
rect -15939 47108 -15892 47172
rect -15828 47108 -15812 47172
rect -15939 47092 -15812 47108
rect -22258 47012 -22131 47028
rect -22258 46948 -22211 47012
rect -22147 46948 -22131 47012
rect -22258 46932 -22131 46948
rect -22258 46868 -22211 46932
rect -22147 46868 -22131 46932
rect -22258 46852 -22131 46868
rect -22258 46788 -22211 46852
rect -22147 46788 -22131 46852
rect -22258 46772 -22131 46788
rect -22258 46708 -22211 46772
rect -22147 46708 -22131 46772
rect -22258 46692 -22131 46708
rect -22258 46628 -22211 46692
rect -22147 46628 -22131 46692
rect -22258 46612 -22131 46628
rect -22258 46548 -22211 46612
rect -22147 46548 -22131 46612
rect -22258 46532 -22131 46548
rect -22258 46468 -22211 46532
rect -22147 46468 -22131 46532
rect -22258 46452 -22131 46468
rect -22258 46388 -22211 46452
rect -22147 46388 -22131 46452
rect -22258 46372 -22131 46388
rect -22258 46308 -22211 46372
rect -22147 46308 -22131 46372
rect -22258 46292 -22131 46308
rect -22258 46228 -22211 46292
rect -22147 46228 -22131 46292
rect -22258 46212 -22131 46228
rect -22258 46148 -22211 46212
rect -22147 46148 -22131 46212
rect -22258 46132 -22131 46148
rect -22258 46068 -22211 46132
rect -22147 46068 -22131 46132
rect -22258 46052 -22131 46068
rect -22258 45988 -22211 46052
rect -22147 45988 -22131 46052
rect -22258 45972 -22131 45988
rect -22258 45908 -22211 45972
rect -22147 45908 -22131 45972
rect -22258 45892 -22131 45908
rect -22258 45828 -22211 45892
rect -22147 45828 -22131 45892
rect -22258 45812 -22131 45828
rect -22258 45748 -22211 45812
rect -22147 45748 -22131 45812
rect -22258 45732 -22131 45748
rect -22258 45668 -22211 45732
rect -22147 45668 -22131 45732
rect -22258 45652 -22131 45668
rect -22258 45588 -22211 45652
rect -22147 45588 -22131 45652
rect -22258 45572 -22131 45588
rect -22258 45508 -22211 45572
rect -22147 45508 -22131 45572
rect -22258 45492 -22131 45508
rect -22258 45428 -22211 45492
rect -22147 45428 -22131 45492
rect -22258 45412 -22131 45428
rect -22258 45348 -22211 45412
rect -22147 45348 -22131 45412
rect -22258 45332 -22131 45348
rect -22258 45268 -22211 45332
rect -22147 45268 -22131 45332
rect -22258 45252 -22131 45268
rect -22258 45188 -22211 45252
rect -22147 45188 -22131 45252
rect -22258 45172 -22131 45188
rect -22258 45108 -22211 45172
rect -22147 45108 -22131 45172
rect -22258 45092 -22131 45108
rect -22258 45028 -22211 45092
rect -22147 45028 -22131 45092
rect -22258 45012 -22131 45028
rect -22258 44948 -22211 45012
rect -22147 44948 -22131 45012
rect -22258 44932 -22131 44948
rect -22258 44868 -22211 44932
rect -22147 44868 -22131 44932
rect -22258 44852 -22131 44868
rect -22258 44788 -22211 44852
rect -22147 44788 -22131 44852
rect -22258 44772 -22131 44788
rect -22258 44708 -22211 44772
rect -22147 44708 -22131 44772
rect -22258 44692 -22131 44708
rect -22258 44628 -22211 44692
rect -22147 44628 -22131 44692
rect -22258 44612 -22131 44628
rect -22258 44548 -22211 44612
rect -22147 44548 -22131 44612
rect -22258 44532 -22131 44548
rect -22258 44468 -22211 44532
rect -22147 44468 -22131 44532
rect -22258 44452 -22131 44468
rect -22258 44388 -22211 44452
rect -22147 44388 -22131 44452
rect -22258 44372 -22131 44388
rect -22258 44308 -22211 44372
rect -22147 44308 -22131 44372
rect -22258 44292 -22131 44308
rect -22258 44228 -22211 44292
rect -22147 44228 -22131 44292
rect -22258 44212 -22131 44228
rect -22258 44148 -22211 44212
rect -22147 44148 -22131 44212
rect -22258 44132 -22131 44148
rect -22258 44068 -22211 44132
rect -22147 44068 -22131 44132
rect -22258 44052 -22131 44068
rect -22258 43988 -22211 44052
rect -22147 43988 -22131 44052
rect -22258 43972 -22131 43988
rect -22258 43908 -22211 43972
rect -22147 43908 -22131 43972
rect -22258 43892 -22131 43908
rect -22258 43828 -22211 43892
rect -22147 43828 -22131 43892
rect -22258 43812 -22131 43828
rect -22258 43748 -22211 43812
rect -22147 43748 -22131 43812
rect -22258 43732 -22131 43748
rect -22258 43668 -22211 43732
rect -22147 43668 -22131 43732
rect -22258 43652 -22131 43668
rect -22258 43588 -22211 43652
rect -22147 43588 -22131 43652
rect -22258 43572 -22131 43588
rect -22258 43508 -22211 43572
rect -22147 43508 -22131 43572
rect -22258 43492 -22131 43508
rect -22258 43428 -22211 43492
rect -22147 43428 -22131 43492
rect -22258 43412 -22131 43428
rect -22258 43348 -22211 43412
rect -22147 43348 -22131 43412
rect -22258 43332 -22131 43348
rect -22258 43268 -22211 43332
rect -22147 43268 -22131 43332
rect -22258 43252 -22131 43268
rect -22258 43188 -22211 43252
rect -22147 43188 -22131 43252
rect -22258 43172 -22131 43188
rect -22258 43108 -22211 43172
rect -22147 43108 -22131 43172
rect -22258 43092 -22131 43108
rect -22258 43028 -22211 43092
rect -22147 43028 -22131 43092
rect -22258 43012 -22131 43028
rect -22258 42948 -22211 43012
rect -22147 42948 -22131 43012
rect -22258 42932 -22131 42948
rect -22258 42868 -22211 42932
rect -22147 42868 -22131 42932
rect -22258 42852 -22131 42868
rect -22258 42788 -22211 42852
rect -22147 42788 -22131 42852
rect -22258 42772 -22131 42788
rect -22258 42708 -22211 42772
rect -22147 42708 -22131 42772
rect -22258 42692 -22131 42708
rect -22258 42628 -22211 42692
rect -22147 42628 -22131 42692
rect -22258 42612 -22131 42628
rect -22258 42548 -22211 42612
rect -22147 42548 -22131 42612
rect -22258 42532 -22131 42548
rect -22258 42468 -22211 42532
rect -22147 42468 -22131 42532
rect -22258 42452 -22131 42468
rect -22258 42388 -22211 42452
rect -22147 42388 -22131 42452
rect -22258 42372 -22131 42388
rect -22258 42308 -22211 42372
rect -22147 42308 -22131 42372
rect -22258 42292 -22131 42308
rect -22258 42228 -22211 42292
rect -22147 42228 -22131 42292
rect -22258 42212 -22131 42228
rect -22258 42148 -22211 42212
rect -22147 42148 -22131 42212
rect -22258 42132 -22131 42148
rect -22258 42068 -22211 42132
rect -22147 42068 -22131 42132
rect -22258 42052 -22131 42068
rect -22258 41988 -22211 42052
rect -22147 41988 -22131 42052
rect -22258 41972 -22131 41988
rect -22258 41908 -22211 41972
rect -22147 41908 -22131 41972
rect -22258 41892 -22131 41908
rect -22258 41828 -22211 41892
rect -22147 41828 -22131 41892
rect -22258 41812 -22131 41828
rect -22258 41748 -22211 41812
rect -22147 41748 -22131 41812
rect -22258 41732 -22131 41748
rect -22258 41668 -22211 41732
rect -22147 41668 -22131 41732
rect -22258 41652 -22131 41668
rect -22258 41588 -22211 41652
rect -22147 41588 -22131 41652
rect -22258 41572 -22131 41588
rect -22258 41508 -22211 41572
rect -22147 41508 -22131 41572
rect -22258 41492 -22131 41508
rect -22258 41428 -22211 41492
rect -22147 41428 -22131 41492
rect -22258 41412 -22131 41428
rect -22258 41348 -22211 41412
rect -22147 41348 -22131 41412
rect -22258 41332 -22131 41348
rect -22258 41268 -22211 41332
rect -22147 41268 -22131 41332
rect -22258 41252 -22131 41268
rect -22258 41188 -22211 41252
rect -22147 41188 -22131 41252
rect -22258 41172 -22131 41188
rect -28577 41092 -28450 41108
rect -28577 41028 -28530 41092
rect -28466 41028 -28450 41092
rect -28577 41012 -28450 41028
rect -28577 40888 -28473 41012
rect -28577 40872 -28450 40888
rect -28577 40808 -28530 40872
rect -28466 40808 -28450 40872
rect -28577 40792 -28450 40808
rect -34896 40712 -34769 40728
rect -34896 40648 -34849 40712
rect -34785 40648 -34769 40712
rect -34896 40632 -34769 40648
rect -34896 40568 -34849 40632
rect -34785 40568 -34769 40632
rect -34896 40552 -34769 40568
rect -34896 40488 -34849 40552
rect -34785 40488 -34769 40552
rect -34896 40472 -34769 40488
rect -34896 40408 -34849 40472
rect -34785 40408 -34769 40472
rect -34896 40392 -34769 40408
rect -34896 40328 -34849 40392
rect -34785 40328 -34769 40392
rect -34896 40312 -34769 40328
rect -34896 40248 -34849 40312
rect -34785 40248 -34769 40312
rect -34896 40232 -34769 40248
rect -34896 40168 -34849 40232
rect -34785 40168 -34769 40232
rect -34896 40152 -34769 40168
rect -34896 40088 -34849 40152
rect -34785 40088 -34769 40152
rect -34896 40072 -34769 40088
rect -34896 40008 -34849 40072
rect -34785 40008 -34769 40072
rect -34896 39992 -34769 40008
rect -34896 39928 -34849 39992
rect -34785 39928 -34769 39992
rect -34896 39912 -34769 39928
rect -34896 39848 -34849 39912
rect -34785 39848 -34769 39912
rect -34896 39832 -34769 39848
rect -34896 39768 -34849 39832
rect -34785 39768 -34769 39832
rect -34896 39752 -34769 39768
rect -34896 39688 -34849 39752
rect -34785 39688 -34769 39752
rect -34896 39672 -34769 39688
rect -34896 39608 -34849 39672
rect -34785 39608 -34769 39672
rect -34896 39592 -34769 39608
rect -34896 39528 -34849 39592
rect -34785 39528 -34769 39592
rect -34896 39512 -34769 39528
rect -34896 39448 -34849 39512
rect -34785 39448 -34769 39512
rect -34896 39432 -34769 39448
rect -34896 39368 -34849 39432
rect -34785 39368 -34769 39432
rect -34896 39352 -34769 39368
rect -34896 39288 -34849 39352
rect -34785 39288 -34769 39352
rect -34896 39272 -34769 39288
rect -34896 39208 -34849 39272
rect -34785 39208 -34769 39272
rect -34896 39192 -34769 39208
rect -34896 39128 -34849 39192
rect -34785 39128 -34769 39192
rect -34896 39112 -34769 39128
rect -34896 39048 -34849 39112
rect -34785 39048 -34769 39112
rect -34896 39032 -34769 39048
rect -34896 38968 -34849 39032
rect -34785 38968 -34769 39032
rect -34896 38952 -34769 38968
rect -34896 38888 -34849 38952
rect -34785 38888 -34769 38952
rect -34896 38872 -34769 38888
rect -34896 38808 -34849 38872
rect -34785 38808 -34769 38872
rect -34896 38792 -34769 38808
rect -34896 38728 -34849 38792
rect -34785 38728 -34769 38792
rect -34896 38712 -34769 38728
rect -34896 38648 -34849 38712
rect -34785 38648 -34769 38712
rect -34896 38632 -34769 38648
rect -34896 38568 -34849 38632
rect -34785 38568 -34769 38632
rect -34896 38552 -34769 38568
rect -34896 38488 -34849 38552
rect -34785 38488 -34769 38552
rect -34896 38472 -34769 38488
rect -34896 38408 -34849 38472
rect -34785 38408 -34769 38472
rect -34896 38392 -34769 38408
rect -34896 38328 -34849 38392
rect -34785 38328 -34769 38392
rect -34896 38312 -34769 38328
rect -34896 38248 -34849 38312
rect -34785 38248 -34769 38312
rect -34896 38232 -34769 38248
rect -34896 38168 -34849 38232
rect -34785 38168 -34769 38232
rect -34896 38152 -34769 38168
rect -34896 38088 -34849 38152
rect -34785 38088 -34769 38152
rect -34896 38072 -34769 38088
rect -34896 38008 -34849 38072
rect -34785 38008 -34769 38072
rect -34896 37992 -34769 38008
rect -34896 37928 -34849 37992
rect -34785 37928 -34769 37992
rect -34896 37912 -34769 37928
rect -34896 37848 -34849 37912
rect -34785 37848 -34769 37912
rect -34896 37832 -34769 37848
rect -34896 37768 -34849 37832
rect -34785 37768 -34769 37832
rect -34896 37752 -34769 37768
rect -34896 37688 -34849 37752
rect -34785 37688 -34769 37752
rect -34896 37672 -34769 37688
rect -34896 37608 -34849 37672
rect -34785 37608 -34769 37672
rect -34896 37592 -34769 37608
rect -34896 37528 -34849 37592
rect -34785 37528 -34769 37592
rect -34896 37512 -34769 37528
rect -34896 37448 -34849 37512
rect -34785 37448 -34769 37512
rect -34896 37432 -34769 37448
rect -34896 37368 -34849 37432
rect -34785 37368 -34769 37432
rect -34896 37352 -34769 37368
rect -34896 37288 -34849 37352
rect -34785 37288 -34769 37352
rect -34896 37272 -34769 37288
rect -34896 37208 -34849 37272
rect -34785 37208 -34769 37272
rect -34896 37192 -34769 37208
rect -34896 37128 -34849 37192
rect -34785 37128 -34769 37192
rect -34896 37112 -34769 37128
rect -34896 37048 -34849 37112
rect -34785 37048 -34769 37112
rect -34896 37032 -34769 37048
rect -34896 36968 -34849 37032
rect -34785 36968 -34769 37032
rect -34896 36952 -34769 36968
rect -34896 36888 -34849 36952
rect -34785 36888 -34769 36952
rect -34896 36872 -34769 36888
rect -34896 36808 -34849 36872
rect -34785 36808 -34769 36872
rect -34896 36792 -34769 36808
rect -34896 36728 -34849 36792
rect -34785 36728 -34769 36792
rect -34896 36712 -34769 36728
rect -34896 36648 -34849 36712
rect -34785 36648 -34769 36712
rect -34896 36632 -34769 36648
rect -34896 36568 -34849 36632
rect -34785 36568 -34769 36632
rect -34896 36552 -34769 36568
rect -34896 36488 -34849 36552
rect -34785 36488 -34769 36552
rect -34896 36472 -34769 36488
rect -34896 36408 -34849 36472
rect -34785 36408 -34769 36472
rect -34896 36392 -34769 36408
rect -34896 36328 -34849 36392
rect -34785 36328 -34769 36392
rect -34896 36312 -34769 36328
rect -34896 36248 -34849 36312
rect -34785 36248 -34769 36312
rect -34896 36232 -34769 36248
rect -34896 36168 -34849 36232
rect -34785 36168 -34769 36232
rect -34896 36152 -34769 36168
rect -34896 36088 -34849 36152
rect -34785 36088 -34769 36152
rect -34896 36072 -34769 36088
rect -34896 36008 -34849 36072
rect -34785 36008 -34769 36072
rect -34896 35992 -34769 36008
rect -34896 35928 -34849 35992
rect -34785 35928 -34769 35992
rect -34896 35912 -34769 35928
rect -34896 35848 -34849 35912
rect -34785 35848 -34769 35912
rect -34896 35832 -34769 35848
rect -34896 35768 -34849 35832
rect -34785 35768 -34769 35832
rect -34896 35752 -34769 35768
rect -34896 35688 -34849 35752
rect -34785 35688 -34769 35752
rect -34896 35672 -34769 35688
rect -34896 35608 -34849 35672
rect -34785 35608 -34769 35672
rect -34896 35592 -34769 35608
rect -34896 35528 -34849 35592
rect -34785 35528 -34769 35592
rect -34896 35512 -34769 35528
rect -34896 35448 -34849 35512
rect -34785 35448 -34769 35512
rect -34896 35432 -34769 35448
rect -34896 35368 -34849 35432
rect -34785 35368 -34769 35432
rect -34896 35352 -34769 35368
rect -34896 35288 -34849 35352
rect -34785 35288 -34769 35352
rect -34896 35272 -34769 35288
rect -34896 35208 -34849 35272
rect -34785 35208 -34769 35272
rect -34896 35192 -34769 35208
rect -34896 35128 -34849 35192
rect -34785 35128 -34769 35192
rect -34896 35112 -34769 35128
rect -34896 35048 -34849 35112
rect -34785 35048 -34769 35112
rect -34896 35032 -34769 35048
rect -34896 34968 -34849 35032
rect -34785 34968 -34769 35032
rect -34896 34952 -34769 34968
rect -34896 34888 -34849 34952
rect -34785 34888 -34769 34952
rect -34896 34872 -34769 34888
rect -41215 34792 -41088 34808
rect -41215 34728 -41168 34792
rect -41104 34728 -41088 34792
rect -41215 34712 -41088 34728
rect -41215 34588 -41111 34712
rect -41215 34572 -41088 34588
rect -41215 34508 -41168 34572
rect -41104 34508 -41088 34572
rect -41215 34492 -41088 34508
rect -47244 34452 -41322 34461
rect -47244 28548 -47235 34452
rect -41331 28548 -41322 34452
rect -47244 28539 -41322 28548
rect -41215 34428 -41168 34492
rect -41104 34428 -41088 34492
rect -38016 34461 -37912 34839
rect -34896 34808 -34849 34872
rect -34785 34808 -34769 34872
rect -34606 40752 -28684 40761
rect -34606 34848 -34597 40752
rect -28693 34848 -28684 40752
rect -34606 34839 -28684 34848
rect -28577 40728 -28530 40792
rect -28466 40728 -28450 40792
rect -25378 40761 -25274 41139
rect -22258 41108 -22211 41172
rect -22147 41108 -22131 41172
rect -21968 47052 -16046 47061
rect -21968 41148 -21959 47052
rect -16055 41148 -16046 47052
rect -21968 41139 -16046 41148
rect -15939 47028 -15892 47092
rect -15828 47028 -15812 47092
rect -12740 47061 -12636 47250
rect -9620 47188 -9516 47250
rect -9620 47172 -9493 47188
rect -9620 47108 -9573 47172
rect -9509 47108 -9493 47172
rect -9620 47092 -9493 47108
rect -15939 47012 -15812 47028
rect -15939 46948 -15892 47012
rect -15828 46948 -15812 47012
rect -15939 46932 -15812 46948
rect -15939 46868 -15892 46932
rect -15828 46868 -15812 46932
rect -15939 46852 -15812 46868
rect -15939 46788 -15892 46852
rect -15828 46788 -15812 46852
rect -15939 46772 -15812 46788
rect -15939 46708 -15892 46772
rect -15828 46708 -15812 46772
rect -15939 46692 -15812 46708
rect -15939 46628 -15892 46692
rect -15828 46628 -15812 46692
rect -15939 46612 -15812 46628
rect -15939 46548 -15892 46612
rect -15828 46548 -15812 46612
rect -15939 46532 -15812 46548
rect -15939 46468 -15892 46532
rect -15828 46468 -15812 46532
rect -15939 46452 -15812 46468
rect -15939 46388 -15892 46452
rect -15828 46388 -15812 46452
rect -15939 46372 -15812 46388
rect -15939 46308 -15892 46372
rect -15828 46308 -15812 46372
rect -15939 46292 -15812 46308
rect -15939 46228 -15892 46292
rect -15828 46228 -15812 46292
rect -15939 46212 -15812 46228
rect -15939 46148 -15892 46212
rect -15828 46148 -15812 46212
rect -15939 46132 -15812 46148
rect -15939 46068 -15892 46132
rect -15828 46068 -15812 46132
rect -15939 46052 -15812 46068
rect -15939 45988 -15892 46052
rect -15828 45988 -15812 46052
rect -15939 45972 -15812 45988
rect -15939 45908 -15892 45972
rect -15828 45908 -15812 45972
rect -15939 45892 -15812 45908
rect -15939 45828 -15892 45892
rect -15828 45828 -15812 45892
rect -15939 45812 -15812 45828
rect -15939 45748 -15892 45812
rect -15828 45748 -15812 45812
rect -15939 45732 -15812 45748
rect -15939 45668 -15892 45732
rect -15828 45668 -15812 45732
rect -15939 45652 -15812 45668
rect -15939 45588 -15892 45652
rect -15828 45588 -15812 45652
rect -15939 45572 -15812 45588
rect -15939 45508 -15892 45572
rect -15828 45508 -15812 45572
rect -15939 45492 -15812 45508
rect -15939 45428 -15892 45492
rect -15828 45428 -15812 45492
rect -15939 45412 -15812 45428
rect -15939 45348 -15892 45412
rect -15828 45348 -15812 45412
rect -15939 45332 -15812 45348
rect -15939 45268 -15892 45332
rect -15828 45268 -15812 45332
rect -15939 45252 -15812 45268
rect -15939 45188 -15892 45252
rect -15828 45188 -15812 45252
rect -15939 45172 -15812 45188
rect -15939 45108 -15892 45172
rect -15828 45108 -15812 45172
rect -15939 45092 -15812 45108
rect -15939 45028 -15892 45092
rect -15828 45028 -15812 45092
rect -15939 45012 -15812 45028
rect -15939 44948 -15892 45012
rect -15828 44948 -15812 45012
rect -15939 44932 -15812 44948
rect -15939 44868 -15892 44932
rect -15828 44868 -15812 44932
rect -15939 44852 -15812 44868
rect -15939 44788 -15892 44852
rect -15828 44788 -15812 44852
rect -15939 44772 -15812 44788
rect -15939 44708 -15892 44772
rect -15828 44708 -15812 44772
rect -15939 44692 -15812 44708
rect -15939 44628 -15892 44692
rect -15828 44628 -15812 44692
rect -15939 44612 -15812 44628
rect -15939 44548 -15892 44612
rect -15828 44548 -15812 44612
rect -15939 44532 -15812 44548
rect -15939 44468 -15892 44532
rect -15828 44468 -15812 44532
rect -15939 44452 -15812 44468
rect -15939 44388 -15892 44452
rect -15828 44388 -15812 44452
rect -15939 44372 -15812 44388
rect -15939 44308 -15892 44372
rect -15828 44308 -15812 44372
rect -15939 44292 -15812 44308
rect -15939 44228 -15892 44292
rect -15828 44228 -15812 44292
rect -15939 44212 -15812 44228
rect -15939 44148 -15892 44212
rect -15828 44148 -15812 44212
rect -15939 44132 -15812 44148
rect -15939 44068 -15892 44132
rect -15828 44068 -15812 44132
rect -15939 44052 -15812 44068
rect -15939 43988 -15892 44052
rect -15828 43988 -15812 44052
rect -15939 43972 -15812 43988
rect -15939 43908 -15892 43972
rect -15828 43908 -15812 43972
rect -15939 43892 -15812 43908
rect -15939 43828 -15892 43892
rect -15828 43828 -15812 43892
rect -15939 43812 -15812 43828
rect -15939 43748 -15892 43812
rect -15828 43748 -15812 43812
rect -15939 43732 -15812 43748
rect -15939 43668 -15892 43732
rect -15828 43668 -15812 43732
rect -15939 43652 -15812 43668
rect -15939 43588 -15892 43652
rect -15828 43588 -15812 43652
rect -15939 43572 -15812 43588
rect -15939 43508 -15892 43572
rect -15828 43508 -15812 43572
rect -15939 43492 -15812 43508
rect -15939 43428 -15892 43492
rect -15828 43428 -15812 43492
rect -15939 43412 -15812 43428
rect -15939 43348 -15892 43412
rect -15828 43348 -15812 43412
rect -15939 43332 -15812 43348
rect -15939 43268 -15892 43332
rect -15828 43268 -15812 43332
rect -15939 43252 -15812 43268
rect -15939 43188 -15892 43252
rect -15828 43188 -15812 43252
rect -15939 43172 -15812 43188
rect -15939 43108 -15892 43172
rect -15828 43108 -15812 43172
rect -15939 43092 -15812 43108
rect -15939 43028 -15892 43092
rect -15828 43028 -15812 43092
rect -15939 43012 -15812 43028
rect -15939 42948 -15892 43012
rect -15828 42948 -15812 43012
rect -15939 42932 -15812 42948
rect -15939 42868 -15892 42932
rect -15828 42868 -15812 42932
rect -15939 42852 -15812 42868
rect -15939 42788 -15892 42852
rect -15828 42788 -15812 42852
rect -15939 42772 -15812 42788
rect -15939 42708 -15892 42772
rect -15828 42708 -15812 42772
rect -15939 42692 -15812 42708
rect -15939 42628 -15892 42692
rect -15828 42628 -15812 42692
rect -15939 42612 -15812 42628
rect -15939 42548 -15892 42612
rect -15828 42548 -15812 42612
rect -15939 42532 -15812 42548
rect -15939 42468 -15892 42532
rect -15828 42468 -15812 42532
rect -15939 42452 -15812 42468
rect -15939 42388 -15892 42452
rect -15828 42388 -15812 42452
rect -15939 42372 -15812 42388
rect -15939 42308 -15892 42372
rect -15828 42308 -15812 42372
rect -15939 42292 -15812 42308
rect -15939 42228 -15892 42292
rect -15828 42228 -15812 42292
rect -15939 42212 -15812 42228
rect -15939 42148 -15892 42212
rect -15828 42148 -15812 42212
rect -15939 42132 -15812 42148
rect -15939 42068 -15892 42132
rect -15828 42068 -15812 42132
rect -15939 42052 -15812 42068
rect -15939 41988 -15892 42052
rect -15828 41988 -15812 42052
rect -15939 41972 -15812 41988
rect -15939 41908 -15892 41972
rect -15828 41908 -15812 41972
rect -15939 41892 -15812 41908
rect -15939 41828 -15892 41892
rect -15828 41828 -15812 41892
rect -15939 41812 -15812 41828
rect -15939 41748 -15892 41812
rect -15828 41748 -15812 41812
rect -15939 41732 -15812 41748
rect -15939 41668 -15892 41732
rect -15828 41668 -15812 41732
rect -15939 41652 -15812 41668
rect -15939 41588 -15892 41652
rect -15828 41588 -15812 41652
rect -15939 41572 -15812 41588
rect -15939 41508 -15892 41572
rect -15828 41508 -15812 41572
rect -15939 41492 -15812 41508
rect -15939 41428 -15892 41492
rect -15828 41428 -15812 41492
rect -15939 41412 -15812 41428
rect -15939 41348 -15892 41412
rect -15828 41348 -15812 41412
rect -15939 41332 -15812 41348
rect -15939 41268 -15892 41332
rect -15828 41268 -15812 41332
rect -15939 41252 -15812 41268
rect -15939 41188 -15892 41252
rect -15828 41188 -15812 41252
rect -15939 41172 -15812 41188
rect -22258 41092 -22131 41108
rect -22258 41028 -22211 41092
rect -22147 41028 -22131 41092
rect -22258 41012 -22131 41028
rect -22258 40888 -22154 41012
rect -22258 40872 -22131 40888
rect -22258 40808 -22211 40872
rect -22147 40808 -22131 40872
rect -22258 40792 -22131 40808
rect -28577 40712 -28450 40728
rect -28577 40648 -28530 40712
rect -28466 40648 -28450 40712
rect -28577 40632 -28450 40648
rect -28577 40568 -28530 40632
rect -28466 40568 -28450 40632
rect -28577 40552 -28450 40568
rect -28577 40488 -28530 40552
rect -28466 40488 -28450 40552
rect -28577 40472 -28450 40488
rect -28577 40408 -28530 40472
rect -28466 40408 -28450 40472
rect -28577 40392 -28450 40408
rect -28577 40328 -28530 40392
rect -28466 40328 -28450 40392
rect -28577 40312 -28450 40328
rect -28577 40248 -28530 40312
rect -28466 40248 -28450 40312
rect -28577 40232 -28450 40248
rect -28577 40168 -28530 40232
rect -28466 40168 -28450 40232
rect -28577 40152 -28450 40168
rect -28577 40088 -28530 40152
rect -28466 40088 -28450 40152
rect -28577 40072 -28450 40088
rect -28577 40008 -28530 40072
rect -28466 40008 -28450 40072
rect -28577 39992 -28450 40008
rect -28577 39928 -28530 39992
rect -28466 39928 -28450 39992
rect -28577 39912 -28450 39928
rect -28577 39848 -28530 39912
rect -28466 39848 -28450 39912
rect -28577 39832 -28450 39848
rect -28577 39768 -28530 39832
rect -28466 39768 -28450 39832
rect -28577 39752 -28450 39768
rect -28577 39688 -28530 39752
rect -28466 39688 -28450 39752
rect -28577 39672 -28450 39688
rect -28577 39608 -28530 39672
rect -28466 39608 -28450 39672
rect -28577 39592 -28450 39608
rect -28577 39528 -28530 39592
rect -28466 39528 -28450 39592
rect -28577 39512 -28450 39528
rect -28577 39448 -28530 39512
rect -28466 39448 -28450 39512
rect -28577 39432 -28450 39448
rect -28577 39368 -28530 39432
rect -28466 39368 -28450 39432
rect -28577 39352 -28450 39368
rect -28577 39288 -28530 39352
rect -28466 39288 -28450 39352
rect -28577 39272 -28450 39288
rect -28577 39208 -28530 39272
rect -28466 39208 -28450 39272
rect -28577 39192 -28450 39208
rect -28577 39128 -28530 39192
rect -28466 39128 -28450 39192
rect -28577 39112 -28450 39128
rect -28577 39048 -28530 39112
rect -28466 39048 -28450 39112
rect -28577 39032 -28450 39048
rect -28577 38968 -28530 39032
rect -28466 38968 -28450 39032
rect -28577 38952 -28450 38968
rect -28577 38888 -28530 38952
rect -28466 38888 -28450 38952
rect -28577 38872 -28450 38888
rect -28577 38808 -28530 38872
rect -28466 38808 -28450 38872
rect -28577 38792 -28450 38808
rect -28577 38728 -28530 38792
rect -28466 38728 -28450 38792
rect -28577 38712 -28450 38728
rect -28577 38648 -28530 38712
rect -28466 38648 -28450 38712
rect -28577 38632 -28450 38648
rect -28577 38568 -28530 38632
rect -28466 38568 -28450 38632
rect -28577 38552 -28450 38568
rect -28577 38488 -28530 38552
rect -28466 38488 -28450 38552
rect -28577 38472 -28450 38488
rect -28577 38408 -28530 38472
rect -28466 38408 -28450 38472
rect -28577 38392 -28450 38408
rect -28577 38328 -28530 38392
rect -28466 38328 -28450 38392
rect -28577 38312 -28450 38328
rect -28577 38248 -28530 38312
rect -28466 38248 -28450 38312
rect -28577 38232 -28450 38248
rect -28577 38168 -28530 38232
rect -28466 38168 -28450 38232
rect -28577 38152 -28450 38168
rect -28577 38088 -28530 38152
rect -28466 38088 -28450 38152
rect -28577 38072 -28450 38088
rect -28577 38008 -28530 38072
rect -28466 38008 -28450 38072
rect -28577 37992 -28450 38008
rect -28577 37928 -28530 37992
rect -28466 37928 -28450 37992
rect -28577 37912 -28450 37928
rect -28577 37848 -28530 37912
rect -28466 37848 -28450 37912
rect -28577 37832 -28450 37848
rect -28577 37768 -28530 37832
rect -28466 37768 -28450 37832
rect -28577 37752 -28450 37768
rect -28577 37688 -28530 37752
rect -28466 37688 -28450 37752
rect -28577 37672 -28450 37688
rect -28577 37608 -28530 37672
rect -28466 37608 -28450 37672
rect -28577 37592 -28450 37608
rect -28577 37528 -28530 37592
rect -28466 37528 -28450 37592
rect -28577 37512 -28450 37528
rect -28577 37448 -28530 37512
rect -28466 37448 -28450 37512
rect -28577 37432 -28450 37448
rect -28577 37368 -28530 37432
rect -28466 37368 -28450 37432
rect -28577 37352 -28450 37368
rect -28577 37288 -28530 37352
rect -28466 37288 -28450 37352
rect -28577 37272 -28450 37288
rect -28577 37208 -28530 37272
rect -28466 37208 -28450 37272
rect -28577 37192 -28450 37208
rect -28577 37128 -28530 37192
rect -28466 37128 -28450 37192
rect -28577 37112 -28450 37128
rect -28577 37048 -28530 37112
rect -28466 37048 -28450 37112
rect -28577 37032 -28450 37048
rect -28577 36968 -28530 37032
rect -28466 36968 -28450 37032
rect -28577 36952 -28450 36968
rect -28577 36888 -28530 36952
rect -28466 36888 -28450 36952
rect -28577 36872 -28450 36888
rect -28577 36808 -28530 36872
rect -28466 36808 -28450 36872
rect -28577 36792 -28450 36808
rect -28577 36728 -28530 36792
rect -28466 36728 -28450 36792
rect -28577 36712 -28450 36728
rect -28577 36648 -28530 36712
rect -28466 36648 -28450 36712
rect -28577 36632 -28450 36648
rect -28577 36568 -28530 36632
rect -28466 36568 -28450 36632
rect -28577 36552 -28450 36568
rect -28577 36488 -28530 36552
rect -28466 36488 -28450 36552
rect -28577 36472 -28450 36488
rect -28577 36408 -28530 36472
rect -28466 36408 -28450 36472
rect -28577 36392 -28450 36408
rect -28577 36328 -28530 36392
rect -28466 36328 -28450 36392
rect -28577 36312 -28450 36328
rect -28577 36248 -28530 36312
rect -28466 36248 -28450 36312
rect -28577 36232 -28450 36248
rect -28577 36168 -28530 36232
rect -28466 36168 -28450 36232
rect -28577 36152 -28450 36168
rect -28577 36088 -28530 36152
rect -28466 36088 -28450 36152
rect -28577 36072 -28450 36088
rect -28577 36008 -28530 36072
rect -28466 36008 -28450 36072
rect -28577 35992 -28450 36008
rect -28577 35928 -28530 35992
rect -28466 35928 -28450 35992
rect -28577 35912 -28450 35928
rect -28577 35848 -28530 35912
rect -28466 35848 -28450 35912
rect -28577 35832 -28450 35848
rect -28577 35768 -28530 35832
rect -28466 35768 -28450 35832
rect -28577 35752 -28450 35768
rect -28577 35688 -28530 35752
rect -28466 35688 -28450 35752
rect -28577 35672 -28450 35688
rect -28577 35608 -28530 35672
rect -28466 35608 -28450 35672
rect -28577 35592 -28450 35608
rect -28577 35528 -28530 35592
rect -28466 35528 -28450 35592
rect -28577 35512 -28450 35528
rect -28577 35448 -28530 35512
rect -28466 35448 -28450 35512
rect -28577 35432 -28450 35448
rect -28577 35368 -28530 35432
rect -28466 35368 -28450 35432
rect -28577 35352 -28450 35368
rect -28577 35288 -28530 35352
rect -28466 35288 -28450 35352
rect -28577 35272 -28450 35288
rect -28577 35208 -28530 35272
rect -28466 35208 -28450 35272
rect -28577 35192 -28450 35208
rect -28577 35128 -28530 35192
rect -28466 35128 -28450 35192
rect -28577 35112 -28450 35128
rect -28577 35048 -28530 35112
rect -28466 35048 -28450 35112
rect -28577 35032 -28450 35048
rect -28577 34968 -28530 35032
rect -28466 34968 -28450 35032
rect -28577 34952 -28450 34968
rect -28577 34888 -28530 34952
rect -28466 34888 -28450 34952
rect -28577 34872 -28450 34888
rect -34896 34792 -34769 34808
rect -34896 34728 -34849 34792
rect -34785 34728 -34769 34792
rect -34896 34712 -34769 34728
rect -34896 34588 -34792 34712
rect -34896 34572 -34769 34588
rect -34896 34508 -34849 34572
rect -34785 34508 -34769 34572
rect -34896 34492 -34769 34508
rect -41215 34412 -41088 34428
rect -41215 34348 -41168 34412
rect -41104 34348 -41088 34412
rect -41215 34332 -41088 34348
rect -41215 34268 -41168 34332
rect -41104 34268 -41088 34332
rect -41215 34252 -41088 34268
rect -41215 34188 -41168 34252
rect -41104 34188 -41088 34252
rect -41215 34172 -41088 34188
rect -41215 34108 -41168 34172
rect -41104 34108 -41088 34172
rect -41215 34092 -41088 34108
rect -41215 34028 -41168 34092
rect -41104 34028 -41088 34092
rect -41215 34012 -41088 34028
rect -41215 33948 -41168 34012
rect -41104 33948 -41088 34012
rect -41215 33932 -41088 33948
rect -41215 33868 -41168 33932
rect -41104 33868 -41088 33932
rect -41215 33852 -41088 33868
rect -41215 33788 -41168 33852
rect -41104 33788 -41088 33852
rect -41215 33772 -41088 33788
rect -41215 33708 -41168 33772
rect -41104 33708 -41088 33772
rect -41215 33692 -41088 33708
rect -41215 33628 -41168 33692
rect -41104 33628 -41088 33692
rect -41215 33612 -41088 33628
rect -41215 33548 -41168 33612
rect -41104 33548 -41088 33612
rect -41215 33532 -41088 33548
rect -41215 33468 -41168 33532
rect -41104 33468 -41088 33532
rect -41215 33452 -41088 33468
rect -41215 33388 -41168 33452
rect -41104 33388 -41088 33452
rect -41215 33372 -41088 33388
rect -41215 33308 -41168 33372
rect -41104 33308 -41088 33372
rect -41215 33292 -41088 33308
rect -41215 33228 -41168 33292
rect -41104 33228 -41088 33292
rect -41215 33212 -41088 33228
rect -41215 33148 -41168 33212
rect -41104 33148 -41088 33212
rect -41215 33132 -41088 33148
rect -41215 33068 -41168 33132
rect -41104 33068 -41088 33132
rect -41215 33052 -41088 33068
rect -41215 32988 -41168 33052
rect -41104 32988 -41088 33052
rect -41215 32972 -41088 32988
rect -41215 32908 -41168 32972
rect -41104 32908 -41088 32972
rect -41215 32892 -41088 32908
rect -41215 32828 -41168 32892
rect -41104 32828 -41088 32892
rect -41215 32812 -41088 32828
rect -41215 32748 -41168 32812
rect -41104 32748 -41088 32812
rect -41215 32732 -41088 32748
rect -41215 32668 -41168 32732
rect -41104 32668 -41088 32732
rect -41215 32652 -41088 32668
rect -41215 32588 -41168 32652
rect -41104 32588 -41088 32652
rect -41215 32572 -41088 32588
rect -41215 32508 -41168 32572
rect -41104 32508 -41088 32572
rect -41215 32492 -41088 32508
rect -41215 32428 -41168 32492
rect -41104 32428 -41088 32492
rect -41215 32412 -41088 32428
rect -41215 32348 -41168 32412
rect -41104 32348 -41088 32412
rect -41215 32332 -41088 32348
rect -41215 32268 -41168 32332
rect -41104 32268 -41088 32332
rect -41215 32252 -41088 32268
rect -41215 32188 -41168 32252
rect -41104 32188 -41088 32252
rect -41215 32172 -41088 32188
rect -41215 32108 -41168 32172
rect -41104 32108 -41088 32172
rect -41215 32092 -41088 32108
rect -41215 32028 -41168 32092
rect -41104 32028 -41088 32092
rect -41215 32012 -41088 32028
rect -41215 31948 -41168 32012
rect -41104 31948 -41088 32012
rect -41215 31932 -41088 31948
rect -41215 31868 -41168 31932
rect -41104 31868 -41088 31932
rect -41215 31852 -41088 31868
rect -41215 31788 -41168 31852
rect -41104 31788 -41088 31852
rect -41215 31772 -41088 31788
rect -41215 31708 -41168 31772
rect -41104 31708 -41088 31772
rect -41215 31692 -41088 31708
rect -41215 31628 -41168 31692
rect -41104 31628 -41088 31692
rect -41215 31612 -41088 31628
rect -41215 31548 -41168 31612
rect -41104 31548 -41088 31612
rect -41215 31532 -41088 31548
rect -41215 31468 -41168 31532
rect -41104 31468 -41088 31532
rect -41215 31452 -41088 31468
rect -41215 31388 -41168 31452
rect -41104 31388 -41088 31452
rect -41215 31372 -41088 31388
rect -41215 31308 -41168 31372
rect -41104 31308 -41088 31372
rect -41215 31292 -41088 31308
rect -41215 31228 -41168 31292
rect -41104 31228 -41088 31292
rect -41215 31212 -41088 31228
rect -41215 31148 -41168 31212
rect -41104 31148 -41088 31212
rect -41215 31132 -41088 31148
rect -41215 31068 -41168 31132
rect -41104 31068 -41088 31132
rect -41215 31052 -41088 31068
rect -41215 30988 -41168 31052
rect -41104 30988 -41088 31052
rect -41215 30972 -41088 30988
rect -41215 30908 -41168 30972
rect -41104 30908 -41088 30972
rect -41215 30892 -41088 30908
rect -41215 30828 -41168 30892
rect -41104 30828 -41088 30892
rect -41215 30812 -41088 30828
rect -41215 30748 -41168 30812
rect -41104 30748 -41088 30812
rect -41215 30732 -41088 30748
rect -41215 30668 -41168 30732
rect -41104 30668 -41088 30732
rect -41215 30652 -41088 30668
rect -41215 30588 -41168 30652
rect -41104 30588 -41088 30652
rect -41215 30572 -41088 30588
rect -41215 30508 -41168 30572
rect -41104 30508 -41088 30572
rect -41215 30492 -41088 30508
rect -41215 30428 -41168 30492
rect -41104 30428 -41088 30492
rect -41215 30412 -41088 30428
rect -41215 30348 -41168 30412
rect -41104 30348 -41088 30412
rect -41215 30332 -41088 30348
rect -41215 30268 -41168 30332
rect -41104 30268 -41088 30332
rect -41215 30252 -41088 30268
rect -41215 30188 -41168 30252
rect -41104 30188 -41088 30252
rect -41215 30172 -41088 30188
rect -41215 30108 -41168 30172
rect -41104 30108 -41088 30172
rect -41215 30092 -41088 30108
rect -41215 30028 -41168 30092
rect -41104 30028 -41088 30092
rect -41215 30012 -41088 30028
rect -41215 29948 -41168 30012
rect -41104 29948 -41088 30012
rect -41215 29932 -41088 29948
rect -41215 29868 -41168 29932
rect -41104 29868 -41088 29932
rect -41215 29852 -41088 29868
rect -41215 29788 -41168 29852
rect -41104 29788 -41088 29852
rect -41215 29772 -41088 29788
rect -41215 29708 -41168 29772
rect -41104 29708 -41088 29772
rect -41215 29692 -41088 29708
rect -41215 29628 -41168 29692
rect -41104 29628 -41088 29692
rect -41215 29612 -41088 29628
rect -41215 29548 -41168 29612
rect -41104 29548 -41088 29612
rect -41215 29532 -41088 29548
rect -41215 29468 -41168 29532
rect -41104 29468 -41088 29532
rect -41215 29452 -41088 29468
rect -41215 29388 -41168 29452
rect -41104 29388 -41088 29452
rect -41215 29372 -41088 29388
rect -41215 29308 -41168 29372
rect -41104 29308 -41088 29372
rect -41215 29292 -41088 29308
rect -41215 29228 -41168 29292
rect -41104 29228 -41088 29292
rect -41215 29212 -41088 29228
rect -41215 29148 -41168 29212
rect -41104 29148 -41088 29212
rect -41215 29132 -41088 29148
rect -41215 29068 -41168 29132
rect -41104 29068 -41088 29132
rect -41215 29052 -41088 29068
rect -41215 28988 -41168 29052
rect -41104 28988 -41088 29052
rect -41215 28972 -41088 28988
rect -41215 28908 -41168 28972
rect -41104 28908 -41088 28972
rect -41215 28892 -41088 28908
rect -41215 28828 -41168 28892
rect -41104 28828 -41088 28892
rect -41215 28812 -41088 28828
rect -41215 28748 -41168 28812
rect -41104 28748 -41088 28812
rect -41215 28732 -41088 28748
rect -41215 28668 -41168 28732
rect -41104 28668 -41088 28732
rect -41215 28652 -41088 28668
rect -41215 28588 -41168 28652
rect -41104 28588 -41088 28652
rect -41215 28572 -41088 28588
rect -44335 28161 -44231 28539
rect -41215 28508 -41168 28572
rect -41104 28508 -41088 28572
rect -40925 34452 -35003 34461
rect -40925 28548 -40916 34452
rect -35012 28548 -35003 34452
rect -40925 28539 -35003 28548
rect -34896 34428 -34849 34492
rect -34785 34428 -34769 34492
rect -31697 34461 -31593 34839
rect -28577 34808 -28530 34872
rect -28466 34808 -28450 34872
rect -28287 40752 -22365 40761
rect -28287 34848 -28278 40752
rect -22374 34848 -22365 40752
rect -28287 34839 -22365 34848
rect -22258 40728 -22211 40792
rect -22147 40728 -22131 40792
rect -19059 40761 -18955 41139
rect -15939 41108 -15892 41172
rect -15828 41108 -15812 41172
rect -15649 47052 -9727 47061
rect -15649 41148 -15640 47052
rect -9736 41148 -9727 47052
rect -15649 41139 -9727 41148
rect -9620 47028 -9573 47092
rect -9509 47028 -9493 47092
rect -6421 47061 -6317 47250
rect -3301 47188 -3197 47250
rect -3301 47172 -3174 47188
rect -3301 47108 -3254 47172
rect -3190 47108 -3174 47172
rect -3301 47092 -3174 47108
rect -9620 47012 -9493 47028
rect -9620 46948 -9573 47012
rect -9509 46948 -9493 47012
rect -9620 46932 -9493 46948
rect -9620 46868 -9573 46932
rect -9509 46868 -9493 46932
rect -9620 46852 -9493 46868
rect -9620 46788 -9573 46852
rect -9509 46788 -9493 46852
rect -9620 46772 -9493 46788
rect -9620 46708 -9573 46772
rect -9509 46708 -9493 46772
rect -9620 46692 -9493 46708
rect -9620 46628 -9573 46692
rect -9509 46628 -9493 46692
rect -9620 46612 -9493 46628
rect -9620 46548 -9573 46612
rect -9509 46548 -9493 46612
rect -9620 46532 -9493 46548
rect -9620 46468 -9573 46532
rect -9509 46468 -9493 46532
rect -9620 46452 -9493 46468
rect -9620 46388 -9573 46452
rect -9509 46388 -9493 46452
rect -9620 46372 -9493 46388
rect -9620 46308 -9573 46372
rect -9509 46308 -9493 46372
rect -9620 46292 -9493 46308
rect -9620 46228 -9573 46292
rect -9509 46228 -9493 46292
rect -9620 46212 -9493 46228
rect -9620 46148 -9573 46212
rect -9509 46148 -9493 46212
rect -9620 46132 -9493 46148
rect -9620 46068 -9573 46132
rect -9509 46068 -9493 46132
rect -9620 46052 -9493 46068
rect -9620 45988 -9573 46052
rect -9509 45988 -9493 46052
rect -9620 45972 -9493 45988
rect -9620 45908 -9573 45972
rect -9509 45908 -9493 45972
rect -9620 45892 -9493 45908
rect -9620 45828 -9573 45892
rect -9509 45828 -9493 45892
rect -9620 45812 -9493 45828
rect -9620 45748 -9573 45812
rect -9509 45748 -9493 45812
rect -9620 45732 -9493 45748
rect -9620 45668 -9573 45732
rect -9509 45668 -9493 45732
rect -9620 45652 -9493 45668
rect -9620 45588 -9573 45652
rect -9509 45588 -9493 45652
rect -9620 45572 -9493 45588
rect -9620 45508 -9573 45572
rect -9509 45508 -9493 45572
rect -9620 45492 -9493 45508
rect -9620 45428 -9573 45492
rect -9509 45428 -9493 45492
rect -9620 45412 -9493 45428
rect -9620 45348 -9573 45412
rect -9509 45348 -9493 45412
rect -9620 45332 -9493 45348
rect -9620 45268 -9573 45332
rect -9509 45268 -9493 45332
rect -9620 45252 -9493 45268
rect -9620 45188 -9573 45252
rect -9509 45188 -9493 45252
rect -9620 45172 -9493 45188
rect -9620 45108 -9573 45172
rect -9509 45108 -9493 45172
rect -9620 45092 -9493 45108
rect -9620 45028 -9573 45092
rect -9509 45028 -9493 45092
rect -9620 45012 -9493 45028
rect -9620 44948 -9573 45012
rect -9509 44948 -9493 45012
rect -9620 44932 -9493 44948
rect -9620 44868 -9573 44932
rect -9509 44868 -9493 44932
rect -9620 44852 -9493 44868
rect -9620 44788 -9573 44852
rect -9509 44788 -9493 44852
rect -9620 44772 -9493 44788
rect -9620 44708 -9573 44772
rect -9509 44708 -9493 44772
rect -9620 44692 -9493 44708
rect -9620 44628 -9573 44692
rect -9509 44628 -9493 44692
rect -9620 44612 -9493 44628
rect -9620 44548 -9573 44612
rect -9509 44548 -9493 44612
rect -9620 44532 -9493 44548
rect -9620 44468 -9573 44532
rect -9509 44468 -9493 44532
rect -9620 44452 -9493 44468
rect -9620 44388 -9573 44452
rect -9509 44388 -9493 44452
rect -9620 44372 -9493 44388
rect -9620 44308 -9573 44372
rect -9509 44308 -9493 44372
rect -9620 44292 -9493 44308
rect -9620 44228 -9573 44292
rect -9509 44228 -9493 44292
rect -9620 44212 -9493 44228
rect -9620 44148 -9573 44212
rect -9509 44148 -9493 44212
rect -9620 44132 -9493 44148
rect -9620 44068 -9573 44132
rect -9509 44068 -9493 44132
rect -9620 44052 -9493 44068
rect -9620 43988 -9573 44052
rect -9509 43988 -9493 44052
rect -9620 43972 -9493 43988
rect -9620 43908 -9573 43972
rect -9509 43908 -9493 43972
rect -9620 43892 -9493 43908
rect -9620 43828 -9573 43892
rect -9509 43828 -9493 43892
rect -9620 43812 -9493 43828
rect -9620 43748 -9573 43812
rect -9509 43748 -9493 43812
rect -9620 43732 -9493 43748
rect -9620 43668 -9573 43732
rect -9509 43668 -9493 43732
rect -9620 43652 -9493 43668
rect -9620 43588 -9573 43652
rect -9509 43588 -9493 43652
rect -9620 43572 -9493 43588
rect -9620 43508 -9573 43572
rect -9509 43508 -9493 43572
rect -9620 43492 -9493 43508
rect -9620 43428 -9573 43492
rect -9509 43428 -9493 43492
rect -9620 43412 -9493 43428
rect -9620 43348 -9573 43412
rect -9509 43348 -9493 43412
rect -9620 43332 -9493 43348
rect -9620 43268 -9573 43332
rect -9509 43268 -9493 43332
rect -9620 43252 -9493 43268
rect -9620 43188 -9573 43252
rect -9509 43188 -9493 43252
rect -9620 43172 -9493 43188
rect -9620 43108 -9573 43172
rect -9509 43108 -9493 43172
rect -9620 43092 -9493 43108
rect -9620 43028 -9573 43092
rect -9509 43028 -9493 43092
rect -9620 43012 -9493 43028
rect -9620 42948 -9573 43012
rect -9509 42948 -9493 43012
rect -9620 42932 -9493 42948
rect -9620 42868 -9573 42932
rect -9509 42868 -9493 42932
rect -9620 42852 -9493 42868
rect -9620 42788 -9573 42852
rect -9509 42788 -9493 42852
rect -9620 42772 -9493 42788
rect -9620 42708 -9573 42772
rect -9509 42708 -9493 42772
rect -9620 42692 -9493 42708
rect -9620 42628 -9573 42692
rect -9509 42628 -9493 42692
rect -9620 42612 -9493 42628
rect -9620 42548 -9573 42612
rect -9509 42548 -9493 42612
rect -9620 42532 -9493 42548
rect -9620 42468 -9573 42532
rect -9509 42468 -9493 42532
rect -9620 42452 -9493 42468
rect -9620 42388 -9573 42452
rect -9509 42388 -9493 42452
rect -9620 42372 -9493 42388
rect -9620 42308 -9573 42372
rect -9509 42308 -9493 42372
rect -9620 42292 -9493 42308
rect -9620 42228 -9573 42292
rect -9509 42228 -9493 42292
rect -9620 42212 -9493 42228
rect -9620 42148 -9573 42212
rect -9509 42148 -9493 42212
rect -9620 42132 -9493 42148
rect -9620 42068 -9573 42132
rect -9509 42068 -9493 42132
rect -9620 42052 -9493 42068
rect -9620 41988 -9573 42052
rect -9509 41988 -9493 42052
rect -9620 41972 -9493 41988
rect -9620 41908 -9573 41972
rect -9509 41908 -9493 41972
rect -9620 41892 -9493 41908
rect -9620 41828 -9573 41892
rect -9509 41828 -9493 41892
rect -9620 41812 -9493 41828
rect -9620 41748 -9573 41812
rect -9509 41748 -9493 41812
rect -9620 41732 -9493 41748
rect -9620 41668 -9573 41732
rect -9509 41668 -9493 41732
rect -9620 41652 -9493 41668
rect -9620 41588 -9573 41652
rect -9509 41588 -9493 41652
rect -9620 41572 -9493 41588
rect -9620 41508 -9573 41572
rect -9509 41508 -9493 41572
rect -9620 41492 -9493 41508
rect -9620 41428 -9573 41492
rect -9509 41428 -9493 41492
rect -9620 41412 -9493 41428
rect -9620 41348 -9573 41412
rect -9509 41348 -9493 41412
rect -9620 41332 -9493 41348
rect -9620 41268 -9573 41332
rect -9509 41268 -9493 41332
rect -9620 41252 -9493 41268
rect -9620 41188 -9573 41252
rect -9509 41188 -9493 41252
rect -9620 41172 -9493 41188
rect -15939 41092 -15812 41108
rect -15939 41028 -15892 41092
rect -15828 41028 -15812 41092
rect -15939 41012 -15812 41028
rect -15939 40888 -15835 41012
rect -15939 40872 -15812 40888
rect -15939 40808 -15892 40872
rect -15828 40808 -15812 40872
rect -15939 40792 -15812 40808
rect -22258 40712 -22131 40728
rect -22258 40648 -22211 40712
rect -22147 40648 -22131 40712
rect -22258 40632 -22131 40648
rect -22258 40568 -22211 40632
rect -22147 40568 -22131 40632
rect -22258 40552 -22131 40568
rect -22258 40488 -22211 40552
rect -22147 40488 -22131 40552
rect -22258 40472 -22131 40488
rect -22258 40408 -22211 40472
rect -22147 40408 -22131 40472
rect -22258 40392 -22131 40408
rect -22258 40328 -22211 40392
rect -22147 40328 -22131 40392
rect -22258 40312 -22131 40328
rect -22258 40248 -22211 40312
rect -22147 40248 -22131 40312
rect -22258 40232 -22131 40248
rect -22258 40168 -22211 40232
rect -22147 40168 -22131 40232
rect -22258 40152 -22131 40168
rect -22258 40088 -22211 40152
rect -22147 40088 -22131 40152
rect -22258 40072 -22131 40088
rect -22258 40008 -22211 40072
rect -22147 40008 -22131 40072
rect -22258 39992 -22131 40008
rect -22258 39928 -22211 39992
rect -22147 39928 -22131 39992
rect -22258 39912 -22131 39928
rect -22258 39848 -22211 39912
rect -22147 39848 -22131 39912
rect -22258 39832 -22131 39848
rect -22258 39768 -22211 39832
rect -22147 39768 -22131 39832
rect -22258 39752 -22131 39768
rect -22258 39688 -22211 39752
rect -22147 39688 -22131 39752
rect -22258 39672 -22131 39688
rect -22258 39608 -22211 39672
rect -22147 39608 -22131 39672
rect -22258 39592 -22131 39608
rect -22258 39528 -22211 39592
rect -22147 39528 -22131 39592
rect -22258 39512 -22131 39528
rect -22258 39448 -22211 39512
rect -22147 39448 -22131 39512
rect -22258 39432 -22131 39448
rect -22258 39368 -22211 39432
rect -22147 39368 -22131 39432
rect -22258 39352 -22131 39368
rect -22258 39288 -22211 39352
rect -22147 39288 -22131 39352
rect -22258 39272 -22131 39288
rect -22258 39208 -22211 39272
rect -22147 39208 -22131 39272
rect -22258 39192 -22131 39208
rect -22258 39128 -22211 39192
rect -22147 39128 -22131 39192
rect -22258 39112 -22131 39128
rect -22258 39048 -22211 39112
rect -22147 39048 -22131 39112
rect -22258 39032 -22131 39048
rect -22258 38968 -22211 39032
rect -22147 38968 -22131 39032
rect -22258 38952 -22131 38968
rect -22258 38888 -22211 38952
rect -22147 38888 -22131 38952
rect -22258 38872 -22131 38888
rect -22258 38808 -22211 38872
rect -22147 38808 -22131 38872
rect -22258 38792 -22131 38808
rect -22258 38728 -22211 38792
rect -22147 38728 -22131 38792
rect -22258 38712 -22131 38728
rect -22258 38648 -22211 38712
rect -22147 38648 -22131 38712
rect -22258 38632 -22131 38648
rect -22258 38568 -22211 38632
rect -22147 38568 -22131 38632
rect -22258 38552 -22131 38568
rect -22258 38488 -22211 38552
rect -22147 38488 -22131 38552
rect -22258 38472 -22131 38488
rect -22258 38408 -22211 38472
rect -22147 38408 -22131 38472
rect -22258 38392 -22131 38408
rect -22258 38328 -22211 38392
rect -22147 38328 -22131 38392
rect -22258 38312 -22131 38328
rect -22258 38248 -22211 38312
rect -22147 38248 -22131 38312
rect -22258 38232 -22131 38248
rect -22258 38168 -22211 38232
rect -22147 38168 -22131 38232
rect -22258 38152 -22131 38168
rect -22258 38088 -22211 38152
rect -22147 38088 -22131 38152
rect -22258 38072 -22131 38088
rect -22258 38008 -22211 38072
rect -22147 38008 -22131 38072
rect -22258 37992 -22131 38008
rect -22258 37928 -22211 37992
rect -22147 37928 -22131 37992
rect -22258 37912 -22131 37928
rect -22258 37848 -22211 37912
rect -22147 37848 -22131 37912
rect -22258 37832 -22131 37848
rect -22258 37768 -22211 37832
rect -22147 37768 -22131 37832
rect -22258 37752 -22131 37768
rect -22258 37688 -22211 37752
rect -22147 37688 -22131 37752
rect -22258 37672 -22131 37688
rect -22258 37608 -22211 37672
rect -22147 37608 -22131 37672
rect -22258 37592 -22131 37608
rect -22258 37528 -22211 37592
rect -22147 37528 -22131 37592
rect -22258 37512 -22131 37528
rect -22258 37448 -22211 37512
rect -22147 37448 -22131 37512
rect -22258 37432 -22131 37448
rect -22258 37368 -22211 37432
rect -22147 37368 -22131 37432
rect -22258 37352 -22131 37368
rect -22258 37288 -22211 37352
rect -22147 37288 -22131 37352
rect -22258 37272 -22131 37288
rect -22258 37208 -22211 37272
rect -22147 37208 -22131 37272
rect -22258 37192 -22131 37208
rect -22258 37128 -22211 37192
rect -22147 37128 -22131 37192
rect -22258 37112 -22131 37128
rect -22258 37048 -22211 37112
rect -22147 37048 -22131 37112
rect -22258 37032 -22131 37048
rect -22258 36968 -22211 37032
rect -22147 36968 -22131 37032
rect -22258 36952 -22131 36968
rect -22258 36888 -22211 36952
rect -22147 36888 -22131 36952
rect -22258 36872 -22131 36888
rect -22258 36808 -22211 36872
rect -22147 36808 -22131 36872
rect -22258 36792 -22131 36808
rect -22258 36728 -22211 36792
rect -22147 36728 -22131 36792
rect -22258 36712 -22131 36728
rect -22258 36648 -22211 36712
rect -22147 36648 -22131 36712
rect -22258 36632 -22131 36648
rect -22258 36568 -22211 36632
rect -22147 36568 -22131 36632
rect -22258 36552 -22131 36568
rect -22258 36488 -22211 36552
rect -22147 36488 -22131 36552
rect -22258 36472 -22131 36488
rect -22258 36408 -22211 36472
rect -22147 36408 -22131 36472
rect -22258 36392 -22131 36408
rect -22258 36328 -22211 36392
rect -22147 36328 -22131 36392
rect -22258 36312 -22131 36328
rect -22258 36248 -22211 36312
rect -22147 36248 -22131 36312
rect -22258 36232 -22131 36248
rect -22258 36168 -22211 36232
rect -22147 36168 -22131 36232
rect -22258 36152 -22131 36168
rect -22258 36088 -22211 36152
rect -22147 36088 -22131 36152
rect -22258 36072 -22131 36088
rect -22258 36008 -22211 36072
rect -22147 36008 -22131 36072
rect -22258 35992 -22131 36008
rect -22258 35928 -22211 35992
rect -22147 35928 -22131 35992
rect -22258 35912 -22131 35928
rect -22258 35848 -22211 35912
rect -22147 35848 -22131 35912
rect -22258 35832 -22131 35848
rect -22258 35768 -22211 35832
rect -22147 35768 -22131 35832
rect -22258 35752 -22131 35768
rect -22258 35688 -22211 35752
rect -22147 35688 -22131 35752
rect -22258 35672 -22131 35688
rect -22258 35608 -22211 35672
rect -22147 35608 -22131 35672
rect -22258 35592 -22131 35608
rect -22258 35528 -22211 35592
rect -22147 35528 -22131 35592
rect -22258 35512 -22131 35528
rect -22258 35448 -22211 35512
rect -22147 35448 -22131 35512
rect -22258 35432 -22131 35448
rect -22258 35368 -22211 35432
rect -22147 35368 -22131 35432
rect -22258 35352 -22131 35368
rect -22258 35288 -22211 35352
rect -22147 35288 -22131 35352
rect -22258 35272 -22131 35288
rect -22258 35208 -22211 35272
rect -22147 35208 -22131 35272
rect -22258 35192 -22131 35208
rect -22258 35128 -22211 35192
rect -22147 35128 -22131 35192
rect -22258 35112 -22131 35128
rect -22258 35048 -22211 35112
rect -22147 35048 -22131 35112
rect -22258 35032 -22131 35048
rect -22258 34968 -22211 35032
rect -22147 34968 -22131 35032
rect -22258 34952 -22131 34968
rect -22258 34888 -22211 34952
rect -22147 34888 -22131 34952
rect -22258 34872 -22131 34888
rect -28577 34792 -28450 34808
rect -28577 34728 -28530 34792
rect -28466 34728 -28450 34792
rect -28577 34712 -28450 34728
rect -28577 34588 -28473 34712
rect -28577 34572 -28450 34588
rect -28577 34508 -28530 34572
rect -28466 34508 -28450 34572
rect -28577 34492 -28450 34508
rect -34896 34412 -34769 34428
rect -34896 34348 -34849 34412
rect -34785 34348 -34769 34412
rect -34896 34332 -34769 34348
rect -34896 34268 -34849 34332
rect -34785 34268 -34769 34332
rect -34896 34252 -34769 34268
rect -34896 34188 -34849 34252
rect -34785 34188 -34769 34252
rect -34896 34172 -34769 34188
rect -34896 34108 -34849 34172
rect -34785 34108 -34769 34172
rect -34896 34092 -34769 34108
rect -34896 34028 -34849 34092
rect -34785 34028 -34769 34092
rect -34896 34012 -34769 34028
rect -34896 33948 -34849 34012
rect -34785 33948 -34769 34012
rect -34896 33932 -34769 33948
rect -34896 33868 -34849 33932
rect -34785 33868 -34769 33932
rect -34896 33852 -34769 33868
rect -34896 33788 -34849 33852
rect -34785 33788 -34769 33852
rect -34896 33772 -34769 33788
rect -34896 33708 -34849 33772
rect -34785 33708 -34769 33772
rect -34896 33692 -34769 33708
rect -34896 33628 -34849 33692
rect -34785 33628 -34769 33692
rect -34896 33612 -34769 33628
rect -34896 33548 -34849 33612
rect -34785 33548 -34769 33612
rect -34896 33532 -34769 33548
rect -34896 33468 -34849 33532
rect -34785 33468 -34769 33532
rect -34896 33452 -34769 33468
rect -34896 33388 -34849 33452
rect -34785 33388 -34769 33452
rect -34896 33372 -34769 33388
rect -34896 33308 -34849 33372
rect -34785 33308 -34769 33372
rect -34896 33292 -34769 33308
rect -34896 33228 -34849 33292
rect -34785 33228 -34769 33292
rect -34896 33212 -34769 33228
rect -34896 33148 -34849 33212
rect -34785 33148 -34769 33212
rect -34896 33132 -34769 33148
rect -34896 33068 -34849 33132
rect -34785 33068 -34769 33132
rect -34896 33052 -34769 33068
rect -34896 32988 -34849 33052
rect -34785 32988 -34769 33052
rect -34896 32972 -34769 32988
rect -34896 32908 -34849 32972
rect -34785 32908 -34769 32972
rect -34896 32892 -34769 32908
rect -34896 32828 -34849 32892
rect -34785 32828 -34769 32892
rect -34896 32812 -34769 32828
rect -34896 32748 -34849 32812
rect -34785 32748 -34769 32812
rect -34896 32732 -34769 32748
rect -34896 32668 -34849 32732
rect -34785 32668 -34769 32732
rect -34896 32652 -34769 32668
rect -34896 32588 -34849 32652
rect -34785 32588 -34769 32652
rect -34896 32572 -34769 32588
rect -34896 32508 -34849 32572
rect -34785 32508 -34769 32572
rect -34896 32492 -34769 32508
rect -34896 32428 -34849 32492
rect -34785 32428 -34769 32492
rect -34896 32412 -34769 32428
rect -34896 32348 -34849 32412
rect -34785 32348 -34769 32412
rect -34896 32332 -34769 32348
rect -34896 32268 -34849 32332
rect -34785 32268 -34769 32332
rect -34896 32252 -34769 32268
rect -34896 32188 -34849 32252
rect -34785 32188 -34769 32252
rect -34896 32172 -34769 32188
rect -34896 32108 -34849 32172
rect -34785 32108 -34769 32172
rect -34896 32092 -34769 32108
rect -34896 32028 -34849 32092
rect -34785 32028 -34769 32092
rect -34896 32012 -34769 32028
rect -34896 31948 -34849 32012
rect -34785 31948 -34769 32012
rect -34896 31932 -34769 31948
rect -34896 31868 -34849 31932
rect -34785 31868 -34769 31932
rect -34896 31852 -34769 31868
rect -34896 31788 -34849 31852
rect -34785 31788 -34769 31852
rect -34896 31772 -34769 31788
rect -34896 31708 -34849 31772
rect -34785 31708 -34769 31772
rect -34896 31692 -34769 31708
rect -34896 31628 -34849 31692
rect -34785 31628 -34769 31692
rect -34896 31612 -34769 31628
rect -34896 31548 -34849 31612
rect -34785 31548 -34769 31612
rect -34896 31532 -34769 31548
rect -34896 31468 -34849 31532
rect -34785 31468 -34769 31532
rect -34896 31452 -34769 31468
rect -34896 31388 -34849 31452
rect -34785 31388 -34769 31452
rect -34896 31372 -34769 31388
rect -34896 31308 -34849 31372
rect -34785 31308 -34769 31372
rect -34896 31292 -34769 31308
rect -34896 31228 -34849 31292
rect -34785 31228 -34769 31292
rect -34896 31212 -34769 31228
rect -34896 31148 -34849 31212
rect -34785 31148 -34769 31212
rect -34896 31132 -34769 31148
rect -34896 31068 -34849 31132
rect -34785 31068 -34769 31132
rect -34896 31052 -34769 31068
rect -34896 30988 -34849 31052
rect -34785 30988 -34769 31052
rect -34896 30972 -34769 30988
rect -34896 30908 -34849 30972
rect -34785 30908 -34769 30972
rect -34896 30892 -34769 30908
rect -34896 30828 -34849 30892
rect -34785 30828 -34769 30892
rect -34896 30812 -34769 30828
rect -34896 30748 -34849 30812
rect -34785 30748 -34769 30812
rect -34896 30732 -34769 30748
rect -34896 30668 -34849 30732
rect -34785 30668 -34769 30732
rect -34896 30652 -34769 30668
rect -34896 30588 -34849 30652
rect -34785 30588 -34769 30652
rect -34896 30572 -34769 30588
rect -34896 30508 -34849 30572
rect -34785 30508 -34769 30572
rect -34896 30492 -34769 30508
rect -34896 30428 -34849 30492
rect -34785 30428 -34769 30492
rect -34896 30412 -34769 30428
rect -34896 30348 -34849 30412
rect -34785 30348 -34769 30412
rect -34896 30332 -34769 30348
rect -34896 30268 -34849 30332
rect -34785 30268 -34769 30332
rect -34896 30252 -34769 30268
rect -34896 30188 -34849 30252
rect -34785 30188 -34769 30252
rect -34896 30172 -34769 30188
rect -34896 30108 -34849 30172
rect -34785 30108 -34769 30172
rect -34896 30092 -34769 30108
rect -34896 30028 -34849 30092
rect -34785 30028 -34769 30092
rect -34896 30012 -34769 30028
rect -34896 29948 -34849 30012
rect -34785 29948 -34769 30012
rect -34896 29932 -34769 29948
rect -34896 29868 -34849 29932
rect -34785 29868 -34769 29932
rect -34896 29852 -34769 29868
rect -34896 29788 -34849 29852
rect -34785 29788 -34769 29852
rect -34896 29772 -34769 29788
rect -34896 29708 -34849 29772
rect -34785 29708 -34769 29772
rect -34896 29692 -34769 29708
rect -34896 29628 -34849 29692
rect -34785 29628 -34769 29692
rect -34896 29612 -34769 29628
rect -34896 29548 -34849 29612
rect -34785 29548 -34769 29612
rect -34896 29532 -34769 29548
rect -34896 29468 -34849 29532
rect -34785 29468 -34769 29532
rect -34896 29452 -34769 29468
rect -34896 29388 -34849 29452
rect -34785 29388 -34769 29452
rect -34896 29372 -34769 29388
rect -34896 29308 -34849 29372
rect -34785 29308 -34769 29372
rect -34896 29292 -34769 29308
rect -34896 29228 -34849 29292
rect -34785 29228 -34769 29292
rect -34896 29212 -34769 29228
rect -34896 29148 -34849 29212
rect -34785 29148 -34769 29212
rect -34896 29132 -34769 29148
rect -34896 29068 -34849 29132
rect -34785 29068 -34769 29132
rect -34896 29052 -34769 29068
rect -34896 28988 -34849 29052
rect -34785 28988 -34769 29052
rect -34896 28972 -34769 28988
rect -34896 28908 -34849 28972
rect -34785 28908 -34769 28972
rect -34896 28892 -34769 28908
rect -34896 28828 -34849 28892
rect -34785 28828 -34769 28892
rect -34896 28812 -34769 28828
rect -34896 28748 -34849 28812
rect -34785 28748 -34769 28812
rect -34896 28732 -34769 28748
rect -34896 28668 -34849 28732
rect -34785 28668 -34769 28732
rect -34896 28652 -34769 28668
rect -34896 28588 -34849 28652
rect -34785 28588 -34769 28652
rect -34896 28572 -34769 28588
rect -41215 28492 -41088 28508
rect -41215 28428 -41168 28492
rect -41104 28428 -41088 28492
rect -41215 28412 -41088 28428
rect -41215 28288 -41111 28412
rect -41215 28272 -41088 28288
rect -41215 28208 -41168 28272
rect -41104 28208 -41088 28272
rect -41215 28192 -41088 28208
rect -47244 28152 -41322 28161
rect -47244 22248 -47235 28152
rect -41331 22248 -41322 28152
rect -47244 22239 -41322 22248
rect -41215 28128 -41168 28192
rect -41104 28128 -41088 28192
rect -38016 28161 -37912 28539
rect -34896 28508 -34849 28572
rect -34785 28508 -34769 28572
rect -34606 34452 -28684 34461
rect -34606 28548 -34597 34452
rect -28693 28548 -28684 34452
rect -34606 28539 -28684 28548
rect -28577 34428 -28530 34492
rect -28466 34428 -28450 34492
rect -25378 34461 -25274 34839
rect -22258 34808 -22211 34872
rect -22147 34808 -22131 34872
rect -21968 40752 -16046 40761
rect -21968 34848 -21959 40752
rect -16055 34848 -16046 40752
rect -21968 34839 -16046 34848
rect -15939 40728 -15892 40792
rect -15828 40728 -15812 40792
rect -12740 40761 -12636 41139
rect -9620 41108 -9573 41172
rect -9509 41108 -9493 41172
rect -9330 47052 -3408 47061
rect -9330 41148 -9321 47052
rect -3417 41148 -3408 47052
rect -9330 41139 -3408 41148
rect -3301 47028 -3254 47092
rect -3190 47028 -3174 47092
rect -102 47061 2 47250
rect 3018 47188 3122 47250
rect 3018 47172 3145 47188
rect 3018 47108 3065 47172
rect 3129 47108 3145 47172
rect 3018 47092 3145 47108
rect -3301 47012 -3174 47028
rect -3301 46948 -3254 47012
rect -3190 46948 -3174 47012
rect -3301 46932 -3174 46948
rect -3301 46868 -3254 46932
rect -3190 46868 -3174 46932
rect -3301 46852 -3174 46868
rect -3301 46788 -3254 46852
rect -3190 46788 -3174 46852
rect -3301 46772 -3174 46788
rect -3301 46708 -3254 46772
rect -3190 46708 -3174 46772
rect -3301 46692 -3174 46708
rect -3301 46628 -3254 46692
rect -3190 46628 -3174 46692
rect -3301 46612 -3174 46628
rect -3301 46548 -3254 46612
rect -3190 46548 -3174 46612
rect -3301 46532 -3174 46548
rect -3301 46468 -3254 46532
rect -3190 46468 -3174 46532
rect -3301 46452 -3174 46468
rect -3301 46388 -3254 46452
rect -3190 46388 -3174 46452
rect -3301 46372 -3174 46388
rect -3301 46308 -3254 46372
rect -3190 46308 -3174 46372
rect -3301 46292 -3174 46308
rect -3301 46228 -3254 46292
rect -3190 46228 -3174 46292
rect -3301 46212 -3174 46228
rect -3301 46148 -3254 46212
rect -3190 46148 -3174 46212
rect -3301 46132 -3174 46148
rect -3301 46068 -3254 46132
rect -3190 46068 -3174 46132
rect -3301 46052 -3174 46068
rect -3301 45988 -3254 46052
rect -3190 45988 -3174 46052
rect -3301 45972 -3174 45988
rect -3301 45908 -3254 45972
rect -3190 45908 -3174 45972
rect -3301 45892 -3174 45908
rect -3301 45828 -3254 45892
rect -3190 45828 -3174 45892
rect -3301 45812 -3174 45828
rect -3301 45748 -3254 45812
rect -3190 45748 -3174 45812
rect -3301 45732 -3174 45748
rect -3301 45668 -3254 45732
rect -3190 45668 -3174 45732
rect -3301 45652 -3174 45668
rect -3301 45588 -3254 45652
rect -3190 45588 -3174 45652
rect -3301 45572 -3174 45588
rect -3301 45508 -3254 45572
rect -3190 45508 -3174 45572
rect -3301 45492 -3174 45508
rect -3301 45428 -3254 45492
rect -3190 45428 -3174 45492
rect -3301 45412 -3174 45428
rect -3301 45348 -3254 45412
rect -3190 45348 -3174 45412
rect -3301 45332 -3174 45348
rect -3301 45268 -3254 45332
rect -3190 45268 -3174 45332
rect -3301 45252 -3174 45268
rect -3301 45188 -3254 45252
rect -3190 45188 -3174 45252
rect -3301 45172 -3174 45188
rect -3301 45108 -3254 45172
rect -3190 45108 -3174 45172
rect -3301 45092 -3174 45108
rect -3301 45028 -3254 45092
rect -3190 45028 -3174 45092
rect -3301 45012 -3174 45028
rect -3301 44948 -3254 45012
rect -3190 44948 -3174 45012
rect -3301 44932 -3174 44948
rect -3301 44868 -3254 44932
rect -3190 44868 -3174 44932
rect -3301 44852 -3174 44868
rect -3301 44788 -3254 44852
rect -3190 44788 -3174 44852
rect -3301 44772 -3174 44788
rect -3301 44708 -3254 44772
rect -3190 44708 -3174 44772
rect -3301 44692 -3174 44708
rect -3301 44628 -3254 44692
rect -3190 44628 -3174 44692
rect -3301 44612 -3174 44628
rect -3301 44548 -3254 44612
rect -3190 44548 -3174 44612
rect -3301 44532 -3174 44548
rect -3301 44468 -3254 44532
rect -3190 44468 -3174 44532
rect -3301 44452 -3174 44468
rect -3301 44388 -3254 44452
rect -3190 44388 -3174 44452
rect -3301 44372 -3174 44388
rect -3301 44308 -3254 44372
rect -3190 44308 -3174 44372
rect -3301 44292 -3174 44308
rect -3301 44228 -3254 44292
rect -3190 44228 -3174 44292
rect -3301 44212 -3174 44228
rect -3301 44148 -3254 44212
rect -3190 44148 -3174 44212
rect -3301 44132 -3174 44148
rect -3301 44068 -3254 44132
rect -3190 44068 -3174 44132
rect -3301 44052 -3174 44068
rect -3301 43988 -3254 44052
rect -3190 43988 -3174 44052
rect -3301 43972 -3174 43988
rect -3301 43908 -3254 43972
rect -3190 43908 -3174 43972
rect -3301 43892 -3174 43908
rect -3301 43828 -3254 43892
rect -3190 43828 -3174 43892
rect -3301 43812 -3174 43828
rect -3301 43748 -3254 43812
rect -3190 43748 -3174 43812
rect -3301 43732 -3174 43748
rect -3301 43668 -3254 43732
rect -3190 43668 -3174 43732
rect -3301 43652 -3174 43668
rect -3301 43588 -3254 43652
rect -3190 43588 -3174 43652
rect -3301 43572 -3174 43588
rect -3301 43508 -3254 43572
rect -3190 43508 -3174 43572
rect -3301 43492 -3174 43508
rect -3301 43428 -3254 43492
rect -3190 43428 -3174 43492
rect -3301 43412 -3174 43428
rect -3301 43348 -3254 43412
rect -3190 43348 -3174 43412
rect -3301 43332 -3174 43348
rect -3301 43268 -3254 43332
rect -3190 43268 -3174 43332
rect -3301 43252 -3174 43268
rect -3301 43188 -3254 43252
rect -3190 43188 -3174 43252
rect -3301 43172 -3174 43188
rect -3301 43108 -3254 43172
rect -3190 43108 -3174 43172
rect -3301 43092 -3174 43108
rect -3301 43028 -3254 43092
rect -3190 43028 -3174 43092
rect -3301 43012 -3174 43028
rect -3301 42948 -3254 43012
rect -3190 42948 -3174 43012
rect -3301 42932 -3174 42948
rect -3301 42868 -3254 42932
rect -3190 42868 -3174 42932
rect -3301 42852 -3174 42868
rect -3301 42788 -3254 42852
rect -3190 42788 -3174 42852
rect -3301 42772 -3174 42788
rect -3301 42708 -3254 42772
rect -3190 42708 -3174 42772
rect -3301 42692 -3174 42708
rect -3301 42628 -3254 42692
rect -3190 42628 -3174 42692
rect -3301 42612 -3174 42628
rect -3301 42548 -3254 42612
rect -3190 42548 -3174 42612
rect -3301 42532 -3174 42548
rect -3301 42468 -3254 42532
rect -3190 42468 -3174 42532
rect -3301 42452 -3174 42468
rect -3301 42388 -3254 42452
rect -3190 42388 -3174 42452
rect -3301 42372 -3174 42388
rect -3301 42308 -3254 42372
rect -3190 42308 -3174 42372
rect -3301 42292 -3174 42308
rect -3301 42228 -3254 42292
rect -3190 42228 -3174 42292
rect -3301 42212 -3174 42228
rect -3301 42148 -3254 42212
rect -3190 42148 -3174 42212
rect -3301 42132 -3174 42148
rect -3301 42068 -3254 42132
rect -3190 42068 -3174 42132
rect -3301 42052 -3174 42068
rect -3301 41988 -3254 42052
rect -3190 41988 -3174 42052
rect -3301 41972 -3174 41988
rect -3301 41908 -3254 41972
rect -3190 41908 -3174 41972
rect -3301 41892 -3174 41908
rect -3301 41828 -3254 41892
rect -3190 41828 -3174 41892
rect -3301 41812 -3174 41828
rect -3301 41748 -3254 41812
rect -3190 41748 -3174 41812
rect -3301 41732 -3174 41748
rect -3301 41668 -3254 41732
rect -3190 41668 -3174 41732
rect -3301 41652 -3174 41668
rect -3301 41588 -3254 41652
rect -3190 41588 -3174 41652
rect -3301 41572 -3174 41588
rect -3301 41508 -3254 41572
rect -3190 41508 -3174 41572
rect -3301 41492 -3174 41508
rect -3301 41428 -3254 41492
rect -3190 41428 -3174 41492
rect -3301 41412 -3174 41428
rect -3301 41348 -3254 41412
rect -3190 41348 -3174 41412
rect -3301 41332 -3174 41348
rect -3301 41268 -3254 41332
rect -3190 41268 -3174 41332
rect -3301 41252 -3174 41268
rect -3301 41188 -3254 41252
rect -3190 41188 -3174 41252
rect -3301 41172 -3174 41188
rect -9620 41092 -9493 41108
rect -9620 41028 -9573 41092
rect -9509 41028 -9493 41092
rect -9620 41012 -9493 41028
rect -9620 40888 -9516 41012
rect -9620 40872 -9493 40888
rect -9620 40808 -9573 40872
rect -9509 40808 -9493 40872
rect -9620 40792 -9493 40808
rect -15939 40712 -15812 40728
rect -15939 40648 -15892 40712
rect -15828 40648 -15812 40712
rect -15939 40632 -15812 40648
rect -15939 40568 -15892 40632
rect -15828 40568 -15812 40632
rect -15939 40552 -15812 40568
rect -15939 40488 -15892 40552
rect -15828 40488 -15812 40552
rect -15939 40472 -15812 40488
rect -15939 40408 -15892 40472
rect -15828 40408 -15812 40472
rect -15939 40392 -15812 40408
rect -15939 40328 -15892 40392
rect -15828 40328 -15812 40392
rect -15939 40312 -15812 40328
rect -15939 40248 -15892 40312
rect -15828 40248 -15812 40312
rect -15939 40232 -15812 40248
rect -15939 40168 -15892 40232
rect -15828 40168 -15812 40232
rect -15939 40152 -15812 40168
rect -15939 40088 -15892 40152
rect -15828 40088 -15812 40152
rect -15939 40072 -15812 40088
rect -15939 40008 -15892 40072
rect -15828 40008 -15812 40072
rect -15939 39992 -15812 40008
rect -15939 39928 -15892 39992
rect -15828 39928 -15812 39992
rect -15939 39912 -15812 39928
rect -15939 39848 -15892 39912
rect -15828 39848 -15812 39912
rect -15939 39832 -15812 39848
rect -15939 39768 -15892 39832
rect -15828 39768 -15812 39832
rect -15939 39752 -15812 39768
rect -15939 39688 -15892 39752
rect -15828 39688 -15812 39752
rect -15939 39672 -15812 39688
rect -15939 39608 -15892 39672
rect -15828 39608 -15812 39672
rect -15939 39592 -15812 39608
rect -15939 39528 -15892 39592
rect -15828 39528 -15812 39592
rect -15939 39512 -15812 39528
rect -15939 39448 -15892 39512
rect -15828 39448 -15812 39512
rect -15939 39432 -15812 39448
rect -15939 39368 -15892 39432
rect -15828 39368 -15812 39432
rect -15939 39352 -15812 39368
rect -15939 39288 -15892 39352
rect -15828 39288 -15812 39352
rect -15939 39272 -15812 39288
rect -15939 39208 -15892 39272
rect -15828 39208 -15812 39272
rect -15939 39192 -15812 39208
rect -15939 39128 -15892 39192
rect -15828 39128 -15812 39192
rect -15939 39112 -15812 39128
rect -15939 39048 -15892 39112
rect -15828 39048 -15812 39112
rect -15939 39032 -15812 39048
rect -15939 38968 -15892 39032
rect -15828 38968 -15812 39032
rect -15939 38952 -15812 38968
rect -15939 38888 -15892 38952
rect -15828 38888 -15812 38952
rect -15939 38872 -15812 38888
rect -15939 38808 -15892 38872
rect -15828 38808 -15812 38872
rect -15939 38792 -15812 38808
rect -15939 38728 -15892 38792
rect -15828 38728 -15812 38792
rect -15939 38712 -15812 38728
rect -15939 38648 -15892 38712
rect -15828 38648 -15812 38712
rect -15939 38632 -15812 38648
rect -15939 38568 -15892 38632
rect -15828 38568 -15812 38632
rect -15939 38552 -15812 38568
rect -15939 38488 -15892 38552
rect -15828 38488 -15812 38552
rect -15939 38472 -15812 38488
rect -15939 38408 -15892 38472
rect -15828 38408 -15812 38472
rect -15939 38392 -15812 38408
rect -15939 38328 -15892 38392
rect -15828 38328 -15812 38392
rect -15939 38312 -15812 38328
rect -15939 38248 -15892 38312
rect -15828 38248 -15812 38312
rect -15939 38232 -15812 38248
rect -15939 38168 -15892 38232
rect -15828 38168 -15812 38232
rect -15939 38152 -15812 38168
rect -15939 38088 -15892 38152
rect -15828 38088 -15812 38152
rect -15939 38072 -15812 38088
rect -15939 38008 -15892 38072
rect -15828 38008 -15812 38072
rect -15939 37992 -15812 38008
rect -15939 37928 -15892 37992
rect -15828 37928 -15812 37992
rect -15939 37912 -15812 37928
rect -15939 37848 -15892 37912
rect -15828 37848 -15812 37912
rect -15939 37832 -15812 37848
rect -15939 37768 -15892 37832
rect -15828 37768 -15812 37832
rect -15939 37752 -15812 37768
rect -15939 37688 -15892 37752
rect -15828 37688 -15812 37752
rect -15939 37672 -15812 37688
rect -15939 37608 -15892 37672
rect -15828 37608 -15812 37672
rect -15939 37592 -15812 37608
rect -15939 37528 -15892 37592
rect -15828 37528 -15812 37592
rect -15939 37512 -15812 37528
rect -15939 37448 -15892 37512
rect -15828 37448 -15812 37512
rect -15939 37432 -15812 37448
rect -15939 37368 -15892 37432
rect -15828 37368 -15812 37432
rect -15939 37352 -15812 37368
rect -15939 37288 -15892 37352
rect -15828 37288 -15812 37352
rect -15939 37272 -15812 37288
rect -15939 37208 -15892 37272
rect -15828 37208 -15812 37272
rect -15939 37192 -15812 37208
rect -15939 37128 -15892 37192
rect -15828 37128 -15812 37192
rect -15939 37112 -15812 37128
rect -15939 37048 -15892 37112
rect -15828 37048 -15812 37112
rect -15939 37032 -15812 37048
rect -15939 36968 -15892 37032
rect -15828 36968 -15812 37032
rect -15939 36952 -15812 36968
rect -15939 36888 -15892 36952
rect -15828 36888 -15812 36952
rect -15939 36872 -15812 36888
rect -15939 36808 -15892 36872
rect -15828 36808 -15812 36872
rect -15939 36792 -15812 36808
rect -15939 36728 -15892 36792
rect -15828 36728 -15812 36792
rect -15939 36712 -15812 36728
rect -15939 36648 -15892 36712
rect -15828 36648 -15812 36712
rect -15939 36632 -15812 36648
rect -15939 36568 -15892 36632
rect -15828 36568 -15812 36632
rect -15939 36552 -15812 36568
rect -15939 36488 -15892 36552
rect -15828 36488 -15812 36552
rect -15939 36472 -15812 36488
rect -15939 36408 -15892 36472
rect -15828 36408 -15812 36472
rect -15939 36392 -15812 36408
rect -15939 36328 -15892 36392
rect -15828 36328 -15812 36392
rect -15939 36312 -15812 36328
rect -15939 36248 -15892 36312
rect -15828 36248 -15812 36312
rect -15939 36232 -15812 36248
rect -15939 36168 -15892 36232
rect -15828 36168 -15812 36232
rect -15939 36152 -15812 36168
rect -15939 36088 -15892 36152
rect -15828 36088 -15812 36152
rect -15939 36072 -15812 36088
rect -15939 36008 -15892 36072
rect -15828 36008 -15812 36072
rect -15939 35992 -15812 36008
rect -15939 35928 -15892 35992
rect -15828 35928 -15812 35992
rect -15939 35912 -15812 35928
rect -15939 35848 -15892 35912
rect -15828 35848 -15812 35912
rect -15939 35832 -15812 35848
rect -15939 35768 -15892 35832
rect -15828 35768 -15812 35832
rect -15939 35752 -15812 35768
rect -15939 35688 -15892 35752
rect -15828 35688 -15812 35752
rect -15939 35672 -15812 35688
rect -15939 35608 -15892 35672
rect -15828 35608 -15812 35672
rect -15939 35592 -15812 35608
rect -15939 35528 -15892 35592
rect -15828 35528 -15812 35592
rect -15939 35512 -15812 35528
rect -15939 35448 -15892 35512
rect -15828 35448 -15812 35512
rect -15939 35432 -15812 35448
rect -15939 35368 -15892 35432
rect -15828 35368 -15812 35432
rect -15939 35352 -15812 35368
rect -15939 35288 -15892 35352
rect -15828 35288 -15812 35352
rect -15939 35272 -15812 35288
rect -15939 35208 -15892 35272
rect -15828 35208 -15812 35272
rect -15939 35192 -15812 35208
rect -15939 35128 -15892 35192
rect -15828 35128 -15812 35192
rect -15939 35112 -15812 35128
rect -15939 35048 -15892 35112
rect -15828 35048 -15812 35112
rect -15939 35032 -15812 35048
rect -15939 34968 -15892 35032
rect -15828 34968 -15812 35032
rect -15939 34952 -15812 34968
rect -15939 34888 -15892 34952
rect -15828 34888 -15812 34952
rect -15939 34872 -15812 34888
rect -22258 34792 -22131 34808
rect -22258 34728 -22211 34792
rect -22147 34728 -22131 34792
rect -22258 34712 -22131 34728
rect -22258 34588 -22154 34712
rect -22258 34572 -22131 34588
rect -22258 34508 -22211 34572
rect -22147 34508 -22131 34572
rect -22258 34492 -22131 34508
rect -28577 34412 -28450 34428
rect -28577 34348 -28530 34412
rect -28466 34348 -28450 34412
rect -28577 34332 -28450 34348
rect -28577 34268 -28530 34332
rect -28466 34268 -28450 34332
rect -28577 34252 -28450 34268
rect -28577 34188 -28530 34252
rect -28466 34188 -28450 34252
rect -28577 34172 -28450 34188
rect -28577 34108 -28530 34172
rect -28466 34108 -28450 34172
rect -28577 34092 -28450 34108
rect -28577 34028 -28530 34092
rect -28466 34028 -28450 34092
rect -28577 34012 -28450 34028
rect -28577 33948 -28530 34012
rect -28466 33948 -28450 34012
rect -28577 33932 -28450 33948
rect -28577 33868 -28530 33932
rect -28466 33868 -28450 33932
rect -28577 33852 -28450 33868
rect -28577 33788 -28530 33852
rect -28466 33788 -28450 33852
rect -28577 33772 -28450 33788
rect -28577 33708 -28530 33772
rect -28466 33708 -28450 33772
rect -28577 33692 -28450 33708
rect -28577 33628 -28530 33692
rect -28466 33628 -28450 33692
rect -28577 33612 -28450 33628
rect -28577 33548 -28530 33612
rect -28466 33548 -28450 33612
rect -28577 33532 -28450 33548
rect -28577 33468 -28530 33532
rect -28466 33468 -28450 33532
rect -28577 33452 -28450 33468
rect -28577 33388 -28530 33452
rect -28466 33388 -28450 33452
rect -28577 33372 -28450 33388
rect -28577 33308 -28530 33372
rect -28466 33308 -28450 33372
rect -28577 33292 -28450 33308
rect -28577 33228 -28530 33292
rect -28466 33228 -28450 33292
rect -28577 33212 -28450 33228
rect -28577 33148 -28530 33212
rect -28466 33148 -28450 33212
rect -28577 33132 -28450 33148
rect -28577 33068 -28530 33132
rect -28466 33068 -28450 33132
rect -28577 33052 -28450 33068
rect -28577 32988 -28530 33052
rect -28466 32988 -28450 33052
rect -28577 32972 -28450 32988
rect -28577 32908 -28530 32972
rect -28466 32908 -28450 32972
rect -28577 32892 -28450 32908
rect -28577 32828 -28530 32892
rect -28466 32828 -28450 32892
rect -28577 32812 -28450 32828
rect -28577 32748 -28530 32812
rect -28466 32748 -28450 32812
rect -28577 32732 -28450 32748
rect -28577 32668 -28530 32732
rect -28466 32668 -28450 32732
rect -28577 32652 -28450 32668
rect -28577 32588 -28530 32652
rect -28466 32588 -28450 32652
rect -28577 32572 -28450 32588
rect -28577 32508 -28530 32572
rect -28466 32508 -28450 32572
rect -28577 32492 -28450 32508
rect -28577 32428 -28530 32492
rect -28466 32428 -28450 32492
rect -28577 32412 -28450 32428
rect -28577 32348 -28530 32412
rect -28466 32348 -28450 32412
rect -28577 32332 -28450 32348
rect -28577 32268 -28530 32332
rect -28466 32268 -28450 32332
rect -28577 32252 -28450 32268
rect -28577 32188 -28530 32252
rect -28466 32188 -28450 32252
rect -28577 32172 -28450 32188
rect -28577 32108 -28530 32172
rect -28466 32108 -28450 32172
rect -28577 32092 -28450 32108
rect -28577 32028 -28530 32092
rect -28466 32028 -28450 32092
rect -28577 32012 -28450 32028
rect -28577 31948 -28530 32012
rect -28466 31948 -28450 32012
rect -28577 31932 -28450 31948
rect -28577 31868 -28530 31932
rect -28466 31868 -28450 31932
rect -28577 31852 -28450 31868
rect -28577 31788 -28530 31852
rect -28466 31788 -28450 31852
rect -28577 31772 -28450 31788
rect -28577 31708 -28530 31772
rect -28466 31708 -28450 31772
rect -28577 31692 -28450 31708
rect -28577 31628 -28530 31692
rect -28466 31628 -28450 31692
rect -28577 31612 -28450 31628
rect -28577 31548 -28530 31612
rect -28466 31548 -28450 31612
rect -28577 31532 -28450 31548
rect -28577 31468 -28530 31532
rect -28466 31468 -28450 31532
rect -28577 31452 -28450 31468
rect -28577 31388 -28530 31452
rect -28466 31388 -28450 31452
rect -28577 31372 -28450 31388
rect -28577 31308 -28530 31372
rect -28466 31308 -28450 31372
rect -28577 31292 -28450 31308
rect -28577 31228 -28530 31292
rect -28466 31228 -28450 31292
rect -28577 31212 -28450 31228
rect -28577 31148 -28530 31212
rect -28466 31148 -28450 31212
rect -28577 31132 -28450 31148
rect -28577 31068 -28530 31132
rect -28466 31068 -28450 31132
rect -28577 31052 -28450 31068
rect -28577 30988 -28530 31052
rect -28466 30988 -28450 31052
rect -28577 30972 -28450 30988
rect -28577 30908 -28530 30972
rect -28466 30908 -28450 30972
rect -28577 30892 -28450 30908
rect -28577 30828 -28530 30892
rect -28466 30828 -28450 30892
rect -28577 30812 -28450 30828
rect -28577 30748 -28530 30812
rect -28466 30748 -28450 30812
rect -28577 30732 -28450 30748
rect -28577 30668 -28530 30732
rect -28466 30668 -28450 30732
rect -28577 30652 -28450 30668
rect -28577 30588 -28530 30652
rect -28466 30588 -28450 30652
rect -28577 30572 -28450 30588
rect -28577 30508 -28530 30572
rect -28466 30508 -28450 30572
rect -28577 30492 -28450 30508
rect -28577 30428 -28530 30492
rect -28466 30428 -28450 30492
rect -28577 30412 -28450 30428
rect -28577 30348 -28530 30412
rect -28466 30348 -28450 30412
rect -28577 30332 -28450 30348
rect -28577 30268 -28530 30332
rect -28466 30268 -28450 30332
rect -28577 30252 -28450 30268
rect -28577 30188 -28530 30252
rect -28466 30188 -28450 30252
rect -28577 30172 -28450 30188
rect -28577 30108 -28530 30172
rect -28466 30108 -28450 30172
rect -28577 30092 -28450 30108
rect -28577 30028 -28530 30092
rect -28466 30028 -28450 30092
rect -28577 30012 -28450 30028
rect -28577 29948 -28530 30012
rect -28466 29948 -28450 30012
rect -28577 29932 -28450 29948
rect -28577 29868 -28530 29932
rect -28466 29868 -28450 29932
rect -28577 29852 -28450 29868
rect -28577 29788 -28530 29852
rect -28466 29788 -28450 29852
rect -28577 29772 -28450 29788
rect -28577 29708 -28530 29772
rect -28466 29708 -28450 29772
rect -28577 29692 -28450 29708
rect -28577 29628 -28530 29692
rect -28466 29628 -28450 29692
rect -28577 29612 -28450 29628
rect -28577 29548 -28530 29612
rect -28466 29548 -28450 29612
rect -28577 29532 -28450 29548
rect -28577 29468 -28530 29532
rect -28466 29468 -28450 29532
rect -28577 29452 -28450 29468
rect -28577 29388 -28530 29452
rect -28466 29388 -28450 29452
rect -28577 29372 -28450 29388
rect -28577 29308 -28530 29372
rect -28466 29308 -28450 29372
rect -28577 29292 -28450 29308
rect -28577 29228 -28530 29292
rect -28466 29228 -28450 29292
rect -28577 29212 -28450 29228
rect -28577 29148 -28530 29212
rect -28466 29148 -28450 29212
rect -28577 29132 -28450 29148
rect -28577 29068 -28530 29132
rect -28466 29068 -28450 29132
rect -28577 29052 -28450 29068
rect -28577 28988 -28530 29052
rect -28466 28988 -28450 29052
rect -28577 28972 -28450 28988
rect -28577 28908 -28530 28972
rect -28466 28908 -28450 28972
rect -28577 28892 -28450 28908
rect -28577 28828 -28530 28892
rect -28466 28828 -28450 28892
rect -28577 28812 -28450 28828
rect -28577 28748 -28530 28812
rect -28466 28748 -28450 28812
rect -28577 28732 -28450 28748
rect -28577 28668 -28530 28732
rect -28466 28668 -28450 28732
rect -28577 28652 -28450 28668
rect -28577 28588 -28530 28652
rect -28466 28588 -28450 28652
rect -28577 28572 -28450 28588
rect -34896 28492 -34769 28508
rect -34896 28428 -34849 28492
rect -34785 28428 -34769 28492
rect -34896 28412 -34769 28428
rect -34896 28288 -34792 28412
rect -34896 28272 -34769 28288
rect -34896 28208 -34849 28272
rect -34785 28208 -34769 28272
rect -34896 28192 -34769 28208
rect -41215 28112 -41088 28128
rect -41215 28048 -41168 28112
rect -41104 28048 -41088 28112
rect -41215 28032 -41088 28048
rect -41215 27968 -41168 28032
rect -41104 27968 -41088 28032
rect -41215 27952 -41088 27968
rect -41215 27888 -41168 27952
rect -41104 27888 -41088 27952
rect -41215 27872 -41088 27888
rect -41215 27808 -41168 27872
rect -41104 27808 -41088 27872
rect -41215 27792 -41088 27808
rect -41215 27728 -41168 27792
rect -41104 27728 -41088 27792
rect -41215 27712 -41088 27728
rect -41215 27648 -41168 27712
rect -41104 27648 -41088 27712
rect -41215 27632 -41088 27648
rect -41215 27568 -41168 27632
rect -41104 27568 -41088 27632
rect -41215 27552 -41088 27568
rect -41215 27488 -41168 27552
rect -41104 27488 -41088 27552
rect -41215 27472 -41088 27488
rect -41215 27408 -41168 27472
rect -41104 27408 -41088 27472
rect -41215 27392 -41088 27408
rect -41215 27328 -41168 27392
rect -41104 27328 -41088 27392
rect -41215 27312 -41088 27328
rect -41215 27248 -41168 27312
rect -41104 27248 -41088 27312
rect -41215 27232 -41088 27248
rect -41215 27168 -41168 27232
rect -41104 27168 -41088 27232
rect -41215 27152 -41088 27168
rect -41215 27088 -41168 27152
rect -41104 27088 -41088 27152
rect -41215 27072 -41088 27088
rect -41215 27008 -41168 27072
rect -41104 27008 -41088 27072
rect -41215 26992 -41088 27008
rect -41215 26928 -41168 26992
rect -41104 26928 -41088 26992
rect -41215 26912 -41088 26928
rect -41215 26848 -41168 26912
rect -41104 26848 -41088 26912
rect -41215 26832 -41088 26848
rect -41215 26768 -41168 26832
rect -41104 26768 -41088 26832
rect -41215 26752 -41088 26768
rect -41215 26688 -41168 26752
rect -41104 26688 -41088 26752
rect -41215 26672 -41088 26688
rect -41215 26608 -41168 26672
rect -41104 26608 -41088 26672
rect -41215 26592 -41088 26608
rect -41215 26528 -41168 26592
rect -41104 26528 -41088 26592
rect -41215 26512 -41088 26528
rect -41215 26448 -41168 26512
rect -41104 26448 -41088 26512
rect -41215 26432 -41088 26448
rect -41215 26368 -41168 26432
rect -41104 26368 -41088 26432
rect -41215 26352 -41088 26368
rect -41215 26288 -41168 26352
rect -41104 26288 -41088 26352
rect -41215 26272 -41088 26288
rect -41215 26208 -41168 26272
rect -41104 26208 -41088 26272
rect -41215 26192 -41088 26208
rect -41215 26128 -41168 26192
rect -41104 26128 -41088 26192
rect -41215 26112 -41088 26128
rect -41215 26048 -41168 26112
rect -41104 26048 -41088 26112
rect -41215 26032 -41088 26048
rect -41215 25968 -41168 26032
rect -41104 25968 -41088 26032
rect -41215 25952 -41088 25968
rect -41215 25888 -41168 25952
rect -41104 25888 -41088 25952
rect -41215 25872 -41088 25888
rect -41215 25808 -41168 25872
rect -41104 25808 -41088 25872
rect -41215 25792 -41088 25808
rect -41215 25728 -41168 25792
rect -41104 25728 -41088 25792
rect -41215 25712 -41088 25728
rect -41215 25648 -41168 25712
rect -41104 25648 -41088 25712
rect -41215 25632 -41088 25648
rect -41215 25568 -41168 25632
rect -41104 25568 -41088 25632
rect -41215 25552 -41088 25568
rect -41215 25488 -41168 25552
rect -41104 25488 -41088 25552
rect -41215 25472 -41088 25488
rect -41215 25408 -41168 25472
rect -41104 25408 -41088 25472
rect -41215 25392 -41088 25408
rect -41215 25328 -41168 25392
rect -41104 25328 -41088 25392
rect -41215 25312 -41088 25328
rect -41215 25248 -41168 25312
rect -41104 25248 -41088 25312
rect -41215 25232 -41088 25248
rect -41215 25168 -41168 25232
rect -41104 25168 -41088 25232
rect -41215 25152 -41088 25168
rect -41215 25088 -41168 25152
rect -41104 25088 -41088 25152
rect -41215 25072 -41088 25088
rect -41215 25008 -41168 25072
rect -41104 25008 -41088 25072
rect -41215 24992 -41088 25008
rect -41215 24928 -41168 24992
rect -41104 24928 -41088 24992
rect -41215 24912 -41088 24928
rect -41215 24848 -41168 24912
rect -41104 24848 -41088 24912
rect -41215 24832 -41088 24848
rect -41215 24768 -41168 24832
rect -41104 24768 -41088 24832
rect -41215 24752 -41088 24768
rect -41215 24688 -41168 24752
rect -41104 24688 -41088 24752
rect -41215 24672 -41088 24688
rect -41215 24608 -41168 24672
rect -41104 24608 -41088 24672
rect -41215 24592 -41088 24608
rect -41215 24528 -41168 24592
rect -41104 24528 -41088 24592
rect -41215 24512 -41088 24528
rect -41215 24448 -41168 24512
rect -41104 24448 -41088 24512
rect -41215 24432 -41088 24448
rect -41215 24368 -41168 24432
rect -41104 24368 -41088 24432
rect -41215 24352 -41088 24368
rect -41215 24288 -41168 24352
rect -41104 24288 -41088 24352
rect -41215 24272 -41088 24288
rect -41215 24208 -41168 24272
rect -41104 24208 -41088 24272
rect -41215 24192 -41088 24208
rect -41215 24128 -41168 24192
rect -41104 24128 -41088 24192
rect -41215 24112 -41088 24128
rect -41215 24048 -41168 24112
rect -41104 24048 -41088 24112
rect -41215 24032 -41088 24048
rect -41215 23968 -41168 24032
rect -41104 23968 -41088 24032
rect -41215 23952 -41088 23968
rect -41215 23888 -41168 23952
rect -41104 23888 -41088 23952
rect -41215 23872 -41088 23888
rect -41215 23808 -41168 23872
rect -41104 23808 -41088 23872
rect -41215 23792 -41088 23808
rect -41215 23728 -41168 23792
rect -41104 23728 -41088 23792
rect -41215 23712 -41088 23728
rect -41215 23648 -41168 23712
rect -41104 23648 -41088 23712
rect -41215 23632 -41088 23648
rect -41215 23568 -41168 23632
rect -41104 23568 -41088 23632
rect -41215 23552 -41088 23568
rect -41215 23488 -41168 23552
rect -41104 23488 -41088 23552
rect -41215 23472 -41088 23488
rect -41215 23408 -41168 23472
rect -41104 23408 -41088 23472
rect -41215 23392 -41088 23408
rect -41215 23328 -41168 23392
rect -41104 23328 -41088 23392
rect -41215 23312 -41088 23328
rect -41215 23248 -41168 23312
rect -41104 23248 -41088 23312
rect -41215 23232 -41088 23248
rect -41215 23168 -41168 23232
rect -41104 23168 -41088 23232
rect -41215 23152 -41088 23168
rect -41215 23088 -41168 23152
rect -41104 23088 -41088 23152
rect -41215 23072 -41088 23088
rect -41215 23008 -41168 23072
rect -41104 23008 -41088 23072
rect -41215 22992 -41088 23008
rect -41215 22928 -41168 22992
rect -41104 22928 -41088 22992
rect -41215 22912 -41088 22928
rect -41215 22848 -41168 22912
rect -41104 22848 -41088 22912
rect -41215 22832 -41088 22848
rect -41215 22768 -41168 22832
rect -41104 22768 -41088 22832
rect -41215 22752 -41088 22768
rect -41215 22688 -41168 22752
rect -41104 22688 -41088 22752
rect -41215 22672 -41088 22688
rect -41215 22608 -41168 22672
rect -41104 22608 -41088 22672
rect -41215 22592 -41088 22608
rect -41215 22528 -41168 22592
rect -41104 22528 -41088 22592
rect -41215 22512 -41088 22528
rect -41215 22448 -41168 22512
rect -41104 22448 -41088 22512
rect -41215 22432 -41088 22448
rect -41215 22368 -41168 22432
rect -41104 22368 -41088 22432
rect -41215 22352 -41088 22368
rect -41215 22288 -41168 22352
rect -41104 22288 -41088 22352
rect -41215 22272 -41088 22288
rect -44335 21861 -44231 22239
rect -41215 22208 -41168 22272
rect -41104 22208 -41088 22272
rect -40925 28152 -35003 28161
rect -40925 22248 -40916 28152
rect -35012 22248 -35003 28152
rect -40925 22239 -35003 22248
rect -34896 28128 -34849 28192
rect -34785 28128 -34769 28192
rect -31697 28161 -31593 28539
rect -28577 28508 -28530 28572
rect -28466 28508 -28450 28572
rect -28287 34452 -22365 34461
rect -28287 28548 -28278 34452
rect -22374 28548 -22365 34452
rect -28287 28539 -22365 28548
rect -22258 34428 -22211 34492
rect -22147 34428 -22131 34492
rect -19059 34461 -18955 34839
rect -15939 34808 -15892 34872
rect -15828 34808 -15812 34872
rect -15649 40752 -9727 40761
rect -15649 34848 -15640 40752
rect -9736 34848 -9727 40752
rect -15649 34839 -9727 34848
rect -9620 40728 -9573 40792
rect -9509 40728 -9493 40792
rect -6421 40761 -6317 41139
rect -3301 41108 -3254 41172
rect -3190 41108 -3174 41172
rect -3011 47052 2911 47061
rect -3011 41148 -3002 47052
rect 2902 41148 2911 47052
rect -3011 41139 2911 41148
rect 3018 47028 3065 47092
rect 3129 47028 3145 47092
rect 6217 47061 6321 47250
rect 9337 47188 9441 47250
rect 9337 47172 9464 47188
rect 9337 47108 9384 47172
rect 9448 47108 9464 47172
rect 9337 47092 9464 47108
rect 3018 47012 3145 47028
rect 3018 46948 3065 47012
rect 3129 46948 3145 47012
rect 3018 46932 3145 46948
rect 3018 46868 3065 46932
rect 3129 46868 3145 46932
rect 3018 46852 3145 46868
rect 3018 46788 3065 46852
rect 3129 46788 3145 46852
rect 3018 46772 3145 46788
rect 3018 46708 3065 46772
rect 3129 46708 3145 46772
rect 3018 46692 3145 46708
rect 3018 46628 3065 46692
rect 3129 46628 3145 46692
rect 3018 46612 3145 46628
rect 3018 46548 3065 46612
rect 3129 46548 3145 46612
rect 3018 46532 3145 46548
rect 3018 46468 3065 46532
rect 3129 46468 3145 46532
rect 3018 46452 3145 46468
rect 3018 46388 3065 46452
rect 3129 46388 3145 46452
rect 3018 46372 3145 46388
rect 3018 46308 3065 46372
rect 3129 46308 3145 46372
rect 3018 46292 3145 46308
rect 3018 46228 3065 46292
rect 3129 46228 3145 46292
rect 3018 46212 3145 46228
rect 3018 46148 3065 46212
rect 3129 46148 3145 46212
rect 3018 46132 3145 46148
rect 3018 46068 3065 46132
rect 3129 46068 3145 46132
rect 3018 46052 3145 46068
rect 3018 45988 3065 46052
rect 3129 45988 3145 46052
rect 3018 45972 3145 45988
rect 3018 45908 3065 45972
rect 3129 45908 3145 45972
rect 3018 45892 3145 45908
rect 3018 45828 3065 45892
rect 3129 45828 3145 45892
rect 3018 45812 3145 45828
rect 3018 45748 3065 45812
rect 3129 45748 3145 45812
rect 3018 45732 3145 45748
rect 3018 45668 3065 45732
rect 3129 45668 3145 45732
rect 3018 45652 3145 45668
rect 3018 45588 3065 45652
rect 3129 45588 3145 45652
rect 3018 45572 3145 45588
rect 3018 45508 3065 45572
rect 3129 45508 3145 45572
rect 3018 45492 3145 45508
rect 3018 45428 3065 45492
rect 3129 45428 3145 45492
rect 3018 45412 3145 45428
rect 3018 45348 3065 45412
rect 3129 45348 3145 45412
rect 3018 45332 3145 45348
rect 3018 45268 3065 45332
rect 3129 45268 3145 45332
rect 3018 45252 3145 45268
rect 3018 45188 3065 45252
rect 3129 45188 3145 45252
rect 3018 45172 3145 45188
rect 3018 45108 3065 45172
rect 3129 45108 3145 45172
rect 3018 45092 3145 45108
rect 3018 45028 3065 45092
rect 3129 45028 3145 45092
rect 3018 45012 3145 45028
rect 3018 44948 3065 45012
rect 3129 44948 3145 45012
rect 3018 44932 3145 44948
rect 3018 44868 3065 44932
rect 3129 44868 3145 44932
rect 3018 44852 3145 44868
rect 3018 44788 3065 44852
rect 3129 44788 3145 44852
rect 3018 44772 3145 44788
rect 3018 44708 3065 44772
rect 3129 44708 3145 44772
rect 3018 44692 3145 44708
rect 3018 44628 3065 44692
rect 3129 44628 3145 44692
rect 3018 44612 3145 44628
rect 3018 44548 3065 44612
rect 3129 44548 3145 44612
rect 3018 44532 3145 44548
rect 3018 44468 3065 44532
rect 3129 44468 3145 44532
rect 3018 44452 3145 44468
rect 3018 44388 3065 44452
rect 3129 44388 3145 44452
rect 3018 44372 3145 44388
rect 3018 44308 3065 44372
rect 3129 44308 3145 44372
rect 3018 44292 3145 44308
rect 3018 44228 3065 44292
rect 3129 44228 3145 44292
rect 3018 44212 3145 44228
rect 3018 44148 3065 44212
rect 3129 44148 3145 44212
rect 3018 44132 3145 44148
rect 3018 44068 3065 44132
rect 3129 44068 3145 44132
rect 3018 44052 3145 44068
rect 3018 43988 3065 44052
rect 3129 43988 3145 44052
rect 3018 43972 3145 43988
rect 3018 43908 3065 43972
rect 3129 43908 3145 43972
rect 3018 43892 3145 43908
rect 3018 43828 3065 43892
rect 3129 43828 3145 43892
rect 3018 43812 3145 43828
rect 3018 43748 3065 43812
rect 3129 43748 3145 43812
rect 3018 43732 3145 43748
rect 3018 43668 3065 43732
rect 3129 43668 3145 43732
rect 3018 43652 3145 43668
rect 3018 43588 3065 43652
rect 3129 43588 3145 43652
rect 3018 43572 3145 43588
rect 3018 43508 3065 43572
rect 3129 43508 3145 43572
rect 3018 43492 3145 43508
rect 3018 43428 3065 43492
rect 3129 43428 3145 43492
rect 3018 43412 3145 43428
rect 3018 43348 3065 43412
rect 3129 43348 3145 43412
rect 3018 43332 3145 43348
rect 3018 43268 3065 43332
rect 3129 43268 3145 43332
rect 3018 43252 3145 43268
rect 3018 43188 3065 43252
rect 3129 43188 3145 43252
rect 3018 43172 3145 43188
rect 3018 43108 3065 43172
rect 3129 43108 3145 43172
rect 3018 43092 3145 43108
rect 3018 43028 3065 43092
rect 3129 43028 3145 43092
rect 3018 43012 3145 43028
rect 3018 42948 3065 43012
rect 3129 42948 3145 43012
rect 3018 42932 3145 42948
rect 3018 42868 3065 42932
rect 3129 42868 3145 42932
rect 3018 42852 3145 42868
rect 3018 42788 3065 42852
rect 3129 42788 3145 42852
rect 3018 42772 3145 42788
rect 3018 42708 3065 42772
rect 3129 42708 3145 42772
rect 3018 42692 3145 42708
rect 3018 42628 3065 42692
rect 3129 42628 3145 42692
rect 3018 42612 3145 42628
rect 3018 42548 3065 42612
rect 3129 42548 3145 42612
rect 3018 42532 3145 42548
rect 3018 42468 3065 42532
rect 3129 42468 3145 42532
rect 3018 42452 3145 42468
rect 3018 42388 3065 42452
rect 3129 42388 3145 42452
rect 3018 42372 3145 42388
rect 3018 42308 3065 42372
rect 3129 42308 3145 42372
rect 3018 42292 3145 42308
rect 3018 42228 3065 42292
rect 3129 42228 3145 42292
rect 3018 42212 3145 42228
rect 3018 42148 3065 42212
rect 3129 42148 3145 42212
rect 3018 42132 3145 42148
rect 3018 42068 3065 42132
rect 3129 42068 3145 42132
rect 3018 42052 3145 42068
rect 3018 41988 3065 42052
rect 3129 41988 3145 42052
rect 3018 41972 3145 41988
rect 3018 41908 3065 41972
rect 3129 41908 3145 41972
rect 3018 41892 3145 41908
rect 3018 41828 3065 41892
rect 3129 41828 3145 41892
rect 3018 41812 3145 41828
rect 3018 41748 3065 41812
rect 3129 41748 3145 41812
rect 3018 41732 3145 41748
rect 3018 41668 3065 41732
rect 3129 41668 3145 41732
rect 3018 41652 3145 41668
rect 3018 41588 3065 41652
rect 3129 41588 3145 41652
rect 3018 41572 3145 41588
rect 3018 41508 3065 41572
rect 3129 41508 3145 41572
rect 3018 41492 3145 41508
rect 3018 41428 3065 41492
rect 3129 41428 3145 41492
rect 3018 41412 3145 41428
rect 3018 41348 3065 41412
rect 3129 41348 3145 41412
rect 3018 41332 3145 41348
rect 3018 41268 3065 41332
rect 3129 41268 3145 41332
rect 3018 41252 3145 41268
rect 3018 41188 3065 41252
rect 3129 41188 3145 41252
rect 3018 41172 3145 41188
rect -3301 41092 -3174 41108
rect -3301 41028 -3254 41092
rect -3190 41028 -3174 41092
rect -3301 41012 -3174 41028
rect -3301 40888 -3197 41012
rect -3301 40872 -3174 40888
rect -3301 40808 -3254 40872
rect -3190 40808 -3174 40872
rect -3301 40792 -3174 40808
rect -9620 40712 -9493 40728
rect -9620 40648 -9573 40712
rect -9509 40648 -9493 40712
rect -9620 40632 -9493 40648
rect -9620 40568 -9573 40632
rect -9509 40568 -9493 40632
rect -9620 40552 -9493 40568
rect -9620 40488 -9573 40552
rect -9509 40488 -9493 40552
rect -9620 40472 -9493 40488
rect -9620 40408 -9573 40472
rect -9509 40408 -9493 40472
rect -9620 40392 -9493 40408
rect -9620 40328 -9573 40392
rect -9509 40328 -9493 40392
rect -9620 40312 -9493 40328
rect -9620 40248 -9573 40312
rect -9509 40248 -9493 40312
rect -9620 40232 -9493 40248
rect -9620 40168 -9573 40232
rect -9509 40168 -9493 40232
rect -9620 40152 -9493 40168
rect -9620 40088 -9573 40152
rect -9509 40088 -9493 40152
rect -9620 40072 -9493 40088
rect -9620 40008 -9573 40072
rect -9509 40008 -9493 40072
rect -9620 39992 -9493 40008
rect -9620 39928 -9573 39992
rect -9509 39928 -9493 39992
rect -9620 39912 -9493 39928
rect -9620 39848 -9573 39912
rect -9509 39848 -9493 39912
rect -9620 39832 -9493 39848
rect -9620 39768 -9573 39832
rect -9509 39768 -9493 39832
rect -9620 39752 -9493 39768
rect -9620 39688 -9573 39752
rect -9509 39688 -9493 39752
rect -9620 39672 -9493 39688
rect -9620 39608 -9573 39672
rect -9509 39608 -9493 39672
rect -9620 39592 -9493 39608
rect -9620 39528 -9573 39592
rect -9509 39528 -9493 39592
rect -9620 39512 -9493 39528
rect -9620 39448 -9573 39512
rect -9509 39448 -9493 39512
rect -9620 39432 -9493 39448
rect -9620 39368 -9573 39432
rect -9509 39368 -9493 39432
rect -9620 39352 -9493 39368
rect -9620 39288 -9573 39352
rect -9509 39288 -9493 39352
rect -9620 39272 -9493 39288
rect -9620 39208 -9573 39272
rect -9509 39208 -9493 39272
rect -9620 39192 -9493 39208
rect -9620 39128 -9573 39192
rect -9509 39128 -9493 39192
rect -9620 39112 -9493 39128
rect -9620 39048 -9573 39112
rect -9509 39048 -9493 39112
rect -9620 39032 -9493 39048
rect -9620 38968 -9573 39032
rect -9509 38968 -9493 39032
rect -9620 38952 -9493 38968
rect -9620 38888 -9573 38952
rect -9509 38888 -9493 38952
rect -9620 38872 -9493 38888
rect -9620 38808 -9573 38872
rect -9509 38808 -9493 38872
rect -9620 38792 -9493 38808
rect -9620 38728 -9573 38792
rect -9509 38728 -9493 38792
rect -9620 38712 -9493 38728
rect -9620 38648 -9573 38712
rect -9509 38648 -9493 38712
rect -9620 38632 -9493 38648
rect -9620 38568 -9573 38632
rect -9509 38568 -9493 38632
rect -9620 38552 -9493 38568
rect -9620 38488 -9573 38552
rect -9509 38488 -9493 38552
rect -9620 38472 -9493 38488
rect -9620 38408 -9573 38472
rect -9509 38408 -9493 38472
rect -9620 38392 -9493 38408
rect -9620 38328 -9573 38392
rect -9509 38328 -9493 38392
rect -9620 38312 -9493 38328
rect -9620 38248 -9573 38312
rect -9509 38248 -9493 38312
rect -9620 38232 -9493 38248
rect -9620 38168 -9573 38232
rect -9509 38168 -9493 38232
rect -9620 38152 -9493 38168
rect -9620 38088 -9573 38152
rect -9509 38088 -9493 38152
rect -9620 38072 -9493 38088
rect -9620 38008 -9573 38072
rect -9509 38008 -9493 38072
rect -9620 37992 -9493 38008
rect -9620 37928 -9573 37992
rect -9509 37928 -9493 37992
rect -9620 37912 -9493 37928
rect -9620 37848 -9573 37912
rect -9509 37848 -9493 37912
rect -9620 37832 -9493 37848
rect -9620 37768 -9573 37832
rect -9509 37768 -9493 37832
rect -9620 37752 -9493 37768
rect -9620 37688 -9573 37752
rect -9509 37688 -9493 37752
rect -9620 37672 -9493 37688
rect -9620 37608 -9573 37672
rect -9509 37608 -9493 37672
rect -9620 37592 -9493 37608
rect -9620 37528 -9573 37592
rect -9509 37528 -9493 37592
rect -9620 37512 -9493 37528
rect -9620 37448 -9573 37512
rect -9509 37448 -9493 37512
rect -9620 37432 -9493 37448
rect -9620 37368 -9573 37432
rect -9509 37368 -9493 37432
rect -9620 37352 -9493 37368
rect -9620 37288 -9573 37352
rect -9509 37288 -9493 37352
rect -9620 37272 -9493 37288
rect -9620 37208 -9573 37272
rect -9509 37208 -9493 37272
rect -9620 37192 -9493 37208
rect -9620 37128 -9573 37192
rect -9509 37128 -9493 37192
rect -9620 37112 -9493 37128
rect -9620 37048 -9573 37112
rect -9509 37048 -9493 37112
rect -9620 37032 -9493 37048
rect -9620 36968 -9573 37032
rect -9509 36968 -9493 37032
rect -9620 36952 -9493 36968
rect -9620 36888 -9573 36952
rect -9509 36888 -9493 36952
rect -9620 36872 -9493 36888
rect -9620 36808 -9573 36872
rect -9509 36808 -9493 36872
rect -9620 36792 -9493 36808
rect -9620 36728 -9573 36792
rect -9509 36728 -9493 36792
rect -9620 36712 -9493 36728
rect -9620 36648 -9573 36712
rect -9509 36648 -9493 36712
rect -9620 36632 -9493 36648
rect -9620 36568 -9573 36632
rect -9509 36568 -9493 36632
rect -9620 36552 -9493 36568
rect -9620 36488 -9573 36552
rect -9509 36488 -9493 36552
rect -9620 36472 -9493 36488
rect -9620 36408 -9573 36472
rect -9509 36408 -9493 36472
rect -9620 36392 -9493 36408
rect -9620 36328 -9573 36392
rect -9509 36328 -9493 36392
rect -9620 36312 -9493 36328
rect -9620 36248 -9573 36312
rect -9509 36248 -9493 36312
rect -9620 36232 -9493 36248
rect -9620 36168 -9573 36232
rect -9509 36168 -9493 36232
rect -9620 36152 -9493 36168
rect -9620 36088 -9573 36152
rect -9509 36088 -9493 36152
rect -9620 36072 -9493 36088
rect -9620 36008 -9573 36072
rect -9509 36008 -9493 36072
rect -9620 35992 -9493 36008
rect -9620 35928 -9573 35992
rect -9509 35928 -9493 35992
rect -9620 35912 -9493 35928
rect -9620 35848 -9573 35912
rect -9509 35848 -9493 35912
rect -9620 35832 -9493 35848
rect -9620 35768 -9573 35832
rect -9509 35768 -9493 35832
rect -9620 35752 -9493 35768
rect -9620 35688 -9573 35752
rect -9509 35688 -9493 35752
rect -9620 35672 -9493 35688
rect -9620 35608 -9573 35672
rect -9509 35608 -9493 35672
rect -9620 35592 -9493 35608
rect -9620 35528 -9573 35592
rect -9509 35528 -9493 35592
rect -9620 35512 -9493 35528
rect -9620 35448 -9573 35512
rect -9509 35448 -9493 35512
rect -9620 35432 -9493 35448
rect -9620 35368 -9573 35432
rect -9509 35368 -9493 35432
rect -9620 35352 -9493 35368
rect -9620 35288 -9573 35352
rect -9509 35288 -9493 35352
rect -9620 35272 -9493 35288
rect -9620 35208 -9573 35272
rect -9509 35208 -9493 35272
rect -9620 35192 -9493 35208
rect -9620 35128 -9573 35192
rect -9509 35128 -9493 35192
rect -9620 35112 -9493 35128
rect -9620 35048 -9573 35112
rect -9509 35048 -9493 35112
rect -9620 35032 -9493 35048
rect -9620 34968 -9573 35032
rect -9509 34968 -9493 35032
rect -9620 34952 -9493 34968
rect -9620 34888 -9573 34952
rect -9509 34888 -9493 34952
rect -9620 34872 -9493 34888
rect -15939 34792 -15812 34808
rect -15939 34728 -15892 34792
rect -15828 34728 -15812 34792
rect -15939 34712 -15812 34728
rect -15939 34588 -15835 34712
rect -15939 34572 -15812 34588
rect -15939 34508 -15892 34572
rect -15828 34508 -15812 34572
rect -15939 34492 -15812 34508
rect -22258 34412 -22131 34428
rect -22258 34348 -22211 34412
rect -22147 34348 -22131 34412
rect -22258 34332 -22131 34348
rect -22258 34268 -22211 34332
rect -22147 34268 -22131 34332
rect -22258 34252 -22131 34268
rect -22258 34188 -22211 34252
rect -22147 34188 -22131 34252
rect -22258 34172 -22131 34188
rect -22258 34108 -22211 34172
rect -22147 34108 -22131 34172
rect -22258 34092 -22131 34108
rect -22258 34028 -22211 34092
rect -22147 34028 -22131 34092
rect -22258 34012 -22131 34028
rect -22258 33948 -22211 34012
rect -22147 33948 -22131 34012
rect -22258 33932 -22131 33948
rect -22258 33868 -22211 33932
rect -22147 33868 -22131 33932
rect -22258 33852 -22131 33868
rect -22258 33788 -22211 33852
rect -22147 33788 -22131 33852
rect -22258 33772 -22131 33788
rect -22258 33708 -22211 33772
rect -22147 33708 -22131 33772
rect -22258 33692 -22131 33708
rect -22258 33628 -22211 33692
rect -22147 33628 -22131 33692
rect -22258 33612 -22131 33628
rect -22258 33548 -22211 33612
rect -22147 33548 -22131 33612
rect -22258 33532 -22131 33548
rect -22258 33468 -22211 33532
rect -22147 33468 -22131 33532
rect -22258 33452 -22131 33468
rect -22258 33388 -22211 33452
rect -22147 33388 -22131 33452
rect -22258 33372 -22131 33388
rect -22258 33308 -22211 33372
rect -22147 33308 -22131 33372
rect -22258 33292 -22131 33308
rect -22258 33228 -22211 33292
rect -22147 33228 -22131 33292
rect -22258 33212 -22131 33228
rect -22258 33148 -22211 33212
rect -22147 33148 -22131 33212
rect -22258 33132 -22131 33148
rect -22258 33068 -22211 33132
rect -22147 33068 -22131 33132
rect -22258 33052 -22131 33068
rect -22258 32988 -22211 33052
rect -22147 32988 -22131 33052
rect -22258 32972 -22131 32988
rect -22258 32908 -22211 32972
rect -22147 32908 -22131 32972
rect -22258 32892 -22131 32908
rect -22258 32828 -22211 32892
rect -22147 32828 -22131 32892
rect -22258 32812 -22131 32828
rect -22258 32748 -22211 32812
rect -22147 32748 -22131 32812
rect -22258 32732 -22131 32748
rect -22258 32668 -22211 32732
rect -22147 32668 -22131 32732
rect -22258 32652 -22131 32668
rect -22258 32588 -22211 32652
rect -22147 32588 -22131 32652
rect -22258 32572 -22131 32588
rect -22258 32508 -22211 32572
rect -22147 32508 -22131 32572
rect -22258 32492 -22131 32508
rect -22258 32428 -22211 32492
rect -22147 32428 -22131 32492
rect -22258 32412 -22131 32428
rect -22258 32348 -22211 32412
rect -22147 32348 -22131 32412
rect -22258 32332 -22131 32348
rect -22258 32268 -22211 32332
rect -22147 32268 -22131 32332
rect -22258 32252 -22131 32268
rect -22258 32188 -22211 32252
rect -22147 32188 -22131 32252
rect -22258 32172 -22131 32188
rect -22258 32108 -22211 32172
rect -22147 32108 -22131 32172
rect -22258 32092 -22131 32108
rect -22258 32028 -22211 32092
rect -22147 32028 -22131 32092
rect -22258 32012 -22131 32028
rect -22258 31948 -22211 32012
rect -22147 31948 -22131 32012
rect -22258 31932 -22131 31948
rect -22258 31868 -22211 31932
rect -22147 31868 -22131 31932
rect -22258 31852 -22131 31868
rect -22258 31788 -22211 31852
rect -22147 31788 -22131 31852
rect -22258 31772 -22131 31788
rect -22258 31708 -22211 31772
rect -22147 31708 -22131 31772
rect -22258 31692 -22131 31708
rect -22258 31628 -22211 31692
rect -22147 31628 -22131 31692
rect -22258 31612 -22131 31628
rect -22258 31548 -22211 31612
rect -22147 31548 -22131 31612
rect -22258 31532 -22131 31548
rect -22258 31468 -22211 31532
rect -22147 31468 -22131 31532
rect -22258 31452 -22131 31468
rect -22258 31388 -22211 31452
rect -22147 31388 -22131 31452
rect -22258 31372 -22131 31388
rect -22258 31308 -22211 31372
rect -22147 31308 -22131 31372
rect -22258 31292 -22131 31308
rect -22258 31228 -22211 31292
rect -22147 31228 -22131 31292
rect -22258 31212 -22131 31228
rect -22258 31148 -22211 31212
rect -22147 31148 -22131 31212
rect -22258 31132 -22131 31148
rect -22258 31068 -22211 31132
rect -22147 31068 -22131 31132
rect -22258 31052 -22131 31068
rect -22258 30988 -22211 31052
rect -22147 30988 -22131 31052
rect -22258 30972 -22131 30988
rect -22258 30908 -22211 30972
rect -22147 30908 -22131 30972
rect -22258 30892 -22131 30908
rect -22258 30828 -22211 30892
rect -22147 30828 -22131 30892
rect -22258 30812 -22131 30828
rect -22258 30748 -22211 30812
rect -22147 30748 -22131 30812
rect -22258 30732 -22131 30748
rect -22258 30668 -22211 30732
rect -22147 30668 -22131 30732
rect -22258 30652 -22131 30668
rect -22258 30588 -22211 30652
rect -22147 30588 -22131 30652
rect -22258 30572 -22131 30588
rect -22258 30508 -22211 30572
rect -22147 30508 -22131 30572
rect -22258 30492 -22131 30508
rect -22258 30428 -22211 30492
rect -22147 30428 -22131 30492
rect -22258 30412 -22131 30428
rect -22258 30348 -22211 30412
rect -22147 30348 -22131 30412
rect -22258 30332 -22131 30348
rect -22258 30268 -22211 30332
rect -22147 30268 -22131 30332
rect -22258 30252 -22131 30268
rect -22258 30188 -22211 30252
rect -22147 30188 -22131 30252
rect -22258 30172 -22131 30188
rect -22258 30108 -22211 30172
rect -22147 30108 -22131 30172
rect -22258 30092 -22131 30108
rect -22258 30028 -22211 30092
rect -22147 30028 -22131 30092
rect -22258 30012 -22131 30028
rect -22258 29948 -22211 30012
rect -22147 29948 -22131 30012
rect -22258 29932 -22131 29948
rect -22258 29868 -22211 29932
rect -22147 29868 -22131 29932
rect -22258 29852 -22131 29868
rect -22258 29788 -22211 29852
rect -22147 29788 -22131 29852
rect -22258 29772 -22131 29788
rect -22258 29708 -22211 29772
rect -22147 29708 -22131 29772
rect -22258 29692 -22131 29708
rect -22258 29628 -22211 29692
rect -22147 29628 -22131 29692
rect -22258 29612 -22131 29628
rect -22258 29548 -22211 29612
rect -22147 29548 -22131 29612
rect -22258 29532 -22131 29548
rect -22258 29468 -22211 29532
rect -22147 29468 -22131 29532
rect -22258 29452 -22131 29468
rect -22258 29388 -22211 29452
rect -22147 29388 -22131 29452
rect -22258 29372 -22131 29388
rect -22258 29308 -22211 29372
rect -22147 29308 -22131 29372
rect -22258 29292 -22131 29308
rect -22258 29228 -22211 29292
rect -22147 29228 -22131 29292
rect -22258 29212 -22131 29228
rect -22258 29148 -22211 29212
rect -22147 29148 -22131 29212
rect -22258 29132 -22131 29148
rect -22258 29068 -22211 29132
rect -22147 29068 -22131 29132
rect -22258 29052 -22131 29068
rect -22258 28988 -22211 29052
rect -22147 28988 -22131 29052
rect -22258 28972 -22131 28988
rect -22258 28908 -22211 28972
rect -22147 28908 -22131 28972
rect -22258 28892 -22131 28908
rect -22258 28828 -22211 28892
rect -22147 28828 -22131 28892
rect -22258 28812 -22131 28828
rect -22258 28748 -22211 28812
rect -22147 28748 -22131 28812
rect -22258 28732 -22131 28748
rect -22258 28668 -22211 28732
rect -22147 28668 -22131 28732
rect -22258 28652 -22131 28668
rect -22258 28588 -22211 28652
rect -22147 28588 -22131 28652
rect -22258 28572 -22131 28588
rect -28577 28492 -28450 28508
rect -28577 28428 -28530 28492
rect -28466 28428 -28450 28492
rect -28577 28412 -28450 28428
rect -28577 28288 -28473 28412
rect -28577 28272 -28450 28288
rect -28577 28208 -28530 28272
rect -28466 28208 -28450 28272
rect -28577 28192 -28450 28208
rect -34896 28112 -34769 28128
rect -34896 28048 -34849 28112
rect -34785 28048 -34769 28112
rect -34896 28032 -34769 28048
rect -34896 27968 -34849 28032
rect -34785 27968 -34769 28032
rect -34896 27952 -34769 27968
rect -34896 27888 -34849 27952
rect -34785 27888 -34769 27952
rect -34896 27872 -34769 27888
rect -34896 27808 -34849 27872
rect -34785 27808 -34769 27872
rect -34896 27792 -34769 27808
rect -34896 27728 -34849 27792
rect -34785 27728 -34769 27792
rect -34896 27712 -34769 27728
rect -34896 27648 -34849 27712
rect -34785 27648 -34769 27712
rect -34896 27632 -34769 27648
rect -34896 27568 -34849 27632
rect -34785 27568 -34769 27632
rect -34896 27552 -34769 27568
rect -34896 27488 -34849 27552
rect -34785 27488 -34769 27552
rect -34896 27472 -34769 27488
rect -34896 27408 -34849 27472
rect -34785 27408 -34769 27472
rect -34896 27392 -34769 27408
rect -34896 27328 -34849 27392
rect -34785 27328 -34769 27392
rect -34896 27312 -34769 27328
rect -34896 27248 -34849 27312
rect -34785 27248 -34769 27312
rect -34896 27232 -34769 27248
rect -34896 27168 -34849 27232
rect -34785 27168 -34769 27232
rect -34896 27152 -34769 27168
rect -34896 27088 -34849 27152
rect -34785 27088 -34769 27152
rect -34896 27072 -34769 27088
rect -34896 27008 -34849 27072
rect -34785 27008 -34769 27072
rect -34896 26992 -34769 27008
rect -34896 26928 -34849 26992
rect -34785 26928 -34769 26992
rect -34896 26912 -34769 26928
rect -34896 26848 -34849 26912
rect -34785 26848 -34769 26912
rect -34896 26832 -34769 26848
rect -34896 26768 -34849 26832
rect -34785 26768 -34769 26832
rect -34896 26752 -34769 26768
rect -34896 26688 -34849 26752
rect -34785 26688 -34769 26752
rect -34896 26672 -34769 26688
rect -34896 26608 -34849 26672
rect -34785 26608 -34769 26672
rect -34896 26592 -34769 26608
rect -34896 26528 -34849 26592
rect -34785 26528 -34769 26592
rect -34896 26512 -34769 26528
rect -34896 26448 -34849 26512
rect -34785 26448 -34769 26512
rect -34896 26432 -34769 26448
rect -34896 26368 -34849 26432
rect -34785 26368 -34769 26432
rect -34896 26352 -34769 26368
rect -34896 26288 -34849 26352
rect -34785 26288 -34769 26352
rect -34896 26272 -34769 26288
rect -34896 26208 -34849 26272
rect -34785 26208 -34769 26272
rect -34896 26192 -34769 26208
rect -34896 26128 -34849 26192
rect -34785 26128 -34769 26192
rect -34896 26112 -34769 26128
rect -34896 26048 -34849 26112
rect -34785 26048 -34769 26112
rect -34896 26032 -34769 26048
rect -34896 25968 -34849 26032
rect -34785 25968 -34769 26032
rect -34896 25952 -34769 25968
rect -34896 25888 -34849 25952
rect -34785 25888 -34769 25952
rect -34896 25872 -34769 25888
rect -34896 25808 -34849 25872
rect -34785 25808 -34769 25872
rect -34896 25792 -34769 25808
rect -34896 25728 -34849 25792
rect -34785 25728 -34769 25792
rect -34896 25712 -34769 25728
rect -34896 25648 -34849 25712
rect -34785 25648 -34769 25712
rect -34896 25632 -34769 25648
rect -34896 25568 -34849 25632
rect -34785 25568 -34769 25632
rect -34896 25552 -34769 25568
rect -34896 25488 -34849 25552
rect -34785 25488 -34769 25552
rect -34896 25472 -34769 25488
rect -34896 25408 -34849 25472
rect -34785 25408 -34769 25472
rect -34896 25392 -34769 25408
rect -34896 25328 -34849 25392
rect -34785 25328 -34769 25392
rect -34896 25312 -34769 25328
rect -34896 25248 -34849 25312
rect -34785 25248 -34769 25312
rect -34896 25232 -34769 25248
rect -34896 25168 -34849 25232
rect -34785 25168 -34769 25232
rect -34896 25152 -34769 25168
rect -34896 25088 -34849 25152
rect -34785 25088 -34769 25152
rect -34896 25072 -34769 25088
rect -34896 25008 -34849 25072
rect -34785 25008 -34769 25072
rect -34896 24992 -34769 25008
rect -34896 24928 -34849 24992
rect -34785 24928 -34769 24992
rect -34896 24912 -34769 24928
rect -34896 24848 -34849 24912
rect -34785 24848 -34769 24912
rect -34896 24832 -34769 24848
rect -34896 24768 -34849 24832
rect -34785 24768 -34769 24832
rect -34896 24752 -34769 24768
rect -34896 24688 -34849 24752
rect -34785 24688 -34769 24752
rect -34896 24672 -34769 24688
rect -34896 24608 -34849 24672
rect -34785 24608 -34769 24672
rect -34896 24592 -34769 24608
rect -34896 24528 -34849 24592
rect -34785 24528 -34769 24592
rect -34896 24512 -34769 24528
rect -34896 24448 -34849 24512
rect -34785 24448 -34769 24512
rect -34896 24432 -34769 24448
rect -34896 24368 -34849 24432
rect -34785 24368 -34769 24432
rect -34896 24352 -34769 24368
rect -34896 24288 -34849 24352
rect -34785 24288 -34769 24352
rect -34896 24272 -34769 24288
rect -34896 24208 -34849 24272
rect -34785 24208 -34769 24272
rect -34896 24192 -34769 24208
rect -34896 24128 -34849 24192
rect -34785 24128 -34769 24192
rect -34896 24112 -34769 24128
rect -34896 24048 -34849 24112
rect -34785 24048 -34769 24112
rect -34896 24032 -34769 24048
rect -34896 23968 -34849 24032
rect -34785 23968 -34769 24032
rect -34896 23952 -34769 23968
rect -34896 23888 -34849 23952
rect -34785 23888 -34769 23952
rect -34896 23872 -34769 23888
rect -34896 23808 -34849 23872
rect -34785 23808 -34769 23872
rect -34896 23792 -34769 23808
rect -34896 23728 -34849 23792
rect -34785 23728 -34769 23792
rect -34896 23712 -34769 23728
rect -34896 23648 -34849 23712
rect -34785 23648 -34769 23712
rect -34896 23632 -34769 23648
rect -34896 23568 -34849 23632
rect -34785 23568 -34769 23632
rect -34896 23552 -34769 23568
rect -34896 23488 -34849 23552
rect -34785 23488 -34769 23552
rect -34896 23472 -34769 23488
rect -34896 23408 -34849 23472
rect -34785 23408 -34769 23472
rect -34896 23392 -34769 23408
rect -34896 23328 -34849 23392
rect -34785 23328 -34769 23392
rect -34896 23312 -34769 23328
rect -34896 23248 -34849 23312
rect -34785 23248 -34769 23312
rect -34896 23232 -34769 23248
rect -34896 23168 -34849 23232
rect -34785 23168 -34769 23232
rect -34896 23152 -34769 23168
rect -34896 23088 -34849 23152
rect -34785 23088 -34769 23152
rect -34896 23072 -34769 23088
rect -34896 23008 -34849 23072
rect -34785 23008 -34769 23072
rect -34896 22992 -34769 23008
rect -34896 22928 -34849 22992
rect -34785 22928 -34769 22992
rect -34896 22912 -34769 22928
rect -34896 22848 -34849 22912
rect -34785 22848 -34769 22912
rect -34896 22832 -34769 22848
rect -34896 22768 -34849 22832
rect -34785 22768 -34769 22832
rect -34896 22752 -34769 22768
rect -34896 22688 -34849 22752
rect -34785 22688 -34769 22752
rect -34896 22672 -34769 22688
rect -34896 22608 -34849 22672
rect -34785 22608 -34769 22672
rect -34896 22592 -34769 22608
rect -34896 22528 -34849 22592
rect -34785 22528 -34769 22592
rect -34896 22512 -34769 22528
rect -34896 22448 -34849 22512
rect -34785 22448 -34769 22512
rect -34896 22432 -34769 22448
rect -34896 22368 -34849 22432
rect -34785 22368 -34769 22432
rect -34896 22352 -34769 22368
rect -34896 22288 -34849 22352
rect -34785 22288 -34769 22352
rect -34896 22272 -34769 22288
rect -41215 22192 -41088 22208
rect -41215 22128 -41168 22192
rect -41104 22128 -41088 22192
rect -41215 22112 -41088 22128
rect -41215 21988 -41111 22112
rect -41215 21972 -41088 21988
rect -41215 21908 -41168 21972
rect -41104 21908 -41088 21972
rect -41215 21892 -41088 21908
rect -47244 21852 -41322 21861
rect -47244 15948 -47235 21852
rect -41331 15948 -41322 21852
rect -47244 15939 -41322 15948
rect -41215 21828 -41168 21892
rect -41104 21828 -41088 21892
rect -38016 21861 -37912 22239
rect -34896 22208 -34849 22272
rect -34785 22208 -34769 22272
rect -34606 28152 -28684 28161
rect -34606 22248 -34597 28152
rect -28693 22248 -28684 28152
rect -34606 22239 -28684 22248
rect -28577 28128 -28530 28192
rect -28466 28128 -28450 28192
rect -25378 28161 -25274 28539
rect -22258 28508 -22211 28572
rect -22147 28508 -22131 28572
rect -21968 34452 -16046 34461
rect -21968 28548 -21959 34452
rect -16055 28548 -16046 34452
rect -21968 28539 -16046 28548
rect -15939 34428 -15892 34492
rect -15828 34428 -15812 34492
rect -12740 34461 -12636 34839
rect -9620 34808 -9573 34872
rect -9509 34808 -9493 34872
rect -9330 40752 -3408 40761
rect -9330 34848 -9321 40752
rect -3417 34848 -3408 40752
rect -9330 34839 -3408 34848
rect -3301 40728 -3254 40792
rect -3190 40728 -3174 40792
rect -102 40761 2 41139
rect 3018 41108 3065 41172
rect 3129 41108 3145 41172
rect 3308 47052 9230 47061
rect 3308 41148 3317 47052
rect 9221 41148 9230 47052
rect 3308 41139 9230 41148
rect 9337 47028 9384 47092
rect 9448 47028 9464 47092
rect 12536 47061 12640 47250
rect 15656 47188 15760 47250
rect 15656 47172 15783 47188
rect 15656 47108 15703 47172
rect 15767 47108 15783 47172
rect 15656 47092 15783 47108
rect 9337 47012 9464 47028
rect 9337 46948 9384 47012
rect 9448 46948 9464 47012
rect 9337 46932 9464 46948
rect 9337 46868 9384 46932
rect 9448 46868 9464 46932
rect 9337 46852 9464 46868
rect 9337 46788 9384 46852
rect 9448 46788 9464 46852
rect 9337 46772 9464 46788
rect 9337 46708 9384 46772
rect 9448 46708 9464 46772
rect 9337 46692 9464 46708
rect 9337 46628 9384 46692
rect 9448 46628 9464 46692
rect 9337 46612 9464 46628
rect 9337 46548 9384 46612
rect 9448 46548 9464 46612
rect 9337 46532 9464 46548
rect 9337 46468 9384 46532
rect 9448 46468 9464 46532
rect 9337 46452 9464 46468
rect 9337 46388 9384 46452
rect 9448 46388 9464 46452
rect 9337 46372 9464 46388
rect 9337 46308 9384 46372
rect 9448 46308 9464 46372
rect 9337 46292 9464 46308
rect 9337 46228 9384 46292
rect 9448 46228 9464 46292
rect 9337 46212 9464 46228
rect 9337 46148 9384 46212
rect 9448 46148 9464 46212
rect 9337 46132 9464 46148
rect 9337 46068 9384 46132
rect 9448 46068 9464 46132
rect 9337 46052 9464 46068
rect 9337 45988 9384 46052
rect 9448 45988 9464 46052
rect 9337 45972 9464 45988
rect 9337 45908 9384 45972
rect 9448 45908 9464 45972
rect 9337 45892 9464 45908
rect 9337 45828 9384 45892
rect 9448 45828 9464 45892
rect 9337 45812 9464 45828
rect 9337 45748 9384 45812
rect 9448 45748 9464 45812
rect 9337 45732 9464 45748
rect 9337 45668 9384 45732
rect 9448 45668 9464 45732
rect 9337 45652 9464 45668
rect 9337 45588 9384 45652
rect 9448 45588 9464 45652
rect 9337 45572 9464 45588
rect 9337 45508 9384 45572
rect 9448 45508 9464 45572
rect 9337 45492 9464 45508
rect 9337 45428 9384 45492
rect 9448 45428 9464 45492
rect 9337 45412 9464 45428
rect 9337 45348 9384 45412
rect 9448 45348 9464 45412
rect 9337 45332 9464 45348
rect 9337 45268 9384 45332
rect 9448 45268 9464 45332
rect 9337 45252 9464 45268
rect 9337 45188 9384 45252
rect 9448 45188 9464 45252
rect 9337 45172 9464 45188
rect 9337 45108 9384 45172
rect 9448 45108 9464 45172
rect 9337 45092 9464 45108
rect 9337 45028 9384 45092
rect 9448 45028 9464 45092
rect 9337 45012 9464 45028
rect 9337 44948 9384 45012
rect 9448 44948 9464 45012
rect 9337 44932 9464 44948
rect 9337 44868 9384 44932
rect 9448 44868 9464 44932
rect 9337 44852 9464 44868
rect 9337 44788 9384 44852
rect 9448 44788 9464 44852
rect 9337 44772 9464 44788
rect 9337 44708 9384 44772
rect 9448 44708 9464 44772
rect 9337 44692 9464 44708
rect 9337 44628 9384 44692
rect 9448 44628 9464 44692
rect 9337 44612 9464 44628
rect 9337 44548 9384 44612
rect 9448 44548 9464 44612
rect 9337 44532 9464 44548
rect 9337 44468 9384 44532
rect 9448 44468 9464 44532
rect 9337 44452 9464 44468
rect 9337 44388 9384 44452
rect 9448 44388 9464 44452
rect 9337 44372 9464 44388
rect 9337 44308 9384 44372
rect 9448 44308 9464 44372
rect 9337 44292 9464 44308
rect 9337 44228 9384 44292
rect 9448 44228 9464 44292
rect 9337 44212 9464 44228
rect 9337 44148 9384 44212
rect 9448 44148 9464 44212
rect 9337 44132 9464 44148
rect 9337 44068 9384 44132
rect 9448 44068 9464 44132
rect 9337 44052 9464 44068
rect 9337 43988 9384 44052
rect 9448 43988 9464 44052
rect 9337 43972 9464 43988
rect 9337 43908 9384 43972
rect 9448 43908 9464 43972
rect 9337 43892 9464 43908
rect 9337 43828 9384 43892
rect 9448 43828 9464 43892
rect 9337 43812 9464 43828
rect 9337 43748 9384 43812
rect 9448 43748 9464 43812
rect 9337 43732 9464 43748
rect 9337 43668 9384 43732
rect 9448 43668 9464 43732
rect 9337 43652 9464 43668
rect 9337 43588 9384 43652
rect 9448 43588 9464 43652
rect 9337 43572 9464 43588
rect 9337 43508 9384 43572
rect 9448 43508 9464 43572
rect 9337 43492 9464 43508
rect 9337 43428 9384 43492
rect 9448 43428 9464 43492
rect 9337 43412 9464 43428
rect 9337 43348 9384 43412
rect 9448 43348 9464 43412
rect 9337 43332 9464 43348
rect 9337 43268 9384 43332
rect 9448 43268 9464 43332
rect 9337 43252 9464 43268
rect 9337 43188 9384 43252
rect 9448 43188 9464 43252
rect 9337 43172 9464 43188
rect 9337 43108 9384 43172
rect 9448 43108 9464 43172
rect 9337 43092 9464 43108
rect 9337 43028 9384 43092
rect 9448 43028 9464 43092
rect 9337 43012 9464 43028
rect 9337 42948 9384 43012
rect 9448 42948 9464 43012
rect 9337 42932 9464 42948
rect 9337 42868 9384 42932
rect 9448 42868 9464 42932
rect 9337 42852 9464 42868
rect 9337 42788 9384 42852
rect 9448 42788 9464 42852
rect 9337 42772 9464 42788
rect 9337 42708 9384 42772
rect 9448 42708 9464 42772
rect 9337 42692 9464 42708
rect 9337 42628 9384 42692
rect 9448 42628 9464 42692
rect 9337 42612 9464 42628
rect 9337 42548 9384 42612
rect 9448 42548 9464 42612
rect 9337 42532 9464 42548
rect 9337 42468 9384 42532
rect 9448 42468 9464 42532
rect 9337 42452 9464 42468
rect 9337 42388 9384 42452
rect 9448 42388 9464 42452
rect 9337 42372 9464 42388
rect 9337 42308 9384 42372
rect 9448 42308 9464 42372
rect 9337 42292 9464 42308
rect 9337 42228 9384 42292
rect 9448 42228 9464 42292
rect 9337 42212 9464 42228
rect 9337 42148 9384 42212
rect 9448 42148 9464 42212
rect 9337 42132 9464 42148
rect 9337 42068 9384 42132
rect 9448 42068 9464 42132
rect 9337 42052 9464 42068
rect 9337 41988 9384 42052
rect 9448 41988 9464 42052
rect 9337 41972 9464 41988
rect 9337 41908 9384 41972
rect 9448 41908 9464 41972
rect 9337 41892 9464 41908
rect 9337 41828 9384 41892
rect 9448 41828 9464 41892
rect 9337 41812 9464 41828
rect 9337 41748 9384 41812
rect 9448 41748 9464 41812
rect 9337 41732 9464 41748
rect 9337 41668 9384 41732
rect 9448 41668 9464 41732
rect 9337 41652 9464 41668
rect 9337 41588 9384 41652
rect 9448 41588 9464 41652
rect 9337 41572 9464 41588
rect 9337 41508 9384 41572
rect 9448 41508 9464 41572
rect 9337 41492 9464 41508
rect 9337 41428 9384 41492
rect 9448 41428 9464 41492
rect 9337 41412 9464 41428
rect 9337 41348 9384 41412
rect 9448 41348 9464 41412
rect 9337 41332 9464 41348
rect 9337 41268 9384 41332
rect 9448 41268 9464 41332
rect 9337 41252 9464 41268
rect 9337 41188 9384 41252
rect 9448 41188 9464 41252
rect 9337 41172 9464 41188
rect 3018 41092 3145 41108
rect 3018 41028 3065 41092
rect 3129 41028 3145 41092
rect 3018 41012 3145 41028
rect 3018 40888 3122 41012
rect 3018 40872 3145 40888
rect 3018 40808 3065 40872
rect 3129 40808 3145 40872
rect 3018 40792 3145 40808
rect -3301 40712 -3174 40728
rect -3301 40648 -3254 40712
rect -3190 40648 -3174 40712
rect -3301 40632 -3174 40648
rect -3301 40568 -3254 40632
rect -3190 40568 -3174 40632
rect -3301 40552 -3174 40568
rect -3301 40488 -3254 40552
rect -3190 40488 -3174 40552
rect -3301 40472 -3174 40488
rect -3301 40408 -3254 40472
rect -3190 40408 -3174 40472
rect -3301 40392 -3174 40408
rect -3301 40328 -3254 40392
rect -3190 40328 -3174 40392
rect -3301 40312 -3174 40328
rect -3301 40248 -3254 40312
rect -3190 40248 -3174 40312
rect -3301 40232 -3174 40248
rect -3301 40168 -3254 40232
rect -3190 40168 -3174 40232
rect -3301 40152 -3174 40168
rect -3301 40088 -3254 40152
rect -3190 40088 -3174 40152
rect -3301 40072 -3174 40088
rect -3301 40008 -3254 40072
rect -3190 40008 -3174 40072
rect -3301 39992 -3174 40008
rect -3301 39928 -3254 39992
rect -3190 39928 -3174 39992
rect -3301 39912 -3174 39928
rect -3301 39848 -3254 39912
rect -3190 39848 -3174 39912
rect -3301 39832 -3174 39848
rect -3301 39768 -3254 39832
rect -3190 39768 -3174 39832
rect -3301 39752 -3174 39768
rect -3301 39688 -3254 39752
rect -3190 39688 -3174 39752
rect -3301 39672 -3174 39688
rect -3301 39608 -3254 39672
rect -3190 39608 -3174 39672
rect -3301 39592 -3174 39608
rect -3301 39528 -3254 39592
rect -3190 39528 -3174 39592
rect -3301 39512 -3174 39528
rect -3301 39448 -3254 39512
rect -3190 39448 -3174 39512
rect -3301 39432 -3174 39448
rect -3301 39368 -3254 39432
rect -3190 39368 -3174 39432
rect -3301 39352 -3174 39368
rect -3301 39288 -3254 39352
rect -3190 39288 -3174 39352
rect -3301 39272 -3174 39288
rect -3301 39208 -3254 39272
rect -3190 39208 -3174 39272
rect -3301 39192 -3174 39208
rect -3301 39128 -3254 39192
rect -3190 39128 -3174 39192
rect -3301 39112 -3174 39128
rect -3301 39048 -3254 39112
rect -3190 39048 -3174 39112
rect -3301 39032 -3174 39048
rect -3301 38968 -3254 39032
rect -3190 38968 -3174 39032
rect -3301 38952 -3174 38968
rect -3301 38888 -3254 38952
rect -3190 38888 -3174 38952
rect -3301 38872 -3174 38888
rect -3301 38808 -3254 38872
rect -3190 38808 -3174 38872
rect -3301 38792 -3174 38808
rect -3301 38728 -3254 38792
rect -3190 38728 -3174 38792
rect -3301 38712 -3174 38728
rect -3301 38648 -3254 38712
rect -3190 38648 -3174 38712
rect -3301 38632 -3174 38648
rect -3301 38568 -3254 38632
rect -3190 38568 -3174 38632
rect -3301 38552 -3174 38568
rect -3301 38488 -3254 38552
rect -3190 38488 -3174 38552
rect -3301 38472 -3174 38488
rect -3301 38408 -3254 38472
rect -3190 38408 -3174 38472
rect -3301 38392 -3174 38408
rect -3301 38328 -3254 38392
rect -3190 38328 -3174 38392
rect -3301 38312 -3174 38328
rect -3301 38248 -3254 38312
rect -3190 38248 -3174 38312
rect -3301 38232 -3174 38248
rect -3301 38168 -3254 38232
rect -3190 38168 -3174 38232
rect -3301 38152 -3174 38168
rect -3301 38088 -3254 38152
rect -3190 38088 -3174 38152
rect -3301 38072 -3174 38088
rect -3301 38008 -3254 38072
rect -3190 38008 -3174 38072
rect -3301 37992 -3174 38008
rect -3301 37928 -3254 37992
rect -3190 37928 -3174 37992
rect -3301 37912 -3174 37928
rect -3301 37848 -3254 37912
rect -3190 37848 -3174 37912
rect -3301 37832 -3174 37848
rect -3301 37768 -3254 37832
rect -3190 37768 -3174 37832
rect -3301 37752 -3174 37768
rect -3301 37688 -3254 37752
rect -3190 37688 -3174 37752
rect -3301 37672 -3174 37688
rect -3301 37608 -3254 37672
rect -3190 37608 -3174 37672
rect -3301 37592 -3174 37608
rect -3301 37528 -3254 37592
rect -3190 37528 -3174 37592
rect -3301 37512 -3174 37528
rect -3301 37448 -3254 37512
rect -3190 37448 -3174 37512
rect -3301 37432 -3174 37448
rect -3301 37368 -3254 37432
rect -3190 37368 -3174 37432
rect -3301 37352 -3174 37368
rect -3301 37288 -3254 37352
rect -3190 37288 -3174 37352
rect -3301 37272 -3174 37288
rect -3301 37208 -3254 37272
rect -3190 37208 -3174 37272
rect -3301 37192 -3174 37208
rect -3301 37128 -3254 37192
rect -3190 37128 -3174 37192
rect -3301 37112 -3174 37128
rect -3301 37048 -3254 37112
rect -3190 37048 -3174 37112
rect -3301 37032 -3174 37048
rect -3301 36968 -3254 37032
rect -3190 36968 -3174 37032
rect -3301 36952 -3174 36968
rect -3301 36888 -3254 36952
rect -3190 36888 -3174 36952
rect -3301 36872 -3174 36888
rect -3301 36808 -3254 36872
rect -3190 36808 -3174 36872
rect -3301 36792 -3174 36808
rect -3301 36728 -3254 36792
rect -3190 36728 -3174 36792
rect -3301 36712 -3174 36728
rect -3301 36648 -3254 36712
rect -3190 36648 -3174 36712
rect -3301 36632 -3174 36648
rect -3301 36568 -3254 36632
rect -3190 36568 -3174 36632
rect -3301 36552 -3174 36568
rect -3301 36488 -3254 36552
rect -3190 36488 -3174 36552
rect -3301 36472 -3174 36488
rect -3301 36408 -3254 36472
rect -3190 36408 -3174 36472
rect -3301 36392 -3174 36408
rect -3301 36328 -3254 36392
rect -3190 36328 -3174 36392
rect -3301 36312 -3174 36328
rect -3301 36248 -3254 36312
rect -3190 36248 -3174 36312
rect -3301 36232 -3174 36248
rect -3301 36168 -3254 36232
rect -3190 36168 -3174 36232
rect -3301 36152 -3174 36168
rect -3301 36088 -3254 36152
rect -3190 36088 -3174 36152
rect -3301 36072 -3174 36088
rect -3301 36008 -3254 36072
rect -3190 36008 -3174 36072
rect -3301 35992 -3174 36008
rect -3301 35928 -3254 35992
rect -3190 35928 -3174 35992
rect -3301 35912 -3174 35928
rect -3301 35848 -3254 35912
rect -3190 35848 -3174 35912
rect -3301 35832 -3174 35848
rect -3301 35768 -3254 35832
rect -3190 35768 -3174 35832
rect -3301 35752 -3174 35768
rect -3301 35688 -3254 35752
rect -3190 35688 -3174 35752
rect -3301 35672 -3174 35688
rect -3301 35608 -3254 35672
rect -3190 35608 -3174 35672
rect -3301 35592 -3174 35608
rect -3301 35528 -3254 35592
rect -3190 35528 -3174 35592
rect -3301 35512 -3174 35528
rect -3301 35448 -3254 35512
rect -3190 35448 -3174 35512
rect -3301 35432 -3174 35448
rect -3301 35368 -3254 35432
rect -3190 35368 -3174 35432
rect -3301 35352 -3174 35368
rect -3301 35288 -3254 35352
rect -3190 35288 -3174 35352
rect -3301 35272 -3174 35288
rect -3301 35208 -3254 35272
rect -3190 35208 -3174 35272
rect -3301 35192 -3174 35208
rect -3301 35128 -3254 35192
rect -3190 35128 -3174 35192
rect -3301 35112 -3174 35128
rect -3301 35048 -3254 35112
rect -3190 35048 -3174 35112
rect -3301 35032 -3174 35048
rect -3301 34968 -3254 35032
rect -3190 34968 -3174 35032
rect -3301 34952 -3174 34968
rect -3301 34888 -3254 34952
rect -3190 34888 -3174 34952
rect -3301 34872 -3174 34888
rect -9620 34792 -9493 34808
rect -9620 34728 -9573 34792
rect -9509 34728 -9493 34792
rect -9620 34712 -9493 34728
rect -9620 34588 -9516 34712
rect -9620 34572 -9493 34588
rect -9620 34508 -9573 34572
rect -9509 34508 -9493 34572
rect -9620 34492 -9493 34508
rect -15939 34412 -15812 34428
rect -15939 34348 -15892 34412
rect -15828 34348 -15812 34412
rect -15939 34332 -15812 34348
rect -15939 34268 -15892 34332
rect -15828 34268 -15812 34332
rect -15939 34252 -15812 34268
rect -15939 34188 -15892 34252
rect -15828 34188 -15812 34252
rect -15939 34172 -15812 34188
rect -15939 34108 -15892 34172
rect -15828 34108 -15812 34172
rect -15939 34092 -15812 34108
rect -15939 34028 -15892 34092
rect -15828 34028 -15812 34092
rect -15939 34012 -15812 34028
rect -15939 33948 -15892 34012
rect -15828 33948 -15812 34012
rect -15939 33932 -15812 33948
rect -15939 33868 -15892 33932
rect -15828 33868 -15812 33932
rect -15939 33852 -15812 33868
rect -15939 33788 -15892 33852
rect -15828 33788 -15812 33852
rect -15939 33772 -15812 33788
rect -15939 33708 -15892 33772
rect -15828 33708 -15812 33772
rect -15939 33692 -15812 33708
rect -15939 33628 -15892 33692
rect -15828 33628 -15812 33692
rect -15939 33612 -15812 33628
rect -15939 33548 -15892 33612
rect -15828 33548 -15812 33612
rect -15939 33532 -15812 33548
rect -15939 33468 -15892 33532
rect -15828 33468 -15812 33532
rect -15939 33452 -15812 33468
rect -15939 33388 -15892 33452
rect -15828 33388 -15812 33452
rect -15939 33372 -15812 33388
rect -15939 33308 -15892 33372
rect -15828 33308 -15812 33372
rect -15939 33292 -15812 33308
rect -15939 33228 -15892 33292
rect -15828 33228 -15812 33292
rect -15939 33212 -15812 33228
rect -15939 33148 -15892 33212
rect -15828 33148 -15812 33212
rect -15939 33132 -15812 33148
rect -15939 33068 -15892 33132
rect -15828 33068 -15812 33132
rect -15939 33052 -15812 33068
rect -15939 32988 -15892 33052
rect -15828 32988 -15812 33052
rect -15939 32972 -15812 32988
rect -15939 32908 -15892 32972
rect -15828 32908 -15812 32972
rect -15939 32892 -15812 32908
rect -15939 32828 -15892 32892
rect -15828 32828 -15812 32892
rect -15939 32812 -15812 32828
rect -15939 32748 -15892 32812
rect -15828 32748 -15812 32812
rect -15939 32732 -15812 32748
rect -15939 32668 -15892 32732
rect -15828 32668 -15812 32732
rect -15939 32652 -15812 32668
rect -15939 32588 -15892 32652
rect -15828 32588 -15812 32652
rect -15939 32572 -15812 32588
rect -15939 32508 -15892 32572
rect -15828 32508 -15812 32572
rect -15939 32492 -15812 32508
rect -15939 32428 -15892 32492
rect -15828 32428 -15812 32492
rect -15939 32412 -15812 32428
rect -15939 32348 -15892 32412
rect -15828 32348 -15812 32412
rect -15939 32332 -15812 32348
rect -15939 32268 -15892 32332
rect -15828 32268 -15812 32332
rect -15939 32252 -15812 32268
rect -15939 32188 -15892 32252
rect -15828 32188 -15812 32252
rect -15939 32172 -15812 32188
rect -15939 32108 -15892 32172
rect -15828 32108 -15812 32172
rect -15939 32092 -15812 32108
rect -15939 32028 -15892 32092
rect -15828 32028 -15812 32092
rect -15939 32012 -15812 32028
rect -15939 31948 -15892 32012
rect -15828 31948 -15812 32012
rect -15939 31932 -15812 31948
rect -15939 31868 -15892 31932
rect -15828 31868 -15812 31932
rect -15939 31852 -15812 31868
rect -15939 31788 -15892 31852
rect -15828 31788 -15812 31852
rect -15939 31772 -15812 31788
rect -15939 31708 -15892 31772
rect -15828 31708 -15812 31772
rect -15939 31692 -15812 31708
rect -15939 31628 -15892 31692
rect -15828 31628 -15812 31692
rect -15939 31612 -15812 31628
rect -15939 31548 -15892 31612
rect -15828 31548 -15812 31612
rect -15939 31532 -15812 31548
rect -15939 31468 -15892 31532
rect -15828 31468 -15812 31532
rect -15939 31452 -15812 31468
rect -15939 31388 -15892 31452
rect -15828 31388 -15812 31452
rect -15939 31372 -15812 31388
rect -15939 31308 -15892 31372
rect -15828 31308 -15812 31372
rect -15939 31292 -15812 31308
rect -15939 31228 -15892 31292
rect -15828 31228 -15812 31292
rect -15939 31212 -15812 31228
rect -15939 31148 -15892 31212
rect -15828 31148 -15812 31212
rect -15939 31132 -15812 31148
rect -15939 31068 -15892 31132
rect -15828 31068 -15812 31132
rect -15939 31052 -15812 31068
rect -15939 30988 -15892 31052
rect -15828 30988 -15812 31052
rect -15939 30972 -15812 30988
rect -15939 30908 -15892 30972
rect -15828 30908 -15812 30972
rect -15939 30892 -15812 30908
rect -15939 30828 -15892 30892
rect -15828 30828 -15812 30892
rect -15939 30812 -15812 30828
rect -15939 30748 -15892 30812
rect -15828 30748 -15812 30812
rect -15939 30732 -15812 30748
rect -15939 30668 -15892 30732
rect -15828 30668 -15812 30732
rect -15939 30652 -15812 30668
rect -15939 30588 -15892 30652
rect -15828 30588 -15812 30652
rect -15939 30572 -15812 30588
rect -15939 30508 -15892 30572
rect -15828 30508 -15812 30572
rect -15939 30492 -15812 30508
rect -15939 30428 -15892 30492
rect -15828 30428 -15812 30492
rect -15939 30412 -15812 30428
rect -15939 30348 -15892 30412
rect -15828 30348 -15812 30412
rect -15939 30332 -15812 30348
rect -15939 30268 -15892 30332
rect -15828 30268 -15812 30332
rect -15939 30252 -15812 30268
rect -15939 30188 -15892 30252
rect -15828 30188 -15812 30252
rect -15939 30172 -15812 30188
rect -15939 30108 -15892 30172
rect -15828 30108 -15812 30172
rect -15939 30092 -15812 30108
rect -15939 30028 -15892 30092
rect -15828 30028 -15812 30092
rect -15939 30012 -15812 30028
rect -15939 29948 -15892 30012
rect -15828 29948 -15812 30012
rect -15939 29932 -15812 29948
rect -15939 29868 -15892 29932
rect -15828 29868 -15812 29932
rect -15939 29852 -15812 29868
rect -15939 29788 -15892 29852
rect -15828 29788 -15812 29852
rect -15939 29772 -15812 29788
rect -15939 29708 -15892 29772
rect -15828 29708 -15812 29772
rect -15939 29692 -15812 29708
rect -15939 29628 -15892 29692
rect -15828 29628 -15812 29692
rect -15939 29612 -15812 29628
rect -15939 29548 -15892 29612
rect -15828 29548 -15812 29612
rect -15939 29532 -15812 29548
rect -15939 29468 -15892 29532
rect -15828 29468 -15812 29532
rect -15939 29452 -15812 29468
rect -15939 29388 -15892 29452
rect -15828 29388 -15812 29452
rect -15939 29372 -15812 29388
rect -15939 29308 -15892 29372
rect -15828 29308 -15812 29372
rect -15939 29292 -15812 29308
rect -15939 29228 -15892 29292
rect -15828 29228 -15812 29292
rect -15939 29212 -15812 29228
rect -15939 29148 -15892 29212
rect -15828 29148 -15812 29212
rect -15939 29132 -15812 29148
rect -15939 29068 -15892 29132
rect -15828 29068 -15812 29132
rect -15939 29052 -15812 29068
rect -15939 28988 -15892 29052
rect -15828 28988 -15812 29052
rect -15939 28972 -15812 28988
rect -15939 28908 -15892 28972
rect -15828 28908 -15812 28972
rect -15939 28892 -15812 28908
rect -15939 28828 -15892 28892
rect -15828 28828 -15812 28892
rect -15939 28812 -15812 28828
rect -15939 28748 -15892 28812
rect -15828 28748 -15812 28812
rect -15939 28732 -15812 28748
rect -15939 28668 -15892 28732
rect -15828 28668 -15812 28732
rect -15939 28652 -15812 28668
rect -15939 28588 -15892 28652
rect -15828 28588 -15812 28652
rect -15939 28572 -15812 28588
rect -22258 28492 -22131 28508
rect -22258 28428 -22211 28492
rect -22147 28428 -22131 28492
rect -22258 28412 -22131 28428
rect -22258 28288 -22154 28412
rect -22258 28272 -22131 28288
rect -22258 28208 -22211 28272
rect -22147 28208 -22131 28272
rect -22258 28192 -22131 28208
rect -28577 28112 -28450 28128
rect -28577 28048 -28530 28112
rect -28466 28048 -28450 28112
rect -28577 28032 -28450 28048
rect -28577 27968 -28530 28032
rect -28466 27968 -28450 28032
rect -28577 27952 -28450 27968
rect -28577 27888 -28530 27952
rect -28466 27888 -28450 27952
rect -28577 27872 -28450 27888
rect -28577 27808 -28530 27872
rect -28466 27808 -28450 27872
rect -28577 27792 -28450 27808
rect -28577 27728 -28530 27792
rect -28466 27728 -28450 27792
rect -28577 27712 -28450 27728
rect -28577 27648 -28530 27712
rect -28466 27648 -28450 27712
rect -28577 27632 -28450 27648
rect -28577 27568 -28530 27632
rect -28466 27568 -28450 27632
rect -28577 27552 -28450 27568
rect -28577 27488 -28530 27552
rect -28466 27488 -28450 27552
rect -28577 27472 -28450 27488
rect -28577 27408 -28530 27472
rect -28466 27408 -28450 27472
rect -28577 27392 -28450 27408
rect -28577 27328 -28530 27392
rect -28466 27328 -28450 27392
rect -28577 27312 -28450 27328
rect -28577 27248 -28530 27312
rect -28466 27248 -28450 27312
rect -28577 27232 -28450 27248
rect -28577 27168 -28530 27232
rect -28466 27168 -28450 27232
rect -28577 27152 -28450 27168
rect -28577 27088 -28530 27152
rect -28466 27088 -28450 27152
rect -28577 27072 -28450 27088
rect -28577 27008 -28530 27072
rect -28466 27008 -28450 27072
rect -28577 26992 -28450 27008
rect -28577 26928 -28530 26992
rect -28466 26928 -28450 26992
rect -28577 26912 -28450 26928
rect -28577 26848 -28530 26912
rect -28466 26848 -28450 26912
rect -28577 26832 -28450 26848
rect -28577 26768 -28530 26832
rect -28466 26768 -28450 26832
rect -28577 26752 -28450 26768
rect -28577 26688 -28530 26752
rect -28466 26688 -28450 26752
rect -28577 26672 -28450 26688
rect -28577 26608 -28530 26672
rect -28466 26608 -28450 26672
rect -28577 26592 -28450 26608
rect -28577 26528 -28530 26592
rect -28466 26528 -28450 26592
rect -28577 26512 -28450 26528
rect -28577 26448 -28530 26512
rect -28466 26448 -28450 26512
rect -28577 26432 -28450 26448
rect -28577 26368 -28530 26432
rect -28466 26368 -28450 26432
rect -28577 26352 -28450 26368
rect -28577 26288 -28530 26352
rect -28466 26288 -28450 26352
rect -28577 26272 -28450 26288
rect -28577 26208 -28530 26272
rect -28466 26208 -28450 26272
rect -28577 26192 -28450 26208
rect -28577 26128 -28530 26192
rect -28466 26128 -28450 26192
rect -28577 26112 -28450 26128
rect -28577 26048 -28530 26112
rect -28466 26048 -28450 26112
rect -28577 26032 -28450 26048
rect -28577 25968 -28530 26032
rect -28466 25968 -28450 26032
rect -28577 25952 -28450 25968
rect -28577 25888 -28530 25952
rect -28466 25888 -28450 25952
rect -28577 25872 -28450 25888
rect -28577 25808 -28530 25872
rect -28466 25808 -28450 25872
rect -28577 25792 -28450 25808
rect -28577 25728 -28530 25792
rect -28466 25728 -28450 25792
rect -28577 25712 -28450 25728
rect -28577 25648 -28530 25712
rect -28466 25648 -28450 25712
rect -28577 25632 -28450 25648
rect -28577 25568 -28530 25632
rect -28466 25568 -28450 25632
rect -28577 25552 -28450 25568
rect -28577 25488 -28530 25552
rect -28466 25488 -28450 25552
rect -28577 25472 -28450 25488
rect -28577 25408 -28530 25472
rect -28466 25408 -28450 25472
rect -28577 25392 -28450 25408
rect -28577 25328 -28530 25392
rect -28466 25328 -28450 25392
rect -28577 25312 -28450 25328
rect -28577 25248 -28530 25312
rect -28466 25248 -28450 25312
rect -28577 25232 -28450 25248
rect -28577 25168 -28530 25232
rect -28466 25168 -28450 25232
rect -28577 25152 -28450 25168
rect -28577 25088 -28530 25152
rect -28466 25088 -28450 25152
rect -28577 25072 -28450 25088
rect -28577 25008 -28530 25072
rect -28466 25008 -28450 25072
rect -28577 24992 -28450 25008
rect -28577 24928 -28530 24992
rect -28466 24928 -28450 24992
rect -28577 24912 -28450 24928
rect -28577 24848 -28530 24912
rect -28466 24848 -28450 24912
rect -28577 24832 -28450 24848
rect -28577 24768 -28530 24832
rect -28466 24768 -28450 24832
rect -28577 24752 -28450 24768
rect -28577 24688 -28530 24752
rect -28466 24688 -28450 24752
rect -28577 24672 -28450 24688
rect -28577 24608 -28530 24672
rect -28466 24608 -28450 24672
rect -28577 24592 -28450 24608
rect -28577 24528 -28530 24592
rect -28466 24528 -28450 24592
rect -28577 24512 -28450 24528
rect -28577 24448 -28530 24512
rect -28466 24448 -28450 24512
rect -28577 24432 -28450 24448
rect -28577 24368 -28530 24432
rect -28466 24368 -28450 24432
rect -28577 24352 -28450 24368
rect -28577 24288 -28530 24352
rect -28466 24288 -28450 24352
rect -28577 24272 -28450 24288
rect -28577 24208 -28530 24272
rect -28466 24208 -28450 24272
rect -28577 24192 -28450 24208
rect -28577 24128 -28530 24192
rect -28466 24128 -28450 24192
rect -28577 24112 -28450 24128
rect -28577 24048 -28530 24112
rect -28466 24048 -28450 24112
rect -28577 24032 -28450 24048
rect -28577 23968 -28530 24032
rect -28466 23968 -28450 24032
rect -28577 23952 -28450 23968
rect -28577 23888 -28530 23952
rect -28466 23888 -28450 23952
rect -28577 23872 -28450 23888
rect -28577 23808 -28530 23872
rect -28466 23808 -28450 23872
rect -28577 23792 -28450 23808
rect -28577 23728 -28530 23792
rect -28466 23728 -28450 23792
rect -28577 23712 -28450 23728
rect -28577 23648 -28530 23712
rect -28466 23648 -28450 23712
rect -28577 23632 -28450 23648
rect -28577 23568 -28530 23632
rect -28466 23568 -28450 23632
rect -28577 23552 -28450 23568
rect -28577 23488 -28530 23552
rect -28466 23488 -28450 23552
rect -28577 23472 -28450 23488
rect -28577 23408 -28530 23472
rect -28466 23408 -28450 23472
rect -28577 23392 -28450 23408
rect -28577 23328 -28530 23392
rect -28466 23328 -28450 23392
rect -28577 23312 -28450 23328
rect -28577 23248 -28530 23312
rect -28466 23248 -28450 23312
rect -28577 23232 -28450 23248
rect -28577 23168 -28530 23232
rect -28466 23168 -28450 23232
rect -28577 23152 -28450 23168
rect -28577 23088 -28530 23152
rect -28466 23088 -28450 23152
rect -28577 23072 -28450 23088
rect -28577 23008 -28530 23072
rect -28466 23008 -28450 23072
rect -28577 22992 -28450 23008
rect -28577 22928 -28530 22992
rect -28466 22928 -28450 22992
rect -28577 22912 -28450 22928
rect -28577 22848 -28530 22912
rect -28466 22848 -28450 22912
rect -28577 22832 -28450 22848
rect -28577 22768 -28530 22832
rect -28466 22768 -28450 22832
rect -28577 22752 -28450 22768
rect -28577 22688 -28530 22752
rect -28466 22688 -28450 22752
rect -28577 22672 -28450 22688
rect -28577 22608 -28530 22672
rect -28466 22608 -28450 22672
rect -28577 22592 -28450 22608
rect -28577 22528 -28530 22592
rect -28466 22528 -28450 22592
rect -28577 22512 -28450 22528
rect -28577 22448 -28530 22512
rect -28466 22448 -28450 22512
rect -28577 22432 -28450 22448
rect -28577 22368 -28530 22432
rect -28466 22368 -28450 22432
rect -28577 22352 -28450 22368
rect -28577 22288 -28530 22352
rect -28466 22288 -28450 22352
rect -28577 22272 -28450 22288
rect -34896 22192 -34769 22208
rect -34896 22128 -34849 22192
rect -34785 22128 -34769 22192
rect -34896 22112 -34769 22128
rect -34896 21988 -34792 22112
rect -34896 21972 -34769 21988
rect -34896 21908 -34849 21972
rect -34785 21908 -34769 21972
rect -34896 21892 -34769 21908
rect -41215 21812 -41088 21828
rect -41215 21748 -41168 21812
rect -41104 21748 -41088 21812
rect -41215 21732 -41088 21748
rect -41215 21668 -41168 21732
rect -41104 21668 -41088 21732
rect -41215 21652 -41088 21668
rect -41215 21588 -41168 21652
rect -41104 21588 -41088 21652
rect -41215 21572 -41088 21588
rect -41215 21508 -41168 21572
rect -41104 21508 -41088 21572
rect -41215 21492 -41088 21508
rect -41215 21428 -41168 21492
rect -41104 21428 -41088 21492
rect -41215 21412 -41088 21428
rect -41215 21348 -41168 21412
rect -41104 21348 -41088 21412
rect -41215 21332 -41088 21348
rect -41215 21268 -41168 21332
rect -41104 21268 -41088 21332
rect -41215 21252 -41088 21268
rect -41215 21188 -41168 21252
rect -41104 21188 -41088 21252
rect -41215 21172 -41088 21188
rect -41215 21108 -41168 21172
rect -41104 21108 -41088 21172
rect -41215 21092 -41088 21108
rect -41215 21028 -41168 21092
rect -41104 21028 -41088 21092
rect -41215 21012 -41088 21028
rect -41215 20948 -41168 21012
rect -41104 20948 -41088 21012
rect -41215 20932 -41088 20948
rect -41215 20868 -41168 20932
rect -41104 20868 -41088 20932
rect -41215 20852 -41088 20868
rect -41215 20788 -41168 20852
rect -41104 20788 -41088 20852
rect -41215 20772 -41088 20788
rect -41215 20708 -41168 20772
rect -41104 20708 -41088 20772
rect -41215 20692 -41088 20708
rect -41215 20628 -41168 20692
rect -41104 20628 -41088 20692
rect -41215 20612 -41088 20628
rect -41215 20548 -41168 20612
rect -41104 20548 -41088 20612
rect -41215 20532 -41088 20548
rect -41215 20468 -41168 20532
rect -41104 20468 -41088 20532
rect -41215 20452 -41088 20468
rect -41215 20388 -41168 20452
rect -41104 20388 -41088 20452
rect -41215 20372 -41088 20388
rect -41215 20308 -41168 20372
rect -41104 20308 -41088 20372
rect -41215 20292 -41088 20308
rect -41215 20228 -41168 20292
rect -41104 20228 -41088 20292
rect -41215 20212 -41088 20228
rect -41215 20148 -41168 20212
rect -41104 20148 -41088 20212
rect -41215 20132 -41088 20148
rect -41215 20068 -41168 20132
rect -41104 20068 -41088 20132
rect -41215 20052 -41088 20068
rect -41215 19988 -41168 20052
rect -41104 19988 -41088 20052
rect -41215 19972 -41088 19988
rect -41215 19908 -41168 19972
rect -41104 19908 -41088 19972
rect -41215 19892 -41088 19908
rect -41215 19828 -41168 19892
rect -41104 19828 -41088 19892
rect -41215 19812 -41088 19828
rect -41215 19748 -41168 19812
rect -41104 19748 -41088 19812
rect -41215 19732 -41088 19748
rect -41215 19668 -41168 19732
rect -41104 19668 -41088 19732
rect -41215 19652 -41088 19668
rect -41215 19588 -41168 19652
rect -41104 19588 -41088 19652
rect -41215 19572 -41088 19588
rect -41215 19508 -41168 19572
rect -41104 19508 -41088 19572
rect -41215 19492 -41088 19508
rect -41215 19428 -41168 19492
rect -41104 19428 -41088 19492
rect -41215 19412 -41088 19428
rect -41215 19348 -41168 19412
rect -41104 19348 -41088 19412
rect -41215 19332 -41088 19348
rect -41215 19268 -41168 19332
rect -41104 19268 -41088 19332
rect -41215 19252 -41088 19268
rect -41215 19188 -41168 19252
rect -41104 19188 -41088 19252
rect -41215 19172 -41088 19188
rect -41215 19108 -41168 19172
rect -41104 19108 -41088 19172
rect -41215 19092 -41088 19108
rect -41215 19028 -41168 19092
rect -41104 19028 -41088 19092
rect -41215 19012 -41088 19028
rect -41215 18948 -41168 19012
rect -41104 18948 -41088 19012
rect -41215 18932 -41088 18948
rect -41215 18868 -41168 18932
rect -41104 18868 -41088 18932
rect -41215 18852 -41088 18868
rect -41215 18788 -41168 18852
rect -41104 18788 -41088 18852
rect -41215 18772 -41088 18788
rect -41215 18708 -41168 18772
rect -41104 18708 -41088 18772
rect -41215 18692 -41088 18708
rect -41215 18628 -41168 18692
rect -41104 18628 -41088 18692
rect -41215 18612 -41088 18628
rect -41215 18548 -41168 18612
rect -41104 18548 -41088 18612
rect -41215 18532 -41088 18548
rect -41215 18468 -41168 18532
rect -41104 18468 -41088 18532
rect -41215 18452 -41088 18468
rect -41215 18388 -41168 18452
rect -41104 18388 -41088 18452
rect -41215 18372 -41088 18388
rect -41215 18308 -41168 18372
rect -41104 18308 -41088 18372
rect -41215 18292 -41088 18308
rect -41215 18228 -41168 18292
rect -41104 18228 -41088 18292
rect -41215 18212 -41088 18228
rect -41215 18148 -41168 18212
rect -41104 18148 -41088 18212
rect -41215 18132 -41088 18148
rect -41215 18068 -41168 18132
rect -41104 18068 -41088 18132
rect -41215 18052 -41088 18068
rect -41215 17988 -41168 18052
rect -41104 17988 -41088 18052
rect -41215 17972 -41088 17988
rect -41215 17908 -41168 17972
rect -41104 17908 -41088 17972
rect -41215 17892 -41088 17908
rect -41215 17828 -41168 17892
rect -41104 17828 -41088 17892
rect -41215 17812 -41088 17828
rect -41215 17748 -41168 17812
rect -41104 17748 -41088 17812
rect -41215 17732 -41088 17748
rect -41215 17668 -41168 17732
rect -41104 17668 -41088 17732
rect -41215 17652 -41088 17668
rect -41215 17588 -41168 17652
rect -41104 17588 -41088 17652
rect -41215 17572 -41088 17588
rect -41215 17508 -41168 17572
rect -41104 17508 -41088 17572
rect -41215 17492 -41088 17508
rect -41215 17428 -41168 17492
rect -41104 17428 -41088 17492
rect -41215 17412 -41088 17428
rect -41215 17348 -41168 17412
rect -41104 17348 -41088 17412
rect -41215 17332 -41088 17348
rect -41215 17268 -41168 17332
rect -41104 17268 -41088 17332
rect -41215 17252 -41088 17268
rect -41215 17188 -41168 17252
rect -41104 17188 -41088 17252
rect -41215 17172 -41088 17188
rect -41215 17108 -41168 17172
rect -41104 17108 -41088 17172
rect -41215 17092 -41088 17108
rect -41215 17028 -41168 17092
rect -41104 17028 -41088 17092
rect -41215 17012 -41088 17028
rect -41215 16948 -41168 17012
rect -41104 16948 -41088 17012
rect -41215 16932 -41088 16948
rect -41215 16868 -41168 16932
rect -41104 16868 -41088 16932
rect -41215 16852 -41088 16868
rect -41215 16788 -41168 16852
rect -41104 16788 -41088 16852
rect -41215 16772 -41088 16788
rect -41215 16708 -41168 16772
rect -41104 16708 -41088 16772
rect -41215 16692 -41088 16708
rect -41215 16628 -41168 16692
rect -41104 16628 -41088 16692
rect -41215 16612 -41088 16628
rect -41215 16548 -41168 16612
rect -41104 16548 -41088 16612
rect -41215 16532 -41088 16548
rect -41215 16468 -41168 16532
rect -41104 16468 -41088 16532
rect -41215 16452 -41088 16468
rect -41215 16388 -41168 16452
rect -41104 16388 -41088 16452
rect -41215 16372 -41088 16388
rect -41215 16308 -41168 16372
rect -41104 16308 -41088 16372
rect -41215 16292 -41088 16308
rect -41215 16228 -41168 16292
rect -41104 16228 -41088 16292
rect -41215 16212 -41088 16228
rect -41215 16148 -41168 16212
rect -41104 16148 -41088 16212
rect -41215 16132 -41088 16148
rect -41215 16068 -41168 16132
rect -41104 16068 -41088 16132
rect -41215 16052 -41088 16068
rect -41215 15988 -41168 16052
rect -41104 15988 -41088 16052
rect -41215 15972 -41088 15988
rect -44335 15561 -44231 15939
rect -41215 15908 -41168 15972
rect -41104 15908 -41088 15972
rect -40925 21852 -35003 21861
rect -40925 15948 -40916 21852
rect -35012 15948 -35003 21852
rect -40925 15939 -35003 15948
rect -34896 21828 -34849 21892
rect -34785 21828 -34769 21892
rect -31697 21861 -31593 22239
rect -28577 22208 -28530 22272
rect -28466 22208 -28450 22272
rect -28287 28152 -22365 28161
rect -28287 22248 -28278 28152
rect -22374 22248 -22365 28152
rect -28287 22239 -22365 22248
rect -22258 28128 -22211 28192
rect -22147 28128 -22131 28192
rect -19059 28161 -18955 28539
rect -15939 28508 -15892 28572
rect -15828 28508 -15812 28572
rect -15649 34452 -9727 34461
rect -15649 28548 -15640 34452
rect -9736 28548 -9727 34452
rect -15649 28539 -9727 28548
rect -9620 34428 -9573 34492
rect -9509 34428 -9493 34492
rect -6421 34461 -6317 34839
rect -3301 34808 -3254 34872
rect -3190 34808 -3174 34872
rect -3011 40752 2911 40761
rect -3011 34848 -3002 40752
rect 2902 34848 2911 40752
rect -3011 34839 2911 34848
rect 3018 40728 3065 40792
rect 3129 40728 3145 40792
rect 6217 40761 6321 41139
rect 9337 41108 9384 41172
rect 9448 41108 9464 41172
rect 9627 47052 15549 47061
rect 9627 41148 9636 47052
rect 15540 41148 15549 47052
rect 9627 41139 15549 41148
rect 15656 47028 15703 47092
rect 15767 47028 15783 47092
rect 18855 47061 18959 47250
rect 21975 47188 22079 47250
rect 21975 47172 22102 47188
rect 21975 47108 22022 47172
rect 22086 47108 22102 47172
rect 21975 47092 22102 47108
rect 15656 47012 15783 47028
rect 15656 46948 15703 47012
rect 15767 46948 15783 47012
rect 15656 46932 15783 46948
rect 15656 46868 15703 46932
rect 15767 46868 15783 46932
rect 15656 46852 15783 46868
rect 15656 46788 15703 46852
rect 15767 46788 15783 46852
rect 15656 46772 15783 46788
rect 15656 46708 15703 46772
rect 15767 46708 15783 46772
rect 15656 46692 15783 46708
rect 15656 46628 15703 46692
rect 15767 46628 15783 46692
rect 15656 46612 15783 46628
rect 15656 46548 15703 46612
rect 15767 46548 15783 46612
rect 15656 46532 15783 46548
rect 15656 46468 15703 46532
rect 15767 46468 15783 46532
rect 15656 46452 15783 46468
rect 15656 46388 15703 46452
rect 15767 46388 15783 46452
rect 15656 46372 15783 46388
rect 15656 46308 15703 46372
rect 15767 46308 15783 46372
rect 15656 46292 15783 46308
rect 15656 46228 15703 46292
rect 15767 46228 15783 46292
rect 15656 46212 15783 46228
rect 15656 46148 15703 46212
rect 15767 46148 15783 46212
rect 15656 46132 15783 46148
rect 15656 46068 15703 46132
rect 15767 46068 15783 46132
rect 15656 46052 15783 46068
rect 15656 45988 15703 46052
rect 15767 45988 15783 46052
rect 15656 45972 15783 45988
rect 15656 45908 15703 45972
rect 15767 45908 15783 45972
rect 15656 45892 15783 45908
rect 15656 45828 15703 45892
rect 15767 45828 15783 45892
rect 15656 45812 15783 45828
rect 15656 45748 15703 45812
rect 15767 45748 15783 45812
rect 15656 45732 15783 45748
rect 15656 45668 15703 45732
rect 15767 45668 15783 45732
rect 15656 45652 15783 45668
rect 15656 45588 15703 45652
rect 15767 45588 15783 45652
rect 15656 45572 15783 45588
rect 15656 45508 15703 45572
rect 15767 45508 15783 45572
rect 15656 45492 15783 45508
rect 15656 45428 15703 45492
rect 15767 45428 15783 45492
rect 15656 45412 15783 45428
rect 15656 45348 15703 45412
rect 15767 45348 15783 45412
rect 15656 45332 15783 45348
rect 15656 45268 15703 45332
rect 15767 45268 15783 45332
rect 15656 45252 15783 45268
rect 15656 45188 15703 45252
rect 15767 45188 15783 45252
rect 15656 45172 15783 45188
rect 15656 45108 15703 45172
rect 15767 45108 15783 45172
rect 15656 45092 15783 45108
rect 15656 45028 15703 45092
rect 15767 45028 15783 45092
rect 15656 45012 15783 45028
rect 15656 44948 15703 45012
rect 15767 44948 15783 45012
rect 15656 44932 15783 44948
rect 15656 44868 15703 44932
rect 15767 44868 15783 44932
rect 15656 44852 15783 44868
rect 15656 44788 15703 44852
rect 15767 44788 15783 44852
rect 15656 44772 15783 44788
rect 15656 44708 15703 44772
rect 15767 44708 15783 44772
rect 15656 44692 15783 44708
rect 15656 44628 15703 44692
rect 15767 44628 15783 44692
rect 15656 44612 15783 44628
rect 15656 44548 15703 44612
rect 15767 44548 15783 44612
rect 15656 44532 15783 44548
rect 15656 44468 15703 44532
rect 15767 44468 15783 44532
rect 15656 44452 15783 44468
rect 15656 44388 15703 44452
rect 15767 44388 15783 44452
rect 15656 44372 15783 44388
rect 15656 44308 15703 44372
rect 15767 44308 15783 44372
rect 15656 44292 15783 44308
rect 15656 44228 15703 44292
rect 15767 44228 15783 44292
rect 15656 44212 15783 44228
rect 15656 44148 15703 44212
rect 15767 44148 15783 44212
rect 15656 44132 15783 44148
rect 15656 44068 15703 44132
rect 15767 44068 15783 44132
rect 15656 44052 15783 44068
rect 15656 43988 15703 44052
rect 15767 43988 15783 44052
rect 15656 43972 15783 43988
rect 15656 43908 15703 43972
rect 15767 43908 15783 43972
rect 15656 43892 15783 43908
rect 15656 43828 15703 43892
rect 15767 43828 15783 43892
rect 15656 43812 15783 43828
rect 15656 43748 15703 43812
rect 15767 43748 15783 43812
rect 15656 43732 15783 43748
rect 15656 43668 15703 43732
rect 15767 43668 15783 43732
rect 15656 43652 15783 43668
rect 15656 43588 15703 43652
rect 15767 43588 15783 43652
rect 15656 43572 15783 43588
rect 15656 43508 15703 43572
rect 15767 43508 15783 43572
rect 15656 43492 15783 43508
rect 15656 43428 15703 43492
rect 15767 43428 15783 43492
rect 15656 43412 15783 43428
rect 15656 43348 15703 43412
rect 15767 43348 15783 43412
rect 15656 43332 15783 43348
rect 15656 43268 15703 43332
rect 15767 43268 15783 43332
rect 15656 43252 15783 43268
rect 15656 43188 15703 43252
rect 15767 43188 15783 43252
rect 15656 43172 15783 43188
rect 15656 43108 15703 43172
rect 15767 43108 15783 43172
rect 15656 43092 15783 43108
rect 15656 43028 15703 43092
rect 15767 43028 15783 43092
rect 15656 43012 15783 43028
rect 15656 42948 15703 43012
rect 15767 42948 15783 43012
rect 15656 42932 15783 42948
rect 15656 42868 15703 42932
rect 15767 42868 15783 42932
rect 15656 42852 15783 42868
rect 15656 42788 15703 42852
rect 15767 42788 15783 42852
rect 15656 42772 15783 42788
rect 15656 42708 15703 42772
rect 15767 42708 15783 42772
rect 15656 42692 15783 42708
rect 15656 42628 15703 42692
rect 15767 42628 15783 42692
rect 15656 42612 15783 42628
rect 15656 42548 15703 42612
rect 15767 42548 15783 42612
rect 15656 42532 15783 42548
rect 15656 42468 15703 42532
rect 15767 42468 15783 42532
rect 15656 42452 15783 42468
rect 15656 42388 15703 42452
rect 15767 42388 15783 42452
rect 15656 42372 15783 42388
rect 15656 42308 15703 42372
rect 15767 42308 15783 42372
rect 15656 42292 15783 42308
rect 15656 42228 15703 42292
rect 15767 42228 15783 42292
rect 15656 42212 15783 42228
rect 15656 42148 15703 42212
rect 15767 42148 15783 42212
rect 15656 42132 15783 42148
rect 15656 42068 15703 42132
rect 15767 42068 15783 42132
rect 15656 42052 15783 42068
rect 15656 41988 15703 42052
rect 15767 41988 15783 42052
rect 15656 41972 15783 41988
rect 15656 41908 15703 41972
rect 15767 41908 15783 41972
rect 15656 41892 15783 41908
rect 15656 41828 15703 41892
rect 15767 41828 15783 41892
rect 15656 41812 15783 41828
rect 15656 41748 15703 41812
rect 15767 41748 15783 41812
rect 15656 41732 15783 41748
rect 15656 41668 15703 41732
rect 15767 41668 15783 41732
rect 15656 41652 15783 41668
rect 15656 41588 15703 41652
rect 15767 41588 15783 41652
rect 15656 41572 15783 41588
rect 15656 41508 15703 41572
rect 15767 41508 15783 41572
rect 15656 41492 15783 41508
rect 15656 41428 15703 41492
rect 15767 41428 15783 41492
rect 15656 41412 15783 41428
rect 15656 41348 15703 41412
rect 15767 41348 15783 41412
rect 15656 41332 15783 41348
rect 15656 41268 15703 41332
rect 15767 41268 15783 41332
rect 15656 41252 15783 41268
rect 15656 41188 15703 41252
rect 15767 41188 15783 41252
rect 15656 41172 15783 41188
rect 9337 41092 9464 41108
rect 9337 41028 9384 41092
rect 9448 41028 9464 41092
rect 9337 41012 9464 41028
rect 9337 40888 9441 41012
rect 9337 40872 9464 40888
rect 9337 40808 9384 40872
rect 9448 40808 9464 40872
rect 9337 40792 9464 40808
rect 3018 40712 3145 40728
rect 3018 40648 3065 40712
rect 3129 40648 3145 40712
rect 3018 40632 3145 40648
rect 3018 40568 3065 40632
rect 3129 40568 3145 40632
rect 3018 40552 3145 40568
rect 3018 40488 3065 40552
rect 3129 40488 3145 40552
rect 3018 40472 3145 40488
rect 3018 40408 3065 40472
rect 3129 40408 3145 40472
rect 3018 40392 3145 40408
rect 3018 40328 3065 40392
rect 3129 40328 3145 40392
rect 3018 40312 3145 40328
rect 3018 40248 3065 40312
rect 3129 40248 3145 40312
rect 3018 40232 3145 40248
rect 3018 40168 3065 40232
rect 3129 40168 3145 40232
rect 3018 40152 3145 40168
rect 3018 40088 3065 40152
rect 3129 40088 3145 40152
rect 3018 40072 3145 40088
rect 3018 40008 3065 40072
rect 3129 40008 3145 40072
rect 3018 39992 3145 40008
rect 3018 39928 3065 39992
rect 3129 39928 3145 39992
rect 3018 39912 3145 39928
rect 3018 39848 3065 39912
rect 3129 39848 3145 39912
rect 3018 39832 3145 39848
rect 3018 39768 3065 39832
rect 3129 39768 3145 39832
rect 3018 39752 3145 39768
rect 3018 39688 3065 39752
rect 3129 39688 3145 39752
rect 3018 39672 3145 39688
rect 3018 39608 3065 39672
rect 3129 39608 3145 39672
rect 3018 39592 3145 39608
rect 3018 39528 3065 39592
rect 3129 39528 3145 39592
rect 3018 39512 3145 39528
rect 3018 39448 3065 39512
rect 3129 39448 3145 39512
rect 3018 39432 3145 39448
rect 3018 39368 3065 39432
rect 3129 39368 3145 39432
rect 3018 39352 3145 39368
rect 3018 39288 3065 39352
rect 3129 39288 3145 39352
rect 3018 39272 3145 39288
rect 3018 39208 3065 39272
rect 3129 39208 3145 39272
rect 3018 39192 3145 39208
rect 3018 39128 3065 39192
rect 3129 39128 3145 39192
rect 3018 39112 3145 39128
rect 3018 39048 3065 39112
rect 3129 39048 3145 39112
rect 3018 39032 3145 39048
rect 3018 38968 3065 39032
rect 3129 38968 3145 39032
rect 3018 38952 3145 38968
rect 3018 38888 3065 38952
rect 3129 38888 3145 38952
rect 3018 38872 3145 38888
rect 3018 38808 3065 38872
rect 3129 38808 3145 38872
rect 3018 38792 3145 38808
rect 3018 38728 3065 38792
rect 3129 38728 3145 38792
rect 3018 38712 3145 38728
rect 3018 38648 3065 38712
rect 3129 38648 3145 38712
rect 3018 38632 3145 38648
rect 3018 38568 3065 38632
rect 3129 38568 3145 38632
rect 3018 38552 3145 38568
rect 3018 38488 3065 38552
rect 3129 38488 3145 38552
rect 3018 38472 3145 38488
rect 3018 38408 3065 38472
rect 3129 38408 3145 38472
rect 3018 38392 3145 38408
rect 3018 38328 3065 38392
rect 3129 38328 3145 38392
rect 3018 38312 3145 38328
rect 3018 38248 3065 38312
rect 3129 38248 3145 38312
rect 3018 38232 3145 38248
rect 3018 38168 3065 38232
rect 3129 38168 3145 38232
rect 3018 38152 3145 38168
rect 3018 38088 3065 38152
rect 3129 38088 3145 38152
rect 3018 38072 3145 38088
rect 3018 38008 3065 38072
rect 3129 38008 3145 38072
rect 3018 37992 3145 38008
rect 3018 37928 3065 37992
rect 3129 37928 3145 37992
rect 3018 37912 3145 37928
rect 3018 37848 3065 37912
rect 3129 37848 3145 37912
rect 3018 37832 3145 37848
rect 3018 37768 3065 37832
rect 3129 37768 3145 37832
rect 3018 37752 3145 37768
rect 3018 37688 3065 37752
rect 3129 37688 3145 37752
rect 3018 37672 3145 37688
rect 3018 37608 3065 37672
rect 3129 37608 3145 37672
rect 3018 37592 3145 37608
rect 3018 37528 3065 37592
rect 3129 37528 3145 37592
rect 3018 37512 3145 37528
rect 3018 37448 3065 37512
rect 3129 37448 3145 37512
rect 3018 37432 3145 37448
rect 3018 37368 3065 37432
rect 3129 37368 3145 37432
rect 3018 37352 3145 37368
rect 3018 37288 3065 37352
rect 3129 37288 3145 37352
rect 3018 37272 3145 37288
rect 3018 37208 3065 37272
rect 3129 37208 3145 37272
rect 3018 37192 3145 37208
rect 3018 37128 3065 37192
rect 3129 37128 3145 37192
rect 3018 37112 3145 37128
rect 3018 37048 3065 37112
rect 3129 37048 3145 37112
rect 3018 37032 3145 37048
rect 3018 36968 3065 37032
rect 3129 36968 3145 37032
rect 3018 36952 3145 36968
rect 3018 36888 3065 36952
rect 3129 36888 3145 36952
rect 3018 36872 3145 36888
rect 3018 36808 3065 36872
rect 3129 36808 3145 36872
rect 3018 36792 3145 36808
rect 3018 36728 3065 36792
rect 3129 36728 3145 36792
rect 3018 36712 3145 36728
rect 3018 36648 3065 36712
rect 3129 36648 3145 36712
rect 3018 36632 3145 36648
rect 3018 36568 3065 36632
rect 3129 36568 3145 36632
rect 3018 36552 3145 36568
rect 3018 36488 3065 36552
rect 3129 36488 3145 36552
rect 3018 36472 3145 36488
rect 3018 36408 3065 36472
rect 3129 36408 3145 36472
rect 3018 36392 3145 36408
rect 3018 36328 3065 36392
rect 3129 36328 3145 36392
rect 3018 36312 3145 36328
rect 3018 36248 3065 36312
rect 3129 36248 3145 36312
rect 3018 36232 3145 36248
rect 3018 36168 3065 36232
rect 3129 36168 3145 36232
rect 3018 36152 3145 36168
rect 3018 36088 3065 36152
rect 3129 36088 3145 36152
rect 3018 36072 3145 36088
rect 3018 36008 3065 36072
rect 3129 36008 3145 36072
rect 3018 35992 3145 36008
rect 3018 35928 3065 35992
rect 3129 35928 3145 35992
rect 3018 35912 3145 35928
rect 3018 35848 3065 35912
rect 3129 35848 3145 35912
rect 3018 35832 3145 35848
rect 3018 35768 3065 35832
rect 3129 35768 3145 35832
rect 3018 35752 3145 35768
rect 3018 35688 3065 35752
rect 3129 35688 3145 35752
rect 3018 35672 3145 35688
rect 3018 35608 3065 35672
rect 3129 35608 3145 35672
rect 3018 35592 3145 35608
rect 3018 35528 3065 35592
rect 3129 35528 3145 35592
rect 3018 35512 3145 35528
rect 3018 35448 3065 35512
rect 3129 35448 3145 35512
rect 3018 35432 3145 35448
rect 3018 35368 3065 35432
rect 3129 35368 3145 35432
rect 3018 35352 3145 35368
rect 3018 35288 3065 35352
rect 3129 35288 3145 35352
rect 3018 35272 3145 35288
rect 3018 35208 3065 35272
rect 3129 35208 3145 35272
rect 3018 35192 3145 35208
rect 3018 35128 3065 35192
rect 3129 35128 3145 35192
rect 3018 35112 3145 35128
rect 3018 35048 3065 35112
rect 3129 35048 3145 35112
rect 3018 35032 3145 35048
rect 3018 34968 3065 35032
rect 3129 34968 3145 35032
rect 3018 34952 3145 34968
rect 3018 34888 3065 34952
rect 3129 34888 3145 34952
rect 3018 34872 3145 34888
rect -3301 34792 -3174 34808
rect -3301 34728 -3254 34792
rect -3190 34728 -3174 34792
rect -3301 34712 -3174 34728
rect -3301 34588 -3197 34712
rect -3301 34572 -3174 34588
rect -3301 34508 -3254 34572
rect -3190 34508 -3174 34572
rect -3301 34492 -3174 34508
rect -9620 34412 -9493 34428
rect -9620 34348 -9573 34412
rect -9509 34348 -9493 34412
rect -9620 34332 -9493 34348
rect -9620 34268 -9573 34332
rect -9509 34268 -9493 34332
rect -9620 34252 -9493 34268
rect -9620 34188 -9573 34252
rect -9509 34188 -9493 34252
rect -9620 34172 -9493 34188
rect -9620 34108 -9573 34172
rect -9509 34108 -9493 34172
rect -9620 34092 -9493 34108
rect -9620 34028 -9573 34092
rect -9509 34028 -9493 34092
rect -9620 34012 -9493 34028
rect -9620 33948 -9573 34012
rect -9509 33948 -9493 34012
rect -9620 33932 -9493 33948
rect -9620 33868 -9573 33932
rect -9509 33868 -9493 33932
rect -9620 33852 -9493 33868
rect -9620 33788 -9573 33852
rect -9509 33788 -9493 33852
rect -9620 33772 -9493 33788
rect -9620 33708 -9573 33772
rect -9509 33708 -9493 33772
rect -9620 33692 -9493 33708
rect -9620 33628 -9573 33692
rect -9509 33628 -9493 33692
rect -9620 33612 -9493 33628
rect -9620 33548 -9573 33612
rect -9509 33548 -9493 33612
rect -9620 33532 -9493 33548
rect -9620 33468 -9573 33532
rect -9509 33468 -9493 33532
rect -9620 33452 -9493 33468
rect -9620 33388 -9573 33452
rect -9509 33388 -9493 33452
rect -9620 33372 -9493 33388
rect -9620 33308 -9573 33372
rect -9509 33308 -9493 33372
rect -9620 33292 -9493 33308
rect -9620 33228 -9573 33292
rect -9509 33228 -9493 33292
rect -9620 33212 -9493 33228
rect -9620 33148 -9573 33212
rect -9509 33148 -9493 33212
rect -9620 33132 -9493 33148
rect -9620 33068 -9573 33132
rect -9509 33068 -9493 33132
rect -9620 33052 -9493 33068
rect -9620 32988 -9573 33052
rect -9509 32988 -9493 33052
rect -9620 32972 -9493 32988
rect -9620 32908 -9573 32972
rect -9509 32908 -9493 32972
rect -9620 32892 -9493 32908
rect -9620 32828 -9573 32892
rect -9509 32828 -9493 32892
rect -9620 32812 -9493 32828
rect -9620 32748 -9573 32812
rect -9509 32748 -9493 32812
rect -9620 32732 -9493 32748
rect -9620 32668 -9573 32732
rect -9509 32668 -9493 32732
rect -9620 32652 -9493 32668
rect -9620 32588 -9573 32652
rect -9509 32588 -9493 32652
rect -9620 32572 -9493 32588
rect -9620 32508 -9573 32572
rect -9509 32508 -9493 32572
rect -9620 32492 -9493 32508
rect -9620 32428 -9573 32492
rect -9509 32428 -9493 32492
rect -9620 32412 -9493 32428
rect -9620 32348 -9573 32412
rect -9509 32348 -9493 32412
rect -9620 32332 -9493 32348
rect -9620 32268 -9573 32332
rect -9509 32268 -9493 32332
rect -9620 32252 -9493 32268
rect -9620 32188 -9573 32252
rect -9509 32188 -9493 32252
rect -9620 32172 -9493 32188
rect -9620 32108 -9573 32172
rect -9509 32108 -9493 32172
rect -9620 32092 -9493 32108
rect -9620 32028 -9573 32092
rect -9509 32028 -9493 32092
rect -9620 32012 -9493 32028
rect -9620 31948 -9573 32012
rect -9509 31948 -9493 32012
rect -9620 31932 -9493 31948
rect -9620 31868 -9573 31932
rect -9509 31868 -9493 31932
rect -9620 31852 -9493 31868
rect -9620 31788 -9573 31852
rect -9509 31788 -9493 31852
rect -9620 31772 -9493 31788
rect -9620 31708 -9573 31772
rect -9509 31708 -9493 31772
rect -9620 31692 -9493 31708
rect -9620 31628 -9573 31692
rect -9509 31628 -9493 31692
rect -9620 31612 -9493 31628
rect -9620 31548 -9573 31612
rect -9509 31548 -9493 31612
rect -9620 31532 -9493 31548
rect -9620 31468 -9573 31532
rect -9509 31468 -9493 31532
rect -9620 31452 -9493 31468
rect -9620 31388 -9573 31452
rect -9509 31388 -9493 31452
rect -9620 31372 -9493 31388
rect -9620 31308 -9573 31372
rect -9509 31308 -9493 31372
rect -9620 31292 -9493 31308
rect -9620 31228 -9573 31292
rect -9509 31228 -9493 31292
rect -9620 31212 -9493 31228
rect -9620 31148 -9573 31212
rect -9509 31148 -9493 31212
rect -9620 31132 -9493 31148
rect -9620 31068 -9573 31132
rect -9509 31068 -9493 31132
rect -9620 31052 -9493 31068
rect -9620 30988 -9573 31052
rect -9509 30988 -9493 31052
rect -9620 30972 -9493 30988
rect -9620 30908 -9573 30972
rect -9509 30908 -9493 30972
rect -9620 30892 -9493 30908
rect -9620 30828 -9573 30892
rect -9509 30828 -9493 30892
rect -9620 30812 -9493 30828
rect -9620 30748 -9573 30812
rect -9509 30748 -9493 30812
rect -9620 30732 -9493 30748
rect -9620 30668 -9573 30732
rect -9509 30668 -9493 30732
rect -9620 30652 -9493 30668
rect -9620 30588 -9573 30652
rect -9509 30588 -9493 30652
rect -9620 30572 -9493 30588
rect -9620 30508 -9573 30572
rect -9509 30508 -9493 30572
rect -9620 30492 -9493 30508
rect -9620 30428 -9573 30492
rect -9509 30428 -9493 30492
rect -9620 30412 -9493 30428
rect -9620 30348 -9573 30412
rect -9509 30348 -9493 30412
rect -9620 30332 -9493 30348
rect -9620 30268 -9573 30332
rect -9509 30268 -9493 30332
rect -9620 30252 -9493 30268
rect -9620 30188 -9573 30252
rect -9509 30188 -9493 30252
rect -9620 30172 -9493 30188
rect -9620 30108 -9573 30172
rect -9509 30108 -9493 30172
rect -9620 30092 -9493 30108
rect -9620 30028 -9573 30092
rect -9509 30028 -9493 30092
rect -9620 30012 -9493 30028
rect -9620 29948 -9573 30012
rect -9509 29948 -9493 30012
rect -9620 29932 -9493 29948
rect -9620 29868 -9573 29932
rect -9509 29868 -9493 29932
rect -9620 29852 -9493 29868
rect -9620 29788 -9573 29852
rect -9509 29788 -9493 29852
rect -9620 29772 -9493 29788
rect -9620 29708 -9573 29772
rect -9509 29708 -9493 29772
rect -9620 29692 -9493 29708
rect -9620 29628 -9573 29692
rect -9509 29628 -9493 29692
rect -9620 29612 -9493 29628
rect -9620 29548 -9573 29612
rect -9509 29548 -9493 29612
rect -9620 29532 -9493 29548
rect -9620 29468 -9573 29532
rect -9509 29468 -9493 29532
rect -9620 29452 -9493 29468
rect -9620 29388 -9573 29452
rect -9509 29388 -9493 29452
rect -9620 29372 -9493 29388
rect -9620 29308 -9573 29372
rect -9509 29308 -9493 29372
rect -9620 29292 -9493 29308
rect -9620 29228 -9573 29292
rect -9509 29228 -9493 29292
rect -9620 29212 -9493 29228
rect -9620 29148 -9573 29212
rect -9509 29148 -9493 29212
rect -9620 29132 -9493 29148
rect -9620 29068 -9573 29132
rect -9509 29068 -9493 29132
rect -9620 29052 -9493 29068
rect -9620 28988 -9573 29052
rect -9509 28988 -9493 29052
rect -9620 28972 -9493 28988
rect -9620 28908 -9573 28972
rect -9509 28908 -9493 28972
rect -9620 28892 -9493 28908
rect -9620 28828 -9573 28892
rect -9509 28828 -9493 28892
rect -9620 28812 -9493 28828
rect -9620 28748 -9573 28812
rect -9509 28748 -9493 28812
rect -9620 28732 -9493 28748
rect -9620 28668 -9573 28732
rect -9509 28668 -9493 28732
rect -9620 28652 -9493 28668
rect -9620 28588 -9573 28652
rect -9509 28588 -9493 28652
rect -9620 28572 -9493 28588
rect -15939 28492 -15812 28508
rect -15939 28428 -15892 28492
rect -15828 28428 -15812 28492
rect -15939 28412 -15812 28428
rect -15939 28288 -15835 28412
rect -15939 28272 -15812 28288
rect -15939 28208 -15892 28272
rect -15828 28208 -15812 28272
rect -15939 28192 -15812 28208
rect -22258 28112 -22131 28128
rect -22258 28048 -22211 28112
rect -22147 28048 -22131 28112
rect -22258 28032 -22131 28048
rect -22258 27968 -22211 28032
rect -22147 27968 -22131 28032
rect -22258 27952 -22131 27968
rect -22258 27888 -22211 27952
rect -22147 27888 -22131 27952
rect -22258 27872 -22131 27888
rect -22258 27808 -22211 27872
rect -22147 27808 -22131 27872
rect -22258 27792 -22131 27808
rect -22258 27728 -22211 27792
rect -22147 27728 -22131 27792
rect -22258 27712 -22131 27728
rect -22258 27648 -22211 27712
rect -22147 27648 -22131 27712
rect -22258 27632 -22131 27648
rect -22258 27568 -22211 27632
rect -22147 27568 -22131 27632
rect -22258 27552 -22131 27568
rect -22258 27488 -22211 27552
rect -22147 27488 -22131 27552
rect -22258 27472 -22131 27488
rect -22258 27408 -22211 27472
rect -22147 27408 -22131 27472
rect -22258 27392 -22131 27408
rect -22258 27328 -22211 27392
rect -22147 27328 -22131 27392
rect -22258 27312 -22131 27328
rect -22258 27248 -22211 27312
rect -22147 27248 -22131 27312
rect -22258 27232 -22131 27248
rect -22258 27168 -22211 27232
rect -22147 27168 -22131 27232
rect -22258 27152 -22131 27168
rect -22258 27088 -22211 27152
rect -22147 27088 -22131 27152
rect -22258 27072 -22131 27088
rect -22258 27008 -22211 27072
rect -22147 27008 -22131 27072
rect -22258 26992 -22131 27008
rect -22258 26928 -22211 26992
rect -22147 26928 -22131 26992
rect -22258 26912 -22131 26928
rect -22258 26848 -22211 26912
rect -22147 26848 -22131 26912
rect -22258 26832 -22131 26848
rect -22258 26768 -22211 26832
rect -22147 26768 -22131 26832
rect -22258 26752 -22131 26768
rect -22258 26688 -22211 26752
rect -22147 26688 -22131 26752
rect -22258 26672 -22131 26688
rect -22258 26608 -22211 26672
rect -22147 26608 -22131 26672
rect -22258 26592 -22131 26608
rect -22258 26528 -22211 26592
rect -22147 26528 -22131 26592
rect -22258 26512 -22131 26528
rect -22258 26448 -22211 26512
rect -22147 26448 -22131 26512
rect -22258 26432 -22131 26448
rect -22258 26368 -22211 26432
rect -22147 26368 -22131 26432
rect -22258 26352 -22131 26368
rect -22258 26288 -22211 26352
rect -22147 26288 -22131 26352
rect -22258 26272 -22131 26288
rect -22258 26208 -22211 26272
rect -22147 26208 -22131 26272
rect -22258 26192 -22131 26208
rect -22258 26128 -22211 26192
rect -22147 26128 -22131 26192
rect -22258 26112 -22131 26128
rect -22258 26048 -22211 26112
rect -22147 26048 -22131 26112
rect -22258 26032 -22131 26048
rect -22258 25968 -22211 26032
rect -22147 25968 -22131 26032
rect -22258 25952 -22131 25968
rect -22258 25888 -22211 25952
rect -22147 25888 -22131 25952
rect -22258 25872 -22131 25888
rect -22258 25808 -22211 25872
rect -22147 25808 -22131 25872
rect -22258 25792 -22131 25808
rect -22258 25728 -22211 25792
rect -22147 25728 -22131 25792
rect -22258 25712 -22131 25728
rect -22258 25648 -22211 25712
rect -22147 25648 -22131 25712
rect -22258 25632 -22131 25648
rect -22258 25568 -22211 25632
rect -22147 25568 -22131 25632
rect -22258 25552 -22131 25568
rect -22258 25488 -22211 25552
rect -22147 25488 -22131 25552
rect -22258 25472 -22131 25488
rect -22258 25408 -22211 25472
rect -22147 25408 -22131 25472
rect -22258 25392 -22131 25408
rect -22258 25328 -22211 25392
rect -22147 25328 -22131 25392
rect -22258 25312 -22131 25328
rect -22258 25248 -22211 25312
rect -22147 25248 -22131 25312
rect -22258 25232 -22131 25248
rect -22258 25168 -22211 25232
rect -22147 25168 -22131 25232
rect -22258 25152 -22131 25168
rect -22258 25088 -22211 25152
rect -22147 25088 -22131 25152
rect -22258 25072 -22131 25088
rect -22258 25008 -22211 25072
rect -22147 25008 -22131 25072
rect -22258 24992 -22131 25008
rect -22258 24928 -22211 24992
rect -22147 24928 -22131 24992
rect -22258 24912 -22131 24928
rect -22258 24848 -22211 24912
rect -22147 24848 -22131 24912
rect -22258 24832 -22131 24848
rect -22258 24768 -22211 24832
rect -22147 24768 -22131 24832
rect -22258 24752 -22131 24768
rect -22258 24688 -22211 24752
rect -22147 24688 -22131 24752
rect -22258 24672 -22131 24688
rect -22258 24608 -22211 24672
rect -22147 24608 -22131 24672
rect -22258 24592 -22131 24608
rect -22258 24528 -22211 24592
rect -22147 24528 -22131 24592
rect -22258 24512 -22131 24528
rect -22258 24448 -22211 24512
rect -22147 24448 -22131 24512
rect -22258 24432 -22131 24448
rect -22258 24368 -22211 24432
rect -22147 24368 -22131 24432
rect -22258 24352 -22131 24368
rect -22258 24288 -22211 24352
rect -22147 24288 -22131 24352
rect -22258 24272 -22131 24288
rect -22258 24208 -22211 24272
rect -22147 24208 -22131 24272
rect -22258 24192 -22131 24208
rect -22258 24128 -22211 24192
rect -22147 24128 -22131 24192
rect -22258 24112 -22131 24128
rect -22258 24048 -22211 24112
rect -22147 24048 -22131 24112
rect -22258 24032 -22131 24048
rect -22258 23968 -22211 24032
rect -22147 23968 -22131 24032
rect -22258 23952 -22131 23968
rect -22258 23888 -22211 23952
rect -22147 23888 -22131 23952
rect -22258 23872 -22131 23888
rect -22258 23808 -22211 23872
rect -22147 23808 -22131 23872
rect -22258 23792 -22131 23808
rect -22258 23728 -22211 23792
rect -22147 23728 -22131 23792
rect -22258 23712 -22131 23728
rect -22258 23648 -22211 23712
rect -22147 23648 -22131 23712
rect -22258 23632 -22131 23648
rect -22258 23568 -22211 23632
rect -22147 23568 -22131 23632
rect -22258 23552 -22131 23568
rect -22258 23488 -22211 23552
rect -22147 23488 -22131 23552
rect -22258 23472 -22131 23488
rect -22258 23408 -22211 23472
rect -22147 23408 -22131 23472
rect -22258 23392 -22131 23408
rect -22258 23328 -22211 23392
rect -22147 23328 -22131 23392
rect -22258 23312 -22131 23328
rect -22258 23248 -22211 23312
rect -22147 23248 -22131 23312
rect -22258 23232 -22131 23248
rect -22258 23168 -22211 23232
rect -22147 23168 -22131 23232
rect -22258 23152 -22131 23168
rect -22258 23088 -22211 23152
rect -22147 23088 -22131 23152
rect -22258 23072 -22131 23088
rect -22258 23008 -22211 23072
rect -22147 23008 -22131 23072
rect -22258 22992 -22131 23008
rect -22258 22928 -22211 22992
rect -22147 22928 -22131 22992
rect -22258 22912 -22131 22928
rect -22258 22848 -22211 22912
rect -22147 22848 -22131 22912
rect -22258 22832 -22131 22848
rect -22258 22768 -22211 22832
rect -22147 22768 -22131 22832
rect -22258 22752 -22131 22768
rect -22258 22688 -22211 22752
rect -22147 22688 -22131 22752
rect -22258 22672 -22131 22688
rect -22258 22608 -22211 22672
rect -22147 22608 -22131 22672
rect -22258 22592 -22131 22608
rect -22258 22528 -22211 22592
rect -22147 22528 -22131 22592
rect -22258 22512 -22131 22528
rect -22258 22448 -22211 22512
rect -22147 22448 -22131 22512
rect -22258 22432 -22131 22448
rect -22258 22368 -22211 22432
rect -22147 22368 -22131 22432
rect -22258 22352 -22131 22368
rect -22258 22288 -22211 22352
rect -22147 22288 -22131 22352
rect -22258 22272 -22131 22288
rect -28577 22192 -28450 22208
rect -28577 22128 -28530 22192
rect -28466 22128 -28450 22192
rect -28577 22112 -28450 22128
rect -28577 21988 -28473 22112
rect -28577 21972 -28450 21988
rect -28577 21908 -28530 21972
rect -28466 21908 -28450 21972
rect -28577 21892 -28450 21908
rect -34896 21812 -34769 21828
rect -34896 21748 -34849 21812
rect -34785 21748 -34769 21812
rect -34896 21732 -34769 21748
rect -34896 21668 -34849 21732
rect -34785 21668 -34769 21732
rect -34896 21652 -34769 21668
rect -34896 21588 -34849 21652
rect -34785 21588 -34769 21652
rect -34896 21572 -34769 21588
rect -34896 21508 -34849 21572
rect -34785 21508 -34769 21572
rect -34896 21492 -34769 21508
rect -34896 21428 -34849 21492
rect -34785 21428 -34769 21492
rect -34896 21412 -34769 21428
rect -34896 21348 -34849 21412
rect -34785 21348 -34769 21412
rect -34896 21332 -34769 21348
rect -34896 21268 -34849 21332
rect -34785 21268 -34769 21332
rect -34896 21252 -34769 21268
rect -34896 21188 -34849 21252
rect -34785 21188 -34769 21252
rect -34896 21172 -34769 21188
rect -34896 21108 -34849 21172
rect -34785 21108 -34769 21172
rect -34896 21092 -34769 21108
rect -34896 21028 -34849 21092
rect -34785 21028 -34769 21092
rect -34896 21012 -34769 21028
rect -34896 20948 -34849 21012
rect -34785 20948 -34769 21012
rect -34896 20932 -34769 20948
rect -34896 20868 -34849 20932
rect -34785 20868 -34769 20932
rect -34896 20852 -34769 20868
rect -34896 20788 -34849 20852
rect -34785 20788 -34769 20852
rect -34896 20772 -34769 20788
rect -34896 20708 -34849 20772
rect -34785 20708 -34769 20772
rect -34896 20692 -34769 20708
rect -34896 20628 -34849 20692
rect -34785 20628 -34769 20692
rect -34896 20612 -34769 20628
rect -34896 20548 -34849 20612
rect -34785 20548 -34769 20612
rect -34896 20532 -34769 20548
rect -34896 20468 -34849 20532
rect -34785 20468 -34769 20532
rect -34896 20452 -34769 20468
rect -34896 20388 -34849 20452
rect -34785 20388 -34769 20452
rect -34896 20372 -34769 20388
rect -34896 20308 -34849 20372
rect -34785 20308 -34769 20372
rect -34896 20292 -34769 20308
rect -34896 20228 -34849 20292
rect -34785 20228 -34769 20292
rect -34896 20212 -34769 20228
rect -34896 20148 -34849 20212
rect -34785 20148 -34769 20212
rect -34896 20132 -34769 20148
rect -34896 20068 -34849 20132
rect -34785 20068 -34769 20132
rect -34896 20052 -34769 20068
rect -34896 19988 -34849 20052
rect -34785 19988 -34769 20052
rect -34896 19972 -34769 19988
rect -34896 19908 -34849 19972
rect -34785 19908 -34769 19972
rect -34896 19892 -34769 19908
rect -34896 19828 -34849 19892
rect -34785 19828 -34769 19892
rect -34896 19812 -34769 19828
rect -34896 19748 -34849 19812
rect -34785 19748 -34769 19812
rect -34896 19732 -34769 19748
rect -34896 19668 -34849 19732
rect -34785 19668 -34769 19732
rect -34896 19652 -34769 19668
rect -34896 19588 -34849 19652
rect -34785 19588 -34769 19652
rect -34896 19572 -34769 19588
rect -34896 19508 -34849 19572
rect -34785 19508 -34769 19572
rect -34896 19492 -34769 19508
rect -34896 19428 -34849 19492
rect -34785 19428 -34769 19492
rect -34896 19412 -34769 19428
rect -34896 19348 -34849 19412
rect -34785 19348 -34769 19412
rect -34896 19332 -34769 19348
rect -34896 19268 -34849 19332
rect -34785 19268 -34769 19332
rect -34896 19252 -34769 19268
rect -34896 19188 -34849 19252
rect -34785 19188 -34769 19252
rect -34896 19172 -34769 19188
rect -34896 19108 -34849 19172
rect -34785 19108 -34769 19172
rect -34896 19092 -34769 19108
rect -34896 19028 -34849 19092
rect -34785 19028 -34769 19092
rect -34896 19012 -34769 19028
rect -34896 18948 -34849 19012
rect -34785 18948 -34769 19012
rect -34896 18932 -34769 18948
rect -34896 18868 -34849 18932
rect -34785 18868 -34769 18932
rect -34896 18852 -34769 18868
rect -34896 18788 -34849 18852
rect -34785 18788 -34769 18852
rect -34896 18772 -34769 18788
rect -34896 18708 -34849 18772
rect -34785 18708 -34769 18772
rect -34896 18692 -34769 18708
rect -34896 18628 -34849 18692
rect -34785 18628 -34769 18692
rect -34896 18612 -34769 18628
rect -34896 18548 -34849 18612
rect -34785 18548 -34769 18612
rect -34896 18532 -34769 18548
rect -34896 18468 -34849 18532
rect -34785 18468 -34769 18532
rect -34896 18452 -34769 18468
rect -34896 18388 -34849 18452
rect -34785 18388 -34769 18452
rect -34896 18372 -34769 18388
rect -34896 18308 -34849 18372
rect -34785 18308 -34769 18372
rect -34896 18292 -34769 18308
rect -34896 18228 -34849 18292
rect -34785 18228 -34769 18292
rect -34896 18212 -34769 18228
rect -34896 18148 -34849 18212
rect -34785 18148 -34769 18212
rect -34896 18132 -34769 18148
rect -34896 18068 -34849 18132
rect -34785 18068 -34769 18132
rect -34896 18052 -34769 18068
rect -34896 17988 -34849 18052
rect -34785 17988 -34769 18052
rect -34896 17972 -34769 17988
rect -34896 17908 -34849 17972
rect -34785 17908 -34769 17972
rect -34896 17892 -34769 17908
rect -34896 17828 -34849 17892
rect -34785 17828 -34769 17892
rect -34896 17812 -34769 17828
rect -34896 17748 -34849 17812
rect -34785 17748 -34769 17812
rect -34896 17732 -34769 17748
rect -34896 17668 -34849 17732
rect -34785 17668 -34769 17732
rect -34896 17652 -34769 17668
rect -34896 17588 -34849 17652
rect -34785 17588 -34769 17652
rect -34896 17572 -34769 17588
rect -34896 17508 -34849 17572
rect -34785 17508 -34769 17572
rect -34896 17492 -34769 17508
rect -34896 17428 -34849 17492
rect -34785 17428 -34769 17492
rect -34896 17412 -34769 17428
rect -34896 17348 -34849 17412
rect -34785 17348 -34769 17412
rect -34896 17332 -34769 17348
rect -34896 17268 -34849 17332
rect -34785 17268 -34769 17332
rect -34896 17252 -34769 17268
rect -34896 17188 -34849 17252
rect -34785 17188 -34769 17252
rect -34896 17172 -34769 17188
rect -34896 17108 -34849 17172
rect -34785 17108 -34769 17172
rect -34896 17092 -34769 17108
rect -34896 17028 -34849 17092
rect -34785 17028 -34769 17092
rect -34896 17012 -34769 17028
rect -34896 16948 -34849 17012
rect -34785 16948 -34769 17012
rect -34896 16932 -34769 16948
rect -34896 16868 -34849 16932
rect -34785 16868 -34769 16932
rect -34896 16852 -34769 16868
rect -34896 16788 -34849 16852
rect -34785 16788 -34769 16852
rect -34896 16772 -34769 16788
rect -34896 16708 -34849 16772
rect -34785 16708 -34769 16772
rect -34896 16692 -34769 16708
rect -34896 16628 -34849 16692
rect -34785 16628 -34769 16692
rect -34896 16612 -34769 16628
rect -34896 16548 -34849 16612
rect -34785 16548 -34769 16612
rect -34896 16532 -34769 16548
rect -34896 16468 -34849 16532
rect -34785 16468 -34769 16532
rect -34896 16452 -34769 16468
rect -34896 16388 -34849 16452
rect -34785 16388 -34769 16452
rect -34896 16372 -34769 16388
rect -34896 16308 -34849 16372
rect -34785 16308 -34769 16372
rect -34896 16292 -34769 16308
rect -34896 16228 -34849 16292
rect -34785 16228 -34769 16292
rect -34896 16212 -34769 16228
rect -34896 16148 -34849 16212
rect -34785 16148 -34769 16212
rect -34896 16132 -34769 16148
rect -34896 16068 -34849 16132
rect -34785 16068 -34769 16132
rect -34896 16052 -34769 16068
rect -34896 15988 -34849 16052
rect -34785 15988 -34769 16052
rect -34896 15972 -34769 15988
rect -41215 15892 -41088 15908
rect -41215 15828 -41168 15892
rect -41104 15828 -41088 15892
rect -41215 15812 -41088 15828
rect -41215 15688 -41111 15812
rect -41215 15672 -41088 15688
rect -41215 15608 -41168 15672
rect -41104 15608 -41088 15672
rect -41215 15592 -41088 15608
rect -47244 15552 -41322 15561
rect -47244 9648 -47235 15552
rect -41331 9648 -41322 15552
rect -47244 9639 -41322 9648
rect -41215 15528 -41168 15592
rect -41104 15528 -41088 15592
rect -38016 15561 -37912 15939
rect -34896 15908 -34849 15972
rect -34785 15908 -34769 15972
rect -34606 21852 -28684 21861
rect -34606 15948 -34597 21852
rect -28693 15948 -28684 21852
rect -34606 15939 -28684 15948
rect -28577 21828 -28530 21892
rect -28466 21828 -28450 21892
rect -25378 21861 -25274 22239
rect -22258 22208 -22211 22272
rect -22147 22208 -22131 22272
rect -21968 28152 -16046 28161
rect -21968 22248 -21959 28152
rect -16055 22248 -16046 28152
rect -21968 22239 -16046 22248
rect -15939 28128 -15892 28192
rect -15828 28128 -15812 28192
rect -12740 28161 -12636 28539
rect -9620 28508 -9573 28572
rect -9509 28508 -9493 28572
rect -9330 34452 -3408 34461
rect -9330 28548 -9321 34452
rect -3417 28548 -3408 34452
rect -9330 28539 -3408 28548
rect -3301 34428 -3254 34492
rect -3190 34428 -3174 34492
rect -102 34461 2 34839
rect 3018 34808 3065 34872
rect 3129 34808 3145 34872
rect 3308 40752 9230 40761
rect 3308 34848 3317 40752
rect 9221 34848 9230 40752
rect 3308 34839 9230 34848
rect 9337 40728 9384 40792
rect 9448 40728 9464 40792
rect 12536 40761 12640 41139
rect 15656 41108 15703 41172
rect 15767 41108 15783 41172
rect 15946 47052 21868 47061
rect 15946 41148 15955 47052
rect 21859 41148 21868 47052
rect 15946 41139 21868 41148
rect 21975 47028 22022 47092
rect 22086 47028 22102 47092
rect 25174 47061 25278 47250
rect 28294 47188 28398 47250
rect 28294 47172 28421 47188
rect 28294 47108 28341 47172
rect 28405 47108 28421 47172
rect 28294 47092 28421 47108
rect 21975 47012 22102 47028
rect 21975 46948 22022 47012
rect 22086 46948 22102 47012
rect 21975 46932 22102 46948
rect 21975 46868 22022 46932
rect 22086 46868 22102 46932
rect 21975 46852 22102 46868
rect 21975 46788 22022 46852
rect 22086 46788 22102 46852
rect 21975 46772 22102 46788
rect 21975 46708 22022 46772
rect 22086 46708 22102 46772
rect 21975 46692 22102 46708
rect 21975 46628 22022 46692
rect 22086 46628 22102 46692
rect 21975 46612 22102 46628
rect 21975 46548 22022 46612
rect 22086 46548 22102 46612
rect 21975 46532 22102 46548
rect 21975 46468 22022 46532
rect 22086 46468 22102 46532
rect 21975 46452 22102 46468
rect 21975 46388 22022 46452
rect 22086 46388 22102 46452
rect 21975 46372 22102 46388
rect 21975 46308 22022 46372
rect 22086 46308 22102 46372
rect 21975 46292 22102 46308
rect 21975 46228 22022 46292
rect 22086 46228 22102 46292
rect 21975 46212 22102 46228
rect 21975 46148 22022 46212
rect 22086 46148 22102 46212
rect 21975 46132 22102 46148
rect 21975 46068 22022 46132
rect 22086 46068 22102 46132
rect 21975 46052 22102 46068
rect 21975 45988 22022 46052
rect 22086 45988 22102 46052
rect 21975 45972 22102 45988
rect 21975 45908 22022 45972
rect 22086 45908 22102 45972
rect 21975 45892 22102 45908
rect 21975 45828 22022 45892
rect 22086 45828 22102 45892
rect 21975 45812 22102 45828
rect 21975 45748 22022 45812
rect 22086 45748 22102 45812
rect 21975 45732 22102 45748
rect 21975 45668 22022 45732
rect 22086 45668 22102 45732
rect 21975 45652 22102 45668
rect 21975 45588 22022 45652
rect 22086 45588 22102 45652
rect 21975 45572 22102 45588
rect 21975 45508 22022 45572
rect 22086 45508 22102 45572
rect 21975 45492 22102 45508
rect 21975 45428 22022 45492
rect 22086 45428 22102 45492
rect 21975 45412 22102 45428
rect 21975 45348 22022 45412
rect 22086 45348 22102 45412
rect 21975 45332 22102 45348
rect 21975 45268 22022 45332
rect 22086 45268 22102 45332
rect 21975 45252 22102 45268
rect 21975 45188 22022 45252
rect 22086 45188 22102 45252
rect 21975 45172 22102 45188
rect 21975 45108 22022 45172
rect 22086 45108 22102 45172
rect 21975 45092 22102 45108
rect 21975 45028 22022 45092
rect 22086 45028 22102 45092
rect 21975 45012 22102 45028
rect 21975 44948 22022 45012
rect 22086 44948 22102 45012
rect 21975 44932 22102 44948
rect 21975 44868 22022 44932
rect 22086 44868 22102 44932
rect 21975 44852 22102 44868
rect 21975 44788 22022 44852
rect 22086 44788 22102 44852
rect 21975 44772 22102 44788
rect 21975 44708 22022 44772
rect 22086 44708 22102 44772
rect 21975 44692 22102 44708
rect 21975 44628 22022 44692
rect 22086 44628 22102 44692
rect 21975 44612 22102 44628
rect 21975 44548 22022 44612
rect 22086 44548 22102 44612
rect 21975 44532 22102 44548
rect 21975 44468 22022 44532
rect 22086 44468 22102 44532
rect 21975 44452 22102 44468
rect 21975 44388 22022 44452
rect 22086 44388 22102 44452
rect 21975 44372 22102 44388
rect 21975 44308 22022 44372
rect 22086 44308 22102 44372
rect 21975 44292 22102 44308
rect 21975 44228 22022 44292
rect 22086 44228 22102 44292
rect 21975 44212 22102 44228
rect 21975 44148 22022 44212
rect 22086 44148 22102 44212
rect 21975 44132 22102 44148
rect 21975 44068 22022 44132
rect 22086 44068 22102 44132
rect 21975 44052 22102 44068
rect 21975 43988 22022 44052
rect 22086 43988 22102 44052
rect 21975 43972 22102 43988
rect 21975 43908 22022 43972
rect 22086 43908 22102 43972
rect 21975 43892 22102 43908
rect 21975 43828 22022 43892
rect 22086 43828 22102 43892
rect 21975 43812 22102 43828
rect 21975 43748 22022 43812
rect 22086 43748 22102 43812
rect 21975 43732 22102 43748
rect 21975 43668 22022 43732
rect 22086 43668 22102 43732
rect 21975 43652 22102 43668
rect 21975 43588 22022 43652
rect 22086 43588 22102 43652
rect 21975 43572 22102 43588
rect 21975 43508 22022 43572
rect 22086 43508 22102 43572
rect 21975 43492 22102 43508
rect 21975 43428 22022 43492
rect 22086 43428 22102 43492
rect 21975 43412 22102 43428
rect 21975 43348 22022 43412
rect 22086 43348 22102 43412
rect 21975 43332 22102 43348
rect 21975 43268 22022 43332
rect 22086 43268 22102 43332
rect 21975 43252 22102 43268
rect 21975 43188 22022 43252
rect 22086 43188 22102 43252
rect 21975 43172 22102 43188
rect 21975 43108 22022 43172
rect 22086 43108 22102 43172
rect 21975 43092 22102 43108
rect 21975 43028 22022 43092
rect 22086 43028 22102 43092
rect 21975 43012 22102 43028
rect 21975 42948 22022 43012
rect 22086 42948 22102 43012
rect 21975 42932 22102 42948
rect 21975 42868 22022 42932
rect 22086 42868 22102 42932
rect 21975 42852 22102 42868
rect 21975 42788 22022 42852
rect 22086 42788 22102 42852
rect 21975 42772 22102 42788
rect 21975 42708 22022 42772
rect 22086 42708 22102 42772
rect 21975 42692 22102 42708
rect 21975 42628 22022 42692
rect 22086 42628 22102 42692
rect 21975 42612 22102 42628
rect 21975 42548 22022 42612
rect 22086 42548 22102 42612
rect 21975 42532 22102 42548
rect 21975 42468 22022 42532
rect 22086 42468 22102 42532
rect 21975 42452 22102 42468
rect 21975 42388 22022 42452
rect 22086 42388 22102 42452
rect 21975 42372 22102 42388
rect 21975 42308 22022 42372
rect 22086 42308 22102 42372
rect 21975 42292 22102 42308
rect 21975 42228 22022 42292
rect 22086 42228 22102 42292
rect 21975 42212 22102 42228
rect 21975 42148 22022 42212
rect 22086 42148 22102 42212
rect 21975 42132 22102 42148
rect 21975 42068 22022 42132
rect 22086 42068 22102 42132
rect 21975 42052 22102 42068
rect 21975 41988 22022 42052
rect 22086 41988 22102 42052
rect 21975 41972 22102 41988
rect 21975 41908 22022 41972
rect 22086 41908 22102 41972
rect 21975 41892 22102 41908
rect 21975 41828 22022 41892
rect 22086 41828 22102 41892
rect 21975 41812 22102 41828
rect 21975 41748 22022 41812
rect 22086 41748 22102 41812
rect 21975 41732 22102 41748
rect 21975 41668 22022 41732
rect 22086 41668 22102 41732
rect 21975 41652 22102 41668
rect 21975 41588 22022 41652
rect 22086 41588 22102 41652
rect 21975 41572 22102 41588
rect 21975 41508 22022 41572
rect 22086 41508 22102 41572
rect 21975 41492 22102 41508
rect 21975 41428 22022 41492
rect 22086 41428 22102 41492
rect 21975 41412 22102 41428
rect 21975 41348 22022 41412
rect 22086 41348 22102 41412
rect 21975 41332 22102 41348
rect 21975 41268 22022 41332
rect 22086 41268 22102 41332
rect 21975 41252 22102 41268
rect 21975 41188 22022 41252
rect 22086 41188 22102 41252
rect 21975 41172 22102 41188
rect 15656 41092 15783 41108
rect 15656 41028 15703 41092
rect 15767 41028 15783 41092
rect 15656 41012 15783 41028
rect 15656 40888 15760 41012
rect 15656 40872 15783 40888
rect 15656 40808 15703 40872
rect 15767 40808 15783 40872
rect 15656 40792 15783 40808
rect 9337 40712 9464 40728
rect 9337 40648 9384 40712
rect 9448 40648 9464 40712
rect 9337 40632 9464 40648
rect 9337 40568 9384 40632
rect 9448 40568 9464 40632
rect 9337 40552 9464 40568
rect 9337 40488 9384 40552
rect 9448 40488 9464 40552
rect 9337 40472 9464 40488
rect 9337 40408 9384 40472
rect 9448 40408 9464 40472
rect 9337 40392 9464 40408
rect 9337 40328 9384 40392
rect 9448 40328 9464 40392
rect 9337 40312 9464 40328
rect 9337 40248 9384 40312
rect 9448 40248 9464 40312
rect 9337 40232 9464 40248
rect 9337 40168 9384 40232
rect 9448 40168 9464 40232
rect 9337 40152 9464 40168
rect 9337 40088 9384 40152
rect 9448 40088 9464 40152
rect 9337 40072 9464 40088
rect 9337 40008 9384 40072
rect 9448 40008 9464 40072
rect 9337 39992 9464 40008
rect 9337 39928 9384 39992
rect 9448 39928 9464 39992
rect 9337 39912 9464 39928
rect 9337 39848 9384 39912
rect 9448 39848 9464 39912
rect 9337 39832 9464 39848
rect 9337 39768 9384 39832
rect 9448 39768 9464 39832
rect 9337 39752 9464 39768
rect 9337 39688 9384 39752
rect 9448 39688 9464 39752
rect 9337 39672 9464 39688
rect 9337 39608 9384 39672
rect 9448 39608 9464 39672
rect 9337 39592 9464 39608
rect 9337 39528 9384 39592
rect 9448 39528 9464 39592
rect 9337 39512 9464 39528
rect 9337 39448 9384 39512
rect 9448 39448 9464 39512
rect 9337 39432 9464 39448
rect 9337 39368 9384 39432
rect 9448 39368 9464 39432
rect 9337 39352 9464 39368
rect 9337 39288 9384 39352
rect 9448 39288 9464 39352
rect 9337 39272 9464 39288
rect 9337 39208 9384 39272
rect 9448 39208 9464 39272
rect 9337 39192 9464 39208
rect 9337 39128 9384 39192
rect 9448 39128 9464 39192
rect 9337 39112 9464 39128
rect 9337 39048 9384 39112
rect 9448 39048 9464 39112
rect 9337 39032 9464 39048
rect 9337 38968 9384 39032
rect 9448 38968 9464 39032
rect 9337 38952 9464 38968
rect 9337 38888 9384 38952
rect 9448 38888 9464 38952
rect 9337 38872 9464 38888
rect 9337 38808 9384 38872
rect 9448 38808 9464 38872
rect 9337 38792 9464 38808
rect 9337 38728 9384 38792
rect 9448 38728 9464 38792
rect 9337 38712 9464 38728
rect 9337 38648 9384 38712
rect 9448 38648 9464 38712
rect 9337 38632 9464 38648
rect 9337 38568 9384 38632
rect 9448 38568 9464 38632
rect 9337 38552 9464 38568
rect 9337 38488 9384 38552
rect 9448 38488 9464 38552
rect 9337 38472 9464 38488
rect 9337 38408 9384 38472
rect 9448 38408 9464 38472
rect 9337 38392 9464 38408
rect 9337 38328 9384 38392
rect 9448 38328 9464 38392
rect 9337 38312 9464 38328
rect 9337 38248 9384 38312
rect 9448 38248 9464 38312
rect 9337 38232 9464 38248
rect 9337 38168 9384 38232
rect 9448 38168 9464 38232
rect 9337 38152 9464 38168
rect 9337 38088 9384 38152
rect 9448 38088 9464 38152
rect 9337 38072 9464 38088
rect 9337 38008 9384 38072
rect 9448 38008 9464 38072
rect 9337 37992 9464 38008
rect 9337 37928 9384 37992
rect 9448 37928 9464 37992
rect 9337 37912 9464 37928
rect 9337 37848 9384 37912
rect 9448 37848 9464 37912
rect 9337 37832 9464 37848
rect 9337 37768 9384 37832
rect 9448 37768 9464 37832
rect 9337 37752 9464 37768
rect 9337 37688 9384 37752
rect 9448 37688 9464 37752
rect 9337 37672 9464 37688
rect 9337 37608 9384 37672
rect 9448 37608 9464 37672
rect 9337 37592 9464 37608
rect 9337 37528 9384 37592
rect 9448 37528 9464 37592
rect 9337 37512 9464 37528
rect 9337 37448 9384 37512
rect 9448 37448 9464 37512
rect 9337 37432 9464 37448
rect 9337 37368 9384 37432
rect 9448 37368 9464 37432
rect 9337 37352 9464 37368
rect 9337 37288 9384 37352
rect 9448 37288 9464 37352
rect 9337 37272 9464 37288
rect 9337 37208 9384 37272
rect 9448 37208 9464 37272
rect 9337 37192 9464 37208
rect 9337 37128 9384 37192
rect 9448 37128 9464 37192
rect 9337 37112 9464 37128
rect 9337 37048 9384 37112
rect 9448 37048 9464 37112
rect 9337 37032 9464 37048
rect 9337 36968 9384 37032
rect 9448 36968 9464 37032
rect 9337 36952 9464 36968
rect 9337 36888 9384 36952
rect 9448 36888 9464 36952
rect 9337 36872 9464 36888
rect 9337 36808 9384 36872
rect 9448 36808 9464 36872
rect 9337 36792 9464 36808
rect 9337 36728 9384 36792
rect 9448 36728 9464 36792
rect 9337 36712 9464 36728
rect 9337 36648 9384 36712
rect 9448 36648 9464 36712
rect 9337 36632 9464 36648
rect 9337 36568 9384 36632
rect 9448 36568 9464 36632
rect 9337 36552 9464 36568
rect 9337 36488 9384 36552
rect 9448 36488 9464 36552
rect 9337 36472 9464 36488
rect 9337 36408 9384 36472
rect 9448 36408 9464 36472
rect 9337 36392 9464 36408
rect 9337 36328 9384 36392
rect 9448 36328 9464 36392
rect 9337 36312 9464 36328
rect 9337 36248 9384 36312
rect 9448 36248 9464 36312
rect 9337 36232 9464 36248
rect 9337 36168 9384 36232
rect 9448 36168 9464 36232
rect 9337 36152 9464 36168
rect 9337 36088 9384 36152
rect 9448 36088 9464 36152
rect 9337 36072 9464 36088
rect 9337 36008 9384 36072
rect 9448 36008 9464 36072
rect 9337 35992 9464 36008
rect 9337 35928 9384 35992
rect 9448 35928 9464 35992
rect 9337 35912 9464 35928
rect 9337 35848 9384 35912
rect 9448 35848 9464 35912
rect 9337 35832 9464 35848
rect 9337 35768 9384 35832
rect 9448 35768 9464 35832
rect 9337 35752 9464 35768
rect 9337 35688 9384 35752
rect 9448 35688 9464 35752
rect 9337 35672 9464 35688
rect 9337 35608 9384 35672
rect 9448 35608 9464 35672
rect 9337 35592 9464 35608
rect 9337 35528 9384 35592
rect 9448 35528 9464 35592
rect 9337 35512 9464 35528
rect 9337 35448 9384 35512
rect 9448 35448 9464 35512
rect 9337 35432 9464 35448
rect 9337 35368 9384 35432
rect 9448 35368 9464 35432
rect 9337 35352 9464 35368
rect 9337 35288 9384 35352
rect 9448 35288 9464 35352
rect 9337 35272 9464 35288
rect 9337 35208 9384 35272
rect 9448 35208 9464 35272
rect 9337 35192 9464 35208
rect 9337 35128 9384 35192
rect 9448 35128 9464 35192
rect 9337 35112 9464 35128
rect 9337 35048 9384 35112
rect 9448 35048 9464 35112
rect 9337 35032 9464 35048
rect 9337 34968 9384 35032
rect 9448 34968 9464 35032
rect 9337 34952 9464 34968
rect 9337 34888 9384 34952
rect 9448 34888 9464 34952
rect 9337 34872 9464 34888
rect 3018 34792 3145 34808
rect 3018 34728 3065 34792
rect 3129 34728 3145 34792
rect 3018 34712 3145 34728
rect 3018 34588 3122 34712
rect 3018 34572 3145 34588
rect 3018 34508 3065 34572
rect 3129 34508 3145 34572
rect 3018 34492 3145 34508
rect -3301 34412 -3174 34428
rect -3301 34348 -3254 34412
rect -3190 34348 -3174 34412
rect -3301 34332 -3174 34348
rect -3301 34268 -3254 34332
rect -3190 34268 -3174 34332
rect -3301 34252 -3174 34268
rect -3301 34188 -3254 34252
rect -3190 34188 -3174 34252
rect -3301 34172 -3174 34188
rect -3301 34108 -3254 34172
rect -3190 34108 -3174 34172
rect -3301 34092 -3174 34108
rect -3301 34028 -3254 34092
rect -3190 34028 -3174 34092
rect -3301 34012 -3174 34028
rect -3301 33948 -3254 34012
rect -3190 33948 -3174 34012
rect -3301 33932 -3174 33948
rect -3301 33868 -3254 33932
rect -3190 33868 -3174 33932
rect -3301 33852 -3174 33868
rect -3301 33788 -3254 33852
rect -3190 33788 -3174 33852
rect -3301 33772 -3174 33788
rect -3301 33708 -3254 33772
rect -3190 33708 -3174 33772
rect -3301 33692 -3174 33708
rect -3301 33628 -3254 33692
rect -3190 33628 -3174 33692
rect -3301 33612 -3174 33628
rect -3301 33548 -3254 33612
rect -3190 33548 -3174 33612
rect -3301 33532 -3174 33548
rect -3301 33468 -3254 33532
rect -3190 33468 -3174 33532
rect -3301 33452 -3174 33468
rect -3301 33388 -3254 33452
rect -3190 33388 -3174 33452
rect -3301 33372 -3174 33388
rect -3301 33308 -3254 33372
rect -3190 33308 -3174 33372
rect -3301 33292 -3174 33308
rect -3301 33228 -3254 33292
rect -3190 33228 -3174 33292
rect -3301 33212 -3174 33228
rect -3301 33148 -3254 33212
rect -3190 33148 -3174 33212
rect -3301 33132 -3174 33148
rect -3301 33068 -3254 33132
rect -3190 33068 -3174 33132
rect -3301 33052 -3174 33068
rect -3301 32988 -3254 33052
rect -3190 32988 -3174 33052
rect -3301 32972 -3174 32988
rect -3301 32908 -3254 32972
rect -3190 32908 -3174 32972
rect -3301 32892 -3174 32908
rect -3301 32828 -3254 32892
rect -3190 32828 -3174 32892
rect -3301 32812 -3174 32828
rect -3301 32748 -3254 32812
rect -3190 32748 -3174 32812
rect -3301 32732 -3174 32748
rect -3301 32668 -3254 32732
rect -3190 32668 -3174 32732
rect -3301 32652 -3174 32668
rect -3301 32588 -3254 32652
rect -3190 32588 -3174 32652
rect -3301 32572 -3174 32588
rect -3301 32508 -3254 32572
rect -3190 32508 -3174 32572
rect -3301 32492 -3174 32508
rect -3301 32428 -3254 32492
rect -3190 32428 -3174 32492
rect -3301 32412 -3174 32428
rect -3301 32348 -3254 32412
rect -3190 32348 -3174 32412
rect -3301 32332 -3174 32348
rect -3301 32268 -3254 32332
rect -3190 32268 -3174 32332
rect -3301 32252 -3174 32268
rect -3301 32188 -3254 32252
rect -3190 32188 -3174 32252
rect -3301 32172 -3174 32188
rect -3301 32108 -3254 32172
rect -3190 32108 -3174 32172
rect -3301 32092 -3174 32108
rect -3301 32028 -3254 32092
rect -3190 32028 -3174 32092
rect -3301 32012 -3174 32028
rect -3301 31948 -3254 32012
rect -3190 31948 -3174 32012
rect -3301 31932 -3174 31948
rect -3301 31868 -3254 31932
rect -3190 31868 -3174 31932
rect -3301 31852 -3174 31868
rect -3301 31788 -3254 31852
rect -3190 31788 -3174 31852
rect -3301 31772 -3174 31788
rect -3301 31708 -3254 31772
rect -3190 31708 -3174 31772
rect -3301 31692 -3174 31708
rect -3301 31628 -3254 31692
rect -3190 31628 -3174 31692
rect -3301 31612 -3174 31628
rect -3301 31548 -3254 31612
rect -3190 31548 -3174 31612
rect -3301 31532 -3174 31548
rect -3301 31468 -3254 31532
rect -3190 31468 -3174 31532
rect -3301 31452 -3174 31468
rect -3301 31388 -3254 31452
rect -3190 31388 -3174 31452
rect -3301 31372 -3174 31388
rect -3301 31308 -3254 31372
rect -3190 31308 -3174 31372
rect -3301 31292 -3174 31308
rect -3301 31228 -3254 31292
rect -3190 31228 -3174 31292
rect -3301 31212 -3174 31228
rect -3301 31148 -3254 31212
rect -3190 31148 -3174 31212
rect -3301 31132 -3174 31148
rect -3301 31068 -3254 31132
rect -3190 31068 -3174 31132
rect -3301 31052 -3174 31068
rect -3301 30988 -3254 31052
rect -3190 30988 -3174 31052
rect -3301 30972 -3174 30988
rect -3301 30908 -3254 30972
rect -3190 30908 -3174 30972
rect -3301 30892 -3174 30908
rect -3301 30828 -3254 30892
rect -3190 30828 -3174 30892
rect -3301 30812 -3174 30828
rect -3301 30748 -3254 30812
rect -3190 30748 -3174 30812
rect -3301 30732 -3174 30748
rect -3301 30668 -3254 30732
rect -3190 30668 -3174 30732
rect -3301 30652 -3174 30668
rect -3301 30588 -3254 30652
rect -3190 30588 -3174 30652
rect -3301 30572 -3174 30588
rect -3301 30508 -3254 30572
rect -3190 30508 -3174 30572
rect -3301 30492 -3174 30508
rect -3301 30428 -3254 30492
rect -3190 30428 -3174 30492
rect -3301 30412 -3174 30428
rect -3301 30348 -3254 30412
rect -3190 30348 -3174 30412
rect -3301 30332 -3174 30348
rect -3301 30268 -3254 30332
rect -3190 30268 -3174 30332
rect -3301 30252 -3174 30268
rect -3301 30188 -3254 30252
rect -3190 30188 -3174 30252
rect -3301 30172 -3174 30188
rect -3301 30108 -3254 30172
rect -3190 30108 -3174 30172
rect -3301 30092 -3174 30108
rect -3301 30028 -3254 30092
rect -3190 30028 -3174 30092
rect -3301 30012 -3174 30028
rect -3301 29948 -3254 30012
rect -3190 29948 -3174 30012
rect -3301 29932 -3174 29948
rect -3301 29868 -3254 29932
rect -3190 29868 -3174 29932
rect -3301 29852 -3174 29868
rect -3301 29788 -3254 29852
rect -3190 29788 -3174 29852
rect -3301 29772 -3174 29788
rect -3301 29708 -3254 29772
rect -3190 29708 -3174 29772
rect -3301 29692 -3174 29708
rect -3301 29628 -3254 29692
rect -3190 29628 -3174 29692
rect -3301 29612 -3174 29628
rect -3301 29548 -3254 29612
rect -3190 29548 -3174 29612
rect -3301 29532 -3174 29548
rect -3301 29468 -3254 29532
rect -3190 29468 -3174 29532
rect -3301 29452 -3174 29468
rect -3301 29388 -3254 29452
rect -3190 29388 -3174 29452
rect -3301 29372 -3174 29388
rect -3301 29308 -3254 29372
rect -3190 29308 -3174 29372
rect -3301 29292 -3174 29308
rect -3301 29228 -3254 29292
rect -3190 29228 -3174 29292
rect -3301 29212 -3174 29228
rect -3301 29148 -3254 29212
rect -3190 29148 -3174 29212
rect -3301 29132 -3174 29148
rect -3301 29068 -3254 29132
rect -3190 29068 -3174 29132
rect -3301 29052 -3174 29068
rect -3301 28988 -3254 29052
rect -3190 28988 -3174 29052
rect -3301 28972 -3174 28988
rect -3301 28908 -3254 28972
rect -3190 28908 -3174 28972
rect -3301 28892 -3174 28908
rect -3301 28828 -3254 28892
rect -3190 28828 -3174 28892
rect -3301 28812 -3174 28828
rect -3301 28748 -3254 28812
rect -3190 28748 -3174 28812
rect -3301 28732 -3174 28748
rect -3301 28668 -3254 28732
rect -3190 28668 -3174 28732
rect -3301 28652 -3174 28668
rect -3301 28588 -3254 28652
rect -3190 28588 -3174 28652
rect -3301 28572 -3174 28588
rect -9620 28492 -9493 28508
rect -9620 28428 -9573 28492
rect -9509 28428 -9493 28492
rect -9620 28412 -9493 28428
rect -9620 28288 -9516 28412
rect -9620 28272 -9493 28288
rect -9620 28208 -9573 28272
rect -9509 28208 -9493 28272
rect -9620 28192 -9493 28208
rect -15939 28112 -15812 28128
rect -15939 28048 -15892 28112
rect -15828 28048 -15812 28112
rect -15939 28032 -15812 28048
rect -15939 27968 -15892 28032
rect -15828 27968 -15812 28032
rect -15939 27952 -15812 27968
rect -15939 27888 -15892 27952
rect -15828 27888 -15812 27952
rect -15939 27872 -15812 27888
rect -15939 27808 -15892 27872
rect -15828 27808 -15812 27872
rect -15939 27792 -15812 27808
rect -15939 27728 -15892 27792
rect -15828 27728 -15812 27792
rect -15939 27712 -15812 27728
rect -15939 27648 -15892 27712
rect -15828 27648 -15812 27712
rect -15939 27632 -15812 27648
rect -15939 27568 -15892 27632
rect -15828 27568 -15812 27632
rect -15939 27552 -15812 27568
rect -15939 27488 -15892 27552
rect -15828 27488 -15812 27552
rect -15939 27472 -15812 27488
rect -15939 27408 -15892 27472
rect -15828 27408 -15812 27472
rect -15939 27392 -15812 27408
rect -15939 27328 -15892 27392
rect -15828 27328 -15812 27392
rect -15939 27312 -15812 27328
rect -15939 27248 -15892 27312
rect -15828 27248 -15812 27312
rect -15939 27232 -15812 27248
rect -15939 27168 -15892 27232
rect -15828 27168 -15812 27232
rect -15939 27152 -15812 27168
rect -15939 27088 -15892 27152
rect -15828 27088 -15812 27152
rect -15939 27072 -15812 27088
rect -15939 27008 -15892 27072
rect -15828 27008 -15812 27072
rect -15939 26992 -15812 27008
rect -15939 26928 -15892 26992
rect -15828 26928 -15812 26992
rect -15939 26912 -15812 26928
rect -15939 26848 -15892 26912
rect -15828 26848 -15812 26912
rect -15939 26832 -15812 26848
rect -15939 26768 -15892 26832
rect -15828 26768 -15812 26832
rect -15939 26752 -15812 26768
rect -15939 26688 -15892 26752
rect -15828 26688 -15812 26752
rect -15939 26672 -15812 26688
rect -15939 26608 -15892 26672
rect -15828 26608 -15812 26672
rect -15939 26592 -15812 26608
rect -15939 26528 -15892 26592
rect -15828 26528 -15812 26592
rect -15939 26512 -15812 26528
rect -15939 26448 -15892 26512
rect -15828 26448 -15812 26512
rect -15939 26432 -15812 26448
rect -15939 26368 -15892 26432
rect -15828 26368 -15812 26432
rect -15939 26352 -15812 26368
rect -15939 26288 -15892 26352
rect -15828 26288 -15812 26352
rect -15939 26272 -15812 26288
rect -15939 26208 -15892 26272
rect -15828 26208 -15812 26272
rect -15939 26192 -15812 26208
rect -15939 26128 -15892 26192
rect -15828 26128 -15812 26192
rect -15939 26112 -15812 26128
rect -15939 26048 -15892 26112
rect -15828 26048 -15812 26112
rect -15939 26032 -15812 26048
rect -15939 25968 -15892 26032
rect -15828 25968 -15812 26032
rect -15939 25952 -15812 25968
rect -15939 25888 -15892 25952
rect -15828 25888 -15812 25952
rect -15939 25872 -15812 25888
rect -15939 25808 -15892 25872
rect -15828 25808 -15812 25872
rect -15939 25792 -15812 25808
rect -15939 25728 -15892 25792
rect -15828 25728 -15812 25792
rect -15939 25712 -15812 25728
rect -15939 25648 -15892 25712
rect -15828 25648 -15812 25712
rect -15939 25632 -15812 25648
rect -15939 25568 -15892 25632
rect -15828 25568 -15812 25632
rect -15939 25552 -15812 25568
rect -15939 25488 -15892 25552
rect -15828 25488 -15812 25552
rect -15939 25472 -15812 25488
rect -15939 25408 -15892 25472
rect -15828 25408 -15812 25472
rect -15939 25392 -15812 25408
rect -15939 25328 -15892 25392
rect -15828 25328 -15812 25392
rect -15939 25312 -15812 25328
rect -15939 25248 -15892 25312
rect -15828 25248 -15812 25312
rect -15939 25232 -15812 25248
rect -15939 25168 -15892 25232
rect -15828 25168 -15812 25232
rect -15939 25152 -15812 25168
rect -15939 25088 -15892 25152
rect -15828 25088 -15812 25152
rect -15939 25072 -15812 25088
rect -15939 25008 -15892 25072
rect -15828 25008 -15812 25072
rect -15939 24992 -15812 25008
rect -15939 24928 -15892 24992
rect -15828 24928 -15812 24992
rect -15939 24912 -15812 24928
rect -15939 24848 -15892 24912
rect -15828 24848 -15812 24912
rect -15939 24832 -15812 24848
rect -15939 24768 -15892 24832
rect -15828 24768 -15812 24832
rect -15939 24752 -15812 24768
rect -15939 24688 -15892 24752
rect -15828 24688 -15812 24752
rect -15939 24672 -15812 24688
rect -15939 24608 -15892 24672
rect -15828 24608 -15812 24672
rect -15939 24592 -15812 24608
rect -15939 24528 -15892 24592
rect -15828 24528 -15812 24592
rect -15939 24512 -15812 24528
rect -15939 24448 -15892 24512
rect -15828 24448 -15812 24512
rect -15939 24432 -15812 24448
rect -15939 24368 -15892 24432
rect -15828 24368 -15812 24432
rect -15939 24352 -15812 24368
rect -15939 24288 -15892 24352
rect -15828 24288 -15812 24352
rect -15939 24272 -15812 24288
rect -15939 24208 -15892 24272
rect -15828 24208 -15812 24272
rect -15939 24192 -15812 24208
rect -15939 24128 -15892 24192
rect -15828 24128 -15812 24192
rect -15939 24112 -15812 24128
rect -15939 24048 -15892 24112
rect -15828 24048 -15812 24112
rect -15939 24032 -15812 24048
rect -15939 23968 -15892 24032
rect -15828 23968 -15812 24032
rect -15939 23952 -15812 23968
rect -15939 23888 -15892 23952
rect -15828 23888 -15812 23952
rect -15939 23872 -15812 23888
rect -15939 23808 -15892 23872
rect -15828 23808 -15812 23872
rect -15939 23792 -15812 23808
rect -15939 23728 -15892 23792
rect -15828 23728 -15812 23792
rect -15939 23712 -15812 23728
rect -15939 23648 -15892 23712
rect -15828 23648 -15812 23712
rect -15939 23632 -15812 23648
rect -15939 23568 -15892 23632
rect -15828 23568 -15812 23632
rect -15939 23552 -15812 23568
rect -15939 23488 -15892 23552
rect -15828 23488 -15812 23552
rect -15939 23472 -15812 23488
rect -15939 23408 -15892 23472
rect -15828 23408 -15812 23472
rect -15939 23392 -15812 23408
rect -15939 23328 -15892 23392
rect -15828 23328 -15812 23392
rect -15939 23312 -15812 23328
rect -15939 23248 -15892 23312
rect -15828 23248 -15812 23312
rect -15939 23232 -15812 23248
rect -15939 23168 -15892 23232
rect -15828 23168 -15812 23232
rect -15939 23152 -15812 23168
rect -15939 23088 -15892 23152
rect -15828 23088 -15812 23152
rect -15939 23072 -15812 23088
rect -15939 23008 -15892 23072
rect -15828 23008 -15812 23072
rect -15939 22992 -15812 23008
rect -15939 22928 -15892 22992
rect -15828 22928 -15812 22992
rect -15939 22912 -15812 22928
rect -15939 22848 -15892 22912
rect -15828 22848 -15812 22912
rect -15939 22832 -15812 22848
rect -15939 22768 -15892 22832
rect -15828 22768 -15812 22832
rect -15939 22752 -15812 22768
rect -15939 22688 -15892 22752
rect -15828 22688 -15812 22752
rect -15939 22672 -15812 22688
rect -15939 22608 -15892 22672
rect -15828 22608 -15812 22672
rect -15939 22592 -15812 22608
rect -15939 22528 -15892 22592
rect -15828 22528 -15812 22592
rect -15939 22512 -15812 22528
rect -15939 22448 -15892 22512
rect -15828 22448 -15812 22512
rect -15939 22432 -15812 22448
rect -15939 22368 -15892 22432
rect -15828 22368 -15812 22432
rect -15939 22352 -15812 22368
rect -15939 22288 -15892 22352
rect -15828 22288 -15812 22352
rect -15939 22272 -15812 22288
rect -22258 22192 -22131 22208
rect -22258 22128 -22211 22192
rect -22147 22128 -22131 22192
rect -22258 22112 -22131 22128
rect -22258 21988 -22154 22112
rect -22258 21972 -22131 21988
rect -22258 21908 -22211 21972
rect -22147 21908 -22131 21972
rect -22258 21892 -22131 21908
rect -28577 21812 -28450 21828
rect -28577 21748 -28530 21812
rect -28466 21748 -28450 21812
rect -28577 21732 -28450 21748
rect -28577 21668 -28530 21732
rect -28466 21668 -28450 21732
rect -28577 21652 -28450 21668
rect -28577 21588 -28530 21652
rect -28466 21588 -28450 21652
rect -28577 21572 -28450 21588
rect -28577 21508 -28530 21572
rect -28466 21508 -28450 21572
rect -28577 21492 -28450 21508
rect -28577 21428 -28530 21492
rect -28466 21428 -28450 21492
rect -28577 21412 -28450 21428
rect -28577 21348 -28530 21412
rect -28466 21348 -28450 21412
rect -28577 21332 -28450 21348
rect -28577 21268 -28530 21332
rect -28466 21268 -28450 21332
rect -28577 21252 -28450 21268
rect -28577 21188 -28530 21252
rect -28466 21188 -28450 21252
rect -28577 21172 -28450 21188
rect -28577 21108 -28530 21172
rect -28466 21108 -28450 21172
rect -28577 21092 -28450 21108
rect -28577 21028 -28530 21092
rect -28466 21028 -28450 21092
rect -28577 21012 -28450 21028
rect -28577 20948 -28530 21012
rect -28466 20948 -28450 21012
rect -28577 20932 -28450 20948
rect -28577 20868 -28530 20932
rect -28466 20868 -28450 20932
rect -28577 20852 -28450 20868
rect -28577 20788 -28530 20852
rect -28466 20788 -28450 20852
rect -28577 20772 -28450 20788
rect -28577 20708 -28530 20772
rect -28466 20708 -28450 20772
rect -28577 20692 -28450 20708
rect -28577 20628 -28530 20692
rect -28466 20628 -28450 20692
rect -28577 20612 -28450 20628
rect -28577 20548 -28530 20612
rect -28466 20548 -28450 20612
rect -28577 20532 -28450 20548
rect -28577 20468 -28530 20532
rect -28466 20468 -28450 20532
rect -28577 20452 -28450 20468
rect -28577 20388 -28530 20452
rect -28466 20388 -28450 20452
rect -28577 20372 -28450 20388
rect -28577 20308 -28530 20372
rect -28466 20308 -28450 20372
rect -28577 20292 -28450 20308
rect -28577 20228 -28530 20292
rect -28466 20228 -28450 20292
rect -28577 20212 -28450 20228
rect -28577 20148 -28530 20212
rect -28466 20148 -28450 20212
rect -28577 20132 -28450 20148
rect -28577 20068 -28530 20132
rect -28466 20068 -28450 20132
rect -28577 20052 -28450 20068
rect -28577 19988 -28530 20052
rect -28466 19988 -28450 20052
rect -28577 19972 -28450 19988
rect -28577 19908 -28530 19972
rect -28466 19908 -28450 19972
rect -28577 19892 -28450 19908
rect -28577 19828 -28530 19892
rect -28466 19828 -28450 19892
rect -28577 19812 -28450 19828
rect -28577 19748 -28530 19812
rect -28466 19748 -28450 19812
rect -28577 19732 -28450 19748
rect -28577 19668 -28530 19732
rect -28466 19668 -28450 19732
rect -28577 19652 -28450 19668
rect -28577 19588 -28530 19652
rect -28466 19588 -28450 19652
rect -28577 19572 -28450 19588
rect -28577 19508 -28530 19572
rect -28466 19508 -28450 19572
rect -28577 19492 -28450 19508
rect -28577 19428 -28530 19492
rect -28466 19428 -28450 19492
rect -28577 19412 -28450 19428
rect -28577 19348 -28530 19412
rect -28466 19348 -28450 19412
rect -28577 19332 -28450 19348
rect -28577 19268 -28530 19332
rect -28466 19268 -28450 19332
rect -28577 19252 -28450 19268
rect -28577 19188 -28530 19252
rect -28466 19188 -28450 19252
rect -28577 19172 -28450 19188
rect -28577 19108 -28530 19172
rect -28466 19108 -28450 19172
rect -28577 19092 -28450 19108
rect -28577 19028 -28530 19092
rect -28466 19028 -28450 19092
rect -28577 19012 -28450 19028
rect -28577 18948 -28530 19012
rect -28466 18948 -28450 19012
rect -28577 18932 -28450 18948
rect -28577 18868 -28530 18932
rect -28466 18868 -28450 18932
rect -28577 18852 -28450 18868
rect -28577 18788 -28530 18852
rect -28466 18788 -28450 18852
rect -28577 18772 -28450 18788
rect -28577 18708 -28530 18772
rect -28466 18708 -28450 18772
rect -28577 18692 -28450 18708
rect -28577 18628 -28530 18692
rect -28466 18628 -28450 18692
rect -28577 18612 -28450 18628
rect -28577 18548 -28530 18612
rect -28466 18548 -28450 18612
rect -28577 18532 -28450 18548
rect -28577 18468 -28530 18532
rect -28466 18468 -28450 18532
rect -28577 18452 -28450 18468
rect -28577 18388 -28530 18452
rect -28466 18388 -28450 18452
rect -28577 18372 -28450 18388
rect -28577 18308 -28530 18372
rect -28466 18308 -28450 18372
rect -28577 18292 -28450 18308
rect -28577 18228 -28530 18292
rect -28466 18228 -28450 18292
rect -28577 18212 -28450 18228
rect -28577 18148 -28530 18212
rect -28466 18148 -28450 18212
rect -28577 18132 -28450 18148
rect -28577 18068 -28530 18132
rect -28466 18068 -28450 18132
rect -28577 18052 -28450 18068
rect -28577 17988 -28530 18052
rect -28466 17988 -28450 18052
rect -28577 17972 -28450 17988
rect -28577 17908 -28530 17972
rect -28466 17908 -28450 17972
rect -28577 17892 -28450 17908
rect -28577 17828 -28530 17892
rect -28466 17828 -28450 17892
rect -28577 17812 -28450 17828
rect -28577 17748 -28530 17812
rect -28466 17748 -28450 17812
rect -28577 17732 -28450 17748
rect -28577 17668 -28530 17732
rect -28466 17668 -28450 17732
rect -28577 17652 -28450 17668
rect -28577 17588 -28530 17652
rect -28466 17588 -28450 17652
rect -28577 17572 -28450 17588
rect -28577 17508 -28530 17572
rect -28466 17508 -28450 17572
rect -28577 17492 -28450 17508
rect -28577 17428 -28530 17492
rect -28466 17428 -28450 17492
rect -28577 17412 -28450 17428
rect -28577 17348 -28530 17412
rect -28466 17348 -28450 17412
rect -28577 17332 -28450 17348
rect -28577 17268 -28530 17332
rect -28466 17268 -28450 17332
rect -28577 17252 -28450 17268
rect -28577 17188 -28530 17252
rect -28466 17188 -28450 17252
rect -28577 17172 -28450 17188
rect -28577 17108 -28530 17172
rect -28466 17108 -28450 17172
rect -28577 17092 -28450 17108
rect -28577 17028 -28530 17092
rect -28466 17028 -28450 17092
rect -28577 17012 -28450 17028
rect -28577 16948 -28530 17012
rect -28466 16948 -28450 17012
rect -28577 16932 -28450 16948
rect -28577 16868 -28530 16932
rect -28466 16868 -28450 16932
rect -28577 16852 -28450 16868
rect -28577 16788 -28530 16852
rect -28466 16788 -28450 16852
rect -28577 16772 -28450 16788
rect -28577 16708 -28530 16772
rect -28466 16708 -28450 16772
rect -28577 16692 -28450 16708
rect -28577 16628 -28530 16692
rect -28466 16628 -28450 16692
rect -28577 16612 -28450 16628
rect -28577 16548 -28530 16612
rect -28466 16548 -28450 16612
rect -28577 16532 -28450 16548
rect -28577 16468 -28530 16532
rect -28466 16468 -28450 16532
rect -28577 16452 -28450 16468
rect -28577 16388 -28530 16452
rect -28466 16388 -28450 16452
rect -28577 16372 -28450 16388
rect -28577 16308 -28530 16372
rect -28466 16308 -28450 16372
rect -28577 16292 -28450 16308
rect -28577 16228 -28530 16292
rect -28466 16228 -28450 16292
rect -28577 16212 -28450 16228
rect -28577 16148 -28530 16212
rect -28466 16148 -28450 16212
rect -28577 16132 -28450 16148
rect -28577 16068 -28530 16132
rect -28466 16068 -28450 16132
rect -28577 16052 -28450 16068
rect -28577 15988 -28530 16052
rect -28466 15988 -28450 16052
rect -28577 15972 -28450 15988
rect -34896 15892 -34769 15908
rect -34896 15828 -34849 15892
rect -34785 15828 -34769 15892
rect -34896 15812 -34769 15828
rect -34896 15688 -34792 15812
rect -34896 15672 -34769 15688
rect -34896 15608 -34849 15672
rect -34785 15608 -34769 15672
rect -34896 15592 -34769 15608
rect -41215 15512 -41088 15528
rect -41215 15448 -41168 15512
rect -41104 15448 -41088 15512
rect -41215 15432 -41088 15448
rect -41215 15368 -41168 15432
rect -41104 15368 -41088 15432
rect -41215 15352 -41088 15368
rect -41215 15288 -41168 15352
rect -41104 15288 -41088 15352
rect -41215 15272 -41088 15288
rect -41215 15208 -41168 15272
rect -41104 15208 -41088 15272
rect -41215 15192 -41088 15208
rect -41215 15128 -41168 15192
rect -41104 15128 -41088 15192
rect -41215 15112 -41088 15128
rect -41215 15048 -41168 15112
rect -41104 15048 -41088 15112
rect -41215 15032 -41088 15048
rect -41215 14968 -41168 15032
rect -41104 14968 -41088 15032
rect -41215 14952 -41088 14968
rect -41215 14888 -41168 14952
rect -41104 14888 -41088 14952
rect -41215 14872 -41088 14888
rect -41215 14808 -41168 14872
rect -41104 14808 -41088 14872
rect -41215 14792 -41088 14808
rect -41215 14728 -41168 14792
rect -41104 14728 -41088 14792
rect -41215 14712 -41088 14728
rect -41215 14648 -41168 14712
rect -41104 14648 -41088 14712
rect -41215 14632 -41088 14648
rect -41215 14568 -41168 14632
rect -41104 14568 -41088 14632
rect -41215 14552 -41088 14568
rect -41215 14488 -41168 14552
rect -41104 14488 -41088 14552
rect -41215 14472 -41088 14488
rect -41215 14408 -41168 14472
rect -41104 14408 -41088 14472
rect -41215 14392 -41088 14408
rect -41215 14328 -41168 14392
rect -41104 14328 -41088 14392
rect -41215 14312 -41088 14328
rect -41215 14248 -41168 14312
rect -41104 14248 -41088 14312
rect -41215 14232 -41088 14248
rect -41215 14168 -41168 14232
rect -41104 14168 -41088 14232
rect -41215 14152 -41088 14168
rect -41215 14088 -41168 14152
rect -41104 14088 -41088 14152
rect -41215 14072 -41088 14088
rect -41215 14008 -41168 14072
rect -41104 14008 -41088 14072
rect -41215 13992 -41088 14008
rect -41215 13928 -41168 13992
rect -41104 13928 -41088 13992
rect -41215 13912 -41088 13928
rect -41215 13848 -41168 13912
rect -41104 13848 -41088 13912
rect -41215 13832 -41088 13848
rect -41215 13768 -41168 13832
rect -41104 13768 -41088 13832
rect -41215 13752 -41088 13768
rect -41215 13688 -41168 13752
rect -41104 13688 -41088 13752
rect -41215 13672 -41088 13688
rect -41215 13608 -41168 13672
rect -41104 13608 -41088 13672
rect -41215 13592 -41088 13608
rect -41215 13528 -41168 13592
rect -41104 13528 -41088 13592
rect -41215 13512 -41088 13528
rect -41215 13448 -41168 13512
rect -41104 13448 -41088 13512
rect -41215 13432 -41088 13448
rect -41215 13368 -41168 13432
rect -41104 13368 -41088 13432
rect -41215 13352 -41088 13368
rect -41215 13288 -41168 13352
rect -41104 13288 -41088 13352
rect -41215 13272 -41088 13288
rect -41215 13208 -41168 13272
rect -41104 13208 -41088 13272
rect -41215 13192 -41088 13208
rect -41215 13128 -41168 13192
rect -41104 13128 -41088 13192
rect -41215 13112 -41088 13128
rect -41215 13048 -41168 13112
rect -41104 13048 -41088 13112
rect -41215 13032 -41088 13048
rect -41215 12968 -41168 13032
rect -41104 12968 -41088 13032
rect -41215 12952 -41088 12968
rect -41215 12888 -41168 12952
rect -41104 12888 -41088 12952
rect -41215 12872 -41088 12888
rect -41215 12808 -41168 12872
rect -41104 12808 -41088 12872
rect -41215 12792 -41088 12808
rect -41215 12728 -41168 12792
rect -41104 12728 -41088 12792
rect -41215 12712 -41088 12728
rect -41215 12648 -41168 12712
rect -41104 12648 -41088 12712
rect -41215 12632 -41088 12648
rect -41215 12568 -41168 12632
rect -41104 12568 -41088 12632
rect -41215 12552 -41088 12568
rect -41215 12488 -41168 12552
rect -41104 12488 -41088 12552
rect -41215 12472 -41088 12488
rect -41215 12408 -41168 12472
rect -41104 12408 -41088 12472
rect -41215 12392 -41088 12408
rect -41215 12328 -41168 12392
rect -41104 12328 -41088 12392
rect -41215 12312 -41088 12328
rect -41215 12248 -41168 12312
rect -41104 12248 -41088 12312
rect -41215 12232 -41088 12248
rect -41215 12168 -41168 12232
rect -41104 12168 -41088 12232
rect -41215 12152 -41088 12168
rect -41215 12088 -41168 12152
rect -41104 12088 -41088 12152
rect -41215 12072 -41088 12088
rect -41215 12008 -41168 12072
rect -41104 12008 -41088 12072
rect -41215 11992 -41088 12008
rect -41215 11928 -41168 11992
rect -41104 11928 -41088 11992
rect -41215 11912 -41088 11928
rect -41215 11848 -41168 11912
rect -41104 11848 -41088 11912
rect -41215 11832 -41088 11848
rect -41215 11768 -41168 11832
rect -41104 11768 -41088 11832
rect -41215 11752 -41088 11768
rect -41215 11688 -41168 11752
rect -41104 11688 -41088 11752
rect -41215 11672 -41088 11688
rect -41215 11608 -41168 11672
rect -41104 11608 -41088 11672
rect -41215 11592 -41088 11608
rect -41215 11528 -41168 11592
rect -41104 11528 -41088 11592
rect -41215 11512 -41088 11528
rect -41215 11448 -41168 11512
rect -41104 11448 -41088 11512
rect -41215 11432 -41088 11448
rect -41215 11368 -41168 11432
rect -41104 11368 -41088 11432
rect -41215 11352 -41088 11368
rect -41215 11288 -41168 11352
rect -41104 11288 -41088 11352
rect -41215 11272 -41088 11288
rect -41215 11208 -41168 11272
rect -41104 11208 -41088 11272
rect -41215 11192 -41088 11208
rect -41215 11128 -41168 11192
rect -41104 11128 -41088 11192
rect -41215 11112 -41088 11128
rect -41215 11048 -41168 11112
rect -41104 11048 -41088 11112
rect -41215 11032 -41088 11048
rect -41215 10968 -41168 11032
rect -41104 10968 -41088 11032
rect -41215 10952 -41088 10968
rect -41215 10888 -41168 10952
rect -41104 10888 -41088 10952
rect -41215 10872 -41088 10888
rect -41215 10808 -41168 10872
rect -41104 10808 -41088 10872
rect -41215 10792 -41088 10808
rect -41215 10728 -41168 10792
rect -41104 10728 -41088 10792
rect -41215 10712 -41088 10728
rect -41215 10648 -41168 10712
rect -41104 10648 -41088 10712
rect -41215 10632 -41088 10648
rect -41215 10568 -41168 10632
rect -41104 10568 -41088 10632
rect -41215 10552 -41088 10568
rect -41215 10488 -41168 10552
rect -41104 10488 -41088 10552
rect -41215 10472 -41088 10488
rect -41215 10408 -41168 10472
rect -41104 10408 -41088 10472
rect -41215 10392 -41088 10408
rect -41215 10328 -41168 10392
rect -41104 10328 -41088 10392
rect -41215 10312 -41088 10328
rect -41215 10248 -41168 10312
rect -41104 10248 -41088 10312
rect -41215 10232 -41088 10248
rect -41215 10168 -41168 10232
rect -41104 10168 -41088 10232
rect -41215 10152 -41088 10168
rect -41215 10088 -41168 10152
rect -41104 10088 -41088 10152
rect -41215 10072 -41088 10088
rect -41215 10008 -41168 10072
rect -41104 10008 -41088 10072
rect -41215 9992 -41088 10008
rect -41215 9928 -41168 9992
rect -41104 9928 -41088 9992
rect -41215 9912 -41088 9928
rect -41215 9848 -41168 9912
rect -41104 9848 -41088 9912
rect -41215 9832 -41088 9848
rect -41215 9768 -41168 9832
rect -41104 9768 -41088 9832
rect -41215 9752 -41088 9768
rect -41215 9688 -41168 9752
rect -41104 9688 -41088 9752
rect -41215 9672 -41088 9688
rect -44335 9261 -44231 9639
rect -41215 9608 -41168 9672
rect -41104 9608 -41088 9672
rect -40925 15552 -35003 15561
rect -40925 9648 -40916 15552
rect -35012 9648 -35003 15552
rect -40925 9639 -35003 9648
rect -34896 15528 -34849 15592
rect -34785 15528 -34769 15592
rect -31697 15561 -31593 15939
rect -28577 15908 -28530 15972
rect -28466 15908 -28450 15972
rect -28287 21852 -22365 21861
rect -28287 15948 -28278 21852
rect -22374 15948 -22365 21852
rect -28287 15939 -22365 15948
rect -22258 21828 -22211 21892
rect -22147 21828 -22131 21892
rect -19059 21861 -18955 22239
rect -15939 22208 -15892 22272
rect -15828 22208 -15812 22272
rect -15649 28152 -9727 28161
rect -15649 22248 -15640 28152
rect -9736 22248 -9727 28152
rect -15649 22239 -9727 22248
rect -9620 28128 -9573 28192
rect -9509 28128 -9493 28192
rect -6421 28161 -6317 28539
rect -3301 28508 -3254 28572
rect -3190 28508 -3174 28572
rect -3011 34452 2911 34461
rect -3011 28548 -3002 34452
rect 2902 28548 2911 34452
rect -3011 28539 2911 28548
rect 3018 34428 3065 34492
rect 3129 34428 3145 34492
rect 6217 34461 6321 34839
rect 9337 34808 9384 34872
rect 9448 34808 9464 34872
rect 9627 40752 15549 40761
rect 9627 34848 9636 40752
rect 15540 34848 15549 40752
rect 9627 34839 15549 34848
rect 15656 40728 15703 40792
rect 15767 40728 15783 40792
rect 18855 40761 18959 41139
rect 21975 41108 22022 41172
rect 22086 41108 22102 41172
rect 22265 47052 28187 47061
rect 22265 41148 22274 47052
rect 28178 41148 28187 47052
rect 22265 41139 28187 41148
rect 28294 47028 28341 47092
rect 28405 47028 28421 47092
rect 31493 47061 31597 47250
rect 34613 47188 34717 47250
rect 34613 47172 34740 47188
rect 34613 47108 34660 47172
rect 34724 47108 34740 47172
rect 34613 47092 34740 47108
rect 28294 47012 28421 47028
rect 28294 46948 28341 47012
rect 28405 46948 28421 47012
rect 28294 46932 28421 46948
rect 28294 46868 28341 46932
rect 28405 46868 28421 46932
rect 28294 46852 28421 46868
rect 28294 46788 28341 46852
rect 28405 46788 28421 46852
rect 28294 46772 28421 46788
rect 28294 46708 28341 46772
rect 28405 46708 28421 46772
rect 28294 46692 28421 46708
rect 28294 46628 28341 46692
rect 28405 46628 28421 46692
rect 28294 46612 28421 46628
rect 28294 46548 28341 46612
rect 28405 46548 28421 46612
rect 28294 46532 28421 46548
rect 28294 46468 28341 46532
rect 28405 46468 28421 46532
rect 28294 46452 28421 46468
rect 28294 46388 28341 46452
rect 28405 46388 28421 46452
rect 28294 46372 28421 46388
rect 28294 46308 28341 46372
rect 28405 46308 28421 46372
rect 28294 46292 28421 46308
rect 28294 46228 28341 46292
rect 28405 46228 28421 46292
rect 28294 46212 28421 46228
rect 28294 46148 28341 46212
rect 28405 46148 28421 46212
rect 28294 46132 28421 46148
rect 28294 46068 28341 46132
rect 28405 46068 28421 46132
rect 28294 46052 28421 46068
rect 28294 45988 28341 46052
rect 28405 45988 28421 46052
rect 28294 45972 28421 45988
rect 28294 45908 28341 45972
rect 28405 45908 28421 45972
rect 28294 45892 28421 45908
rect 28294 45828 28341 45892
rect 28405 45828 28421 45892
rect 28294 45812 28421 45828
rect 28294 45748 28341 45812
rect 28405 45748 28421 45812
rect 28294 45732 28421 45748
rect 28294 45668 28341 45732
rect 28405 45668 28421 45732
rect 28294 45652 28421 45668
rect 28294 45588 28341 45652
rect 28405 45588 28421 45652
rect 28294 45572 28421 45588
rect 28294 45508 28341 45572
rect 28405 45508 28421 45572
rect 28294 45492 28421 45508
rect 28294 45428 28341 45492
rect 28405 45428 28421 45492
rect 28294 45412 28421 45428
rect 28294 45348 28341 45412
rect 28405 45348 28421 45412
rect 28294 45332 28421 45348
rect 28294 45268 28341 45332
rect 28405 45268 28421 45332
rect 28294 45252 28421 45268
rect 28294 45188 28341 45252
rect 28405 45188 28421 45252
rect 28294 45172 28421 45188
rect 28294 45108 28341 45172
rect 28405 45108 28421 45172
rect 28294 45092 28421 45108
rect 28294 45028 28341 45092
rect 28405 45028 28421 45092
rect 28294 45012 28421 45028
rect 28294 44948 28341 45012
rect 28405 44948 28421 45012
rect 28294 44932 28421 44948
rect 28294 44868 28341 44932
rect 28405 44868 28421 44932
rect 28294 44852 28421 44868
rect 28294 44788 28341 44852
rect 28405 44788 28421 44852
rect 28294 44772 28421 44788
rect 28294 44708 28341 44772
rect 28405 44708 28421 44772
rect 28294 44692 28421 44708
rect 28294 44628 28341 44692
rect 28405 44628 28421 44692
rect 28294 44612 28421 44628
rect 28294 44548 28341 44612
rect 28405 44548 28421 44612
rect 28294 44532 28421 44548
rect 28294 44468 28341 44532
rect 28405 44468 28421 44532
rect 28294 44452 28421 44468
rect 28294 44388 28341 44452
rect 28405 44388 28421 44452
rect 28294 44372 28421 44388
rect 28294 44308 28341 44372
rect 28405 44308 28421 44372
rect 28294 44292 28421 44308
rect 28294 44228 28341 44292
rect 28405 44228 28421 44292
rect 28294 44212 28421 44228
rect 28294 44148 28341 44212
rect 28405 44148 28421 44212
rect 28294 44132 28421 44148
rect 28294 44068 28341 44132
rect 28405 44068 28421 44132
rect 28294 44052 28421 44068
rect 28294 43988 28341 44052
rect 28405 43988 28421 44052
rect 28294 43972 28421 43988
rect 28294 43908 28341 43972
rect 28405 43908 28421 43972
rect 28294 43892 28421 43908
rect 28294 43828 28341 43892
rect 28405 43828 28421 43892
rect 28294 43812 28421 43828
rect 28294 43748 28341 43812
rect 28405 43748 28421 43812
rect 28294 43732 28421 43748
rect 28294 43668 28341 43732
rect 28405 43668 28421 43732
rect 28294 43652 28421 43668
rect 28294 43588 28341 43652
rect 28405 43588 28421 43652
rect 28294 43572 28421 43588
rect 28294 43508 28341 43572
rect 28405 43508 28421 43572
rect 28294 43492 28421 43508
rect 28294 43428 28341 43492
rect 28405 43428 28421 43492
rect 28294 43412 28421 43428
rect 28294 43348 28341 43412
rect 28405 43348 28421 43412
rect 28294 43332 28421 43348
rect 28294 43268 28341 43332
rect 28405 43268 28421 43332
rect 28294 43252 28421 43268
rect 28294 43188 28341 43252
rect 28405 43188 28421 43252
rect 28294 43172 28421 43188
rect 28294 43108 28341 43172
rect 28405 43108 28421 43172
rect 28294 43092 28421 43108
rect 28294 43028 28341 43092
rect 28405 43028 28421 43092
rect 28294 43012 28421 43028
rect 28294 42948 28341 43012
rect 28405 42948 28421 43012
rect 28294 42932 28421 42948
rect 28294 42868 28341 42932
rect 28405 42868 28421 42932
rect 28294 42852 28421 42868
rect 28294 42788 28341 42852
rect 28405 42788 28421 42852
rect 28294 42772 28421 42788
rect 28294 42708 28341 42772
rect 28405 42708 28421 42772
rect 28294 42692 28421 42708
rect 28294 42628 28341 42692
rect 28405 42628 28421 42692
rect 28294 42612 28421 42628
rect 28294 42548 28341 42612
rect 28405 42548 28421 42612
rect 28294 42532 28421 42548
rect 28294 42468 28341 42532
rect 28405 42468 28421 42532
rect 28294 42452 28421 42468
rect 28294 42388 28341 42452
rect 28405 42388 28421 42452
rect 28294 42372 28421 42388
rect 28294 42308 28341 42372
rect 28405 42308 28421 42372
rect 28294 42292 28421 42308
rect 28294 42228 28341 42292
rect 28405 42228 28421 42292
rect 28294 42212 28421 42228
rect 28294 42148 28341 42212
rect 28405 42148 28421 42212
rect 28294 42132 28421 42148
rect 28294 42068 28341 42132
rect 28405 42068 28421 42132
rect 28294 42052 28421 42068
rect 28294 41988 28341 42052
rect 28405 41988 28421 42052
rect 28294 41972 28421 41988
rect 28294 41908 28341 41972
rect 28405 41908 28421 41972
rect 28294 41892 28421 41908
rect 28294 41828 28341 41892
rect 28405 41828 28421 41892
rect 28294 41812 28421 41828
rect 28294 41748 28341 41812
rect 28405 41748 28421 41812
rect 28294 41732 28421 41748
rect 28294 41668 28341 41732
rect 28405 41668 28421 41732
rect 28294 41652 28421 41668
rect 28294 41588 28341 41652
rect 28405 41588 28421 41652
rect 28294 41572 28421 41588
rect 28294 41508 28341 41572
rect 28405 41508 28421 41572
rect 28294 41492 28421 41508
rect 28294 41428 28341 41492
rect 28405 41428 28421 41492
rect 28294 41412 28421 41428
rect 28294 41348 28341 41412
rect 28405 41348 28421 41412
rect 28294 41332 28421 41348
rect 28294 41268 28341 41332
rect 28405 41268 28421 41332
rect 28294 41252 28421 41268
rect 28294 41188 28341 41252
rect 28405 41188 28421 41252
rect 28294 41172 28421 41188
rect 21975 41092 22102 41108
rect 21975 41028 22022 41092
rect 22086 41028 22102 41092
rect 21975 41012 22102 41028
rect 21975 40888 22079 41012
rect 21975 40872 22102 40888
rect 21975 40808 22022 40872
rect 22086 40808 22102 40872
rect 21975 40792 22102 40808
rect 15656 40712 15783 40728
rect 15656 40648 15703 40712
rect 15767 40648 15783 40712
rect 15656 40632 15783 40648
rect 15656 40568 15703 40632
rect 15767 40568 15783 40632
rect 15656 40552 15783 40568
rect 15656 40488 15703 40552
rect 15767 40488 15783 40552
rect 15656 40472 15783 40488
rect 15656 40408 15703 40472
rect 15767 40408 15783 40472
rect 15656 40392 15783 40408
rect 15656 40328 15703 40392
rect 15767 40328 15783 40392
rect 15656 40312 15783 40328
rect 15656 40248 15703 40312
rect 15767 40248 15783 40312
rect 15656 40232 15783 40248
rect 15656 40168 15703 40232
rect 15767 40168 15783 40232
rect 15656 40152 15783 40168
rect 15656 40088 15703 40152
rect 15767 40088 15783 40152
rect 15656 40072 15783 40088
rect 15656 40008 15703 40072
rect 15767 40008 15783 40072
rect 15656 39992 15783 40008
rect 15656 39928 15703 39992
rect 15767 39928 15783 39992
rect 15656 39912 15783 39928
rect 15656 39848 15703 39912
rect 15767 39848 15783 39912
rect 15656 39832 15783 39848
rect 15656 39768 15703 39832
rect 15767 39768 15783 39832
rect 15656 39752 15783 39768
rect 15656 39688 15703 39752
rect 15767 39688 15783 39752
rect 15656 39672 15783 39688
rect 15656 39608 15703 39672
rect 15767 39608 15783 39672
rect 15656 39592 15783 39608
rect 15656 39528 15703 39592
rect 15767 39528 15783 39592
rect 15656 39512 15783 39528
rect 15656 39448 15703 39512
rect 15767 39448 15783 39512
rect 15656 39432 15783 39448
rect 15656 39368 15703 39432
rect 15767 39368 15783 39432
rect 15656 39352 15783 39368
rect 15656 39288 15703 39352
rect 15767 39288 15783 39352
rect 15656 39272 15783 39288
rect 15656 39208 15703 39272
rect 15767 39208 15783 39272
rect 15656 39192 15783 39208
rect 15656 39128 15703 39192
rect 15767 39128 15783 39192
rect 15656 39112 15783 39128
rect 15656 39048 15703 39112
rect 15767 39048 15783 39112
rect 15656 39032 15783 39048
rect 15656 38968 15703 39032
rect 15767 38968 15783 39032
rect 15656 38952 15783 38968
rect 15656 38888 15703 38952
rect 15767 38888 15783 38952
rect 15656 38872 15783 38888
rect 15656 38808 15703 38872
rect 15767 38808 15783 38872
rect 15656 38792 15783 38808
rect 15656 38728 15703 38792
rect 15767 38728 15783 38792
rect 15656 38712 15783 38728
rect 15656 38648 15703 38712
rect 15767 38648 15783 38712
rect 15656 38632 15783 38648
rect 15656 38568 15703 38632
rect 15767 38568 15783 38632
rect 15656 38552 15783 38568
rect 15656 38488 15703 38552
rect 15767 38488 15783 38552
rect 15656 38472 15783 38488
rect 15656 38408 15703 38472
rect 15767 38408 15783 38472
rect 15656 38392 15783 38408
rect 15656 38328 15703 38392
rect 15767 38328 15783 38392
rect 15656 38312 15783 38328
rect 15656 38248 15703 38312
rect 15767 38248 15783 38312
rect 15656 38232 15783 38248
rect 15656 38168 15703 38232
rect 15767 38168 15783 38232
rect 15656 38152 15783 38168
rect 15656 38088 15703 38152
rect 15767 38088 15783 38152
rect 15656 38072 15783 38088
rect 15656 38008 15703 38072
rect 15767 38008 15783 38072
rect 15656 37992 15783 38008
rect 15656 37928 15703 37992
rect 15767 37928 15783 37992
rect 15656 37912 15783 37928
rect 15656 37848 15703 37912
rect 15767 37848 15783 37912
rect 15656 37832 15783 37848
rect 15656 37768 15703 37832
rect 15767 37768 15783 37832
rect 15656 37752 15783 37768
rect 15656 37688 15703 37752
rect 15767 37688 15783 37752
rect 15656 37672 15783 37688
rect 15656 37608 15703 37672
rect 15767 37608 15783 37672
rect 15656 37592 15783 37608
rect 15656 37528 15703 37592
rect 15767 37528 15783 37592
rect 15656 37512 15783 37528
rect 15656 37448 15703 37512
rect 15767 37448 15783 37512
rect 15656 37432 15783 37448
rect 15656 37368 15703 37432
rect 15767 37368 15783 37432
rect 15656 37352 15783 37368
rect 15656 37288 15703 37352
rect 15767 37288 15783 37352
rect 15656 37272 15783 37288
rect 15656 37208 15703 37272
rect 15767 37208 15783 37272
rect 15656 37192 15783 37208
rect 15656 37128 15703 37192
rect 15767 37128 15783 37192
rect 15656 37112 15783 37128
rect 15656 37048 15703 37112
rect 15767 37048 15783 37112
rect 15656 37032 15783 37048
rect 15656 36968 15703 37032
rect 15767 36968 15783 37032
rect 15656 36952 15783 36968
rect 15656 36888 15703 36952
rect 15767 36888 15783 36952
rect 15656 36872 15783 36888
rect 15656 36808 15703 36872
rect 15767 36808 15783 36872
rect 15656 36792 15783 36808
rect 15656 36728 15703 36792
rect 15767 36728 15783 36792
rect 15656 36712 15783 36728
rect 15656 36648 15703 36712
rect 15767 36648 15783 36712
rect 15656 36632 15783 36648
rect 15656 36568 15703 36632
rect 15767 36568 15783 36632
rect 15656 36552 15783 36568
rect 15656 36488 15703 36552
rect 15767 36488 15783 36552
rect 15656 36472 15783 36488
rect 15656 36408 15703 36472
rect 15767 36408 15783 36472
rect 15656 36392 15783 36408
rect 15656 36328 15703 36392
rect 15767 36328 15783 36392
rect 15656 36312 15783 36328
rect 15656 36248 15703 36312
rect 15767 36248 15783 36312
rect 15656 36232 15783 36248
rect 15656 36168 15703 36232
rect 15767 36168 15783 36232
rect 15656 36152 15783 36168
rect 15656 36088 15703 36152
rect 15767 36088 15783 36152
rect 15656 36072 15783 36088
rect 15656 36008 15703 36072
rect 15767 36008 15783 36072
rect 15656 35992 15783 36008
rect 15656 35928 15703 35992
rect 15767 35928 15783 35992
rect 15656 35912 15783 35928
rect 15656 35848 15703 35912
rect 15767 35848 15783 35912
rect 15656 35832 15783 35848
rect 15656 35768 15703 35832
rect 15767 35768 15783 35832
rect 15656 35752 15783 35768
rect 15656 35688 15703 35752
rect 15767 35688 15783 35752
rect 15656 35672 15783 35688
rect 15656 35608 15703 35672
rect 15767 35608 15783 35672
rect 15656 35592 15783 35608
rect 15656 35528 15703 35592
rect 15767 35528 15783 35592
rect 15656 35512 15783 35528
rect 15656 35448 15703 35512
rect 15767 35448 15783 35512
rect 15656 35432 15783 35448
rect 15656 35368 15703 35432
rect 15767 35368 15783 35432
rect 15656 35352 15783 35368
rect 15656 35288 15703 35352
rect 15767 35288 15783 35352
rect 15656 35272 15783 35288
rect 15656 35208 15703 35272
rect 15767 35208 15783 35272
rect 15656 35192 15783 35208
rect 15656 35128 15703 35192
rect 15767 35128 15783 35192
rect 15656 35112 15783 35128
rect 15656 35048 15703 35112
rect 15767 35048 15783 35112
rect 15656 35032 15783 35048
rect 15656 34968 15703 35032
rect 15767 34968 15783 35032
rect 15656 34952 15783 34968
rect 15656 34888 15703 34952
rect 15767 34888 15783 34952
rect 15656 34872 15783 34888
rect 9337 34792 9464 34808
rect 9337 34728 9384 34792
rect 9448 34728 9464 34792
rect 9337 34712 9464 34728
rect 9337 34588 9441 34712
rect 9337 34572 9464 34588
rect 9337 34508 9384 34572
rect 9448 34508 9464 34572
rect 9337 34492 9464 34508
rect 3018 34412 3145 34428
rect 3018 34348 3065 34412
rect 3129 34348 3145 34412
rect 3018 34332 3145 34348
rect 3018 34268 3065 34332
rect 3129 34268 3145 34332
rect 3018 34252 3145 34268
rect 3018 34188 3065 34252
rect 3129 34188 3145 34252
rect 3018 34172 3145 34188
rect 3018 34108 3065 34172
rect 3129 34108 3145 34172
rect 3018 34092 3145 34108
rect 3018 34028 3065 34092
rect 3129 34028 3145 34092
rect 3018 34012 3145 34028
rect 3018 33948 3065 34012
rect 3129 33948 3145 34012
rect 3018 33932 3145 33948
rect 3018 33868 3065 33932
rect 3129 33868 3145 33932
rect 3018 33852 3145 33868
rect 3018 33788 3065 33852
rect 3129 33788 3145 33852
rect 3018 33772 3145 33788
rect 3018 33708 3065 33772
rect 3129 33708 3145 33772
rect 3018 33692 3145 33708
rect 3018 33628 3065 33692
rect 3129 33628 3145 33692
rect 3018 33612 3145 33628
rect 3018 33548 3065 33612
rect 3129 33548 3145 33612
rect 3018 33532 3145 33548
rect 3018 33468 3065 33532
rect 3129 33468 3145 33532
rect 3018 33452 3145 33468
rect 3018 33388 3065 33452
rect 3129 33388 3145 33452
rect 3018 33372 3145 33388
rect 3018 33308 3065 33372
rect 3129 33308 3145 33372
rect 3018 33292 3145 33308
rect 3018 33228 3065 33292
rect 3129 33228 3145 33292
rect 3018 33212 3145 33228
rect 3018 33148 3065 33212
rect 3129 33148 3145 33212
rect 3018 33132 3145 33148
rect 3018 33068 3065 33132
rect 3129 33068 3145 33132
rect 3018 33052 3145 33068
rect 3018 32988 3065 33052
rect 3129 32988 3145 33052
rect 3018 32972 3145 32988
rect 3018 32908 3065 32972
rect 3129 32908 3145 32972
rect 3018 32892 3145 32908
rect 3018 32828 3065 32892
rect 3129 32828 3145 32892
rect 3018 32812 3145 32828
rect 3018 32748 3065 32812
rect 3129 32748 3145 32812
rect 3018 32732 3145 32748
rect 3018 32668 3065 32732
rect 3129 32668 3145 32732
rect 3018 32652 3145 32668
rect 3018 32588 3065 32652
rect 3129 32588 3145 32652
rect 3018 32572 3145 32588
rect 3018 32508 3065 32572
rect 3129 32508 3145 32572
rect 3018 32492 3145 32508
rect 3018 32428 3065 32492
rect 3129 32428 3145 32492
rect 3018 32412 3145 32428
rect 3018 32348 3065 32412
rect 3129 32348 3145 32412
rect 3018 32332 3145 32348
rect 3018 32268 3065 32332
rect 3129 32268 3145 32332
rect 3018 32252 3145 32268
rect 3018 32188 3065 32252
rect 3129 32188 3145 32252
rect 3018 32172 3145 32188
rect 3018 32108 3065 32172
rect 3129 32108 3145 32172
rect 3018 32092 3145 32108
rect 3018 32028 3065 32092
rect 3129 32028 3145 32092
rect 3018 32012 3145 32028
rect 3018 31948 3065 32012
rect 3129 31948 3145 32012
rect 3018 31932 3145 31948
rect 3018 31868 3065 31932
rect 3129 31868 3145 31932
rect 3018 31852 3145 31868
rect 3018 31788 3065 31852
rect 3129 31788 3145 31852
rect 3018 31772 3145 31788
rect 3018 31708 3065 31772
rect 3129 31708 3145 31772
rect 3018 31692 3145 31708
rect 3018 31628 3065 31692
rect 3129 31628 3145 31692
rect 3018 31612 3145 31628
rect 3018 31548 3065 31612
rect 3129 31548 3145 31612
rect 3018 31532 3145 31548
rect 3018 31468 3065 31532
rect 3129 31468 3145 31532
rect 3018 31452 3145 31468
rect 3018 31388 3065 31452
rect 3129 31388 3145 31452
rect 3018 31372 3145 31388
rect 3018 31308 3065 31372
rect 3129 31308 3145 31372
rect 3018 31292 3145 31308
rect 3018 31228 3065 31292
rect 3129 31228 3145 31292
rect 3018 31212 3145 31228
rect 3018 31148 3065 31212
rect 3129 31148 3145 31212
rect 3018 31132 3145 31148
rect 3018 31068 3065 31132
rect 3129 31068 3145 31132
rect 3018 31052 3145 31068
rect 3018 30988 3065 31052
rect 3129 30988 3145 31052
rect 3018 30972 3145 30988
rect 3018 30908 3065 30972
rect 3129 30908 3145 30972
rect 3018 30892 3145 30908
rect 3018 30828 3065 30892
rect 3129 30828 3145 30892
rect 3018 30812 3145 30828
rect 3018 30748 3065 30812
rect 3129 30748 3145 30812
rect 3018 30732 3145 30748
rect 3018 30668 3065 30732
rect 3129 30668 3145 30732
rect 3018 30652 3145 30668
rect 3018 30588 3065 30652
rect 3129 30588 3145 30652
rect 3018 30572 3145 30588
rect 3018 30508 3065 30572
rect 3129 30508 3145 30572
rect 3018 30492 3145 30508
rect 3018 30428 3065 30492
rect 3129 30428 3145 30492
rect 3018 30412 3145 30428
rect 3018 30348 3065 30412
rect 3129 30348 3145 30412
rect 3018 30332 3145 30348
rect 3018 30268 3065 30332
rect 3129 30268 3145 30332
rect 3018 30252 3145 30268
rect 3018 30188 3065 30252
rect 3129 30188 3145 30252
rect 3018 30172 3145 30188
rect 3018 30108 3065 30172
rect 3129 30108 3145 30172
rect 3018 30092 3145 30108
rect 3018 30028 3065 30092
rect 3129 30028 3145 30092
rect 3018 30012 3145 30028
rect 3018 29948 3065 30012
rect 3129 29948 3145 30012
rect 3018 29932 3145 29948
rect 3018 29868 3065 29932
rect 3129 29868 3145 29932
rect 3018 29852 3145 29868
rect 3018 29788 3065 29852
rect 3129 29788 3145 29852
rect 3018 29772 3145 29788
rect 3018 29708 3065 29772
rect 3129 29708 3145 29772
rect 3018 29692 3145 29708
rect 3018 29628 3065 29692
rect 3129 29628 3145 29692
rect 3018 29612 3145 29628
rect 3018 29548 3065 29612
rect 3129 29548 3145 29612
rect 3018 29532 3145 29548
rect 3018 29468 3065 29532
rect 3129 29468 3145 29532
rect 3018 29452 3145 29468
rect 3018 29388 3065 29452
rect 3129 29388 3145 29452
rect 3018 29372 3145 29388
rect 3018 29308 3065 29372
rect 3129 29308 3145 29372
rect 3018 29292 3145 29308
rect 3018 29228 3065 29292
rect 3129 29228 3145 29292
rect 3018 29212 3145 29228
rect 3018 29148 3065 29212
rect 3129 29148 3145 29212
rect 3018 29132 3145 29148
rect 3018 29068 3065 29132
rect 3129 29068 3145 29132
rect 3018 29052 3145 29068
rect 3018 28988 3065 29052
rect 3129 28988 3145 29052
rect 3018 28972 3145 28988
rect 3018 28908 3065 28972
rect 3129 28908 3145 28972
rect 3018 28892 3145 28908
rect 3018 28828 3065 28892
rect 3129 28828 3145 28892
rect 3018 28812 3145 28828
rect 3018 28748 3065 28812
rect 3129 28748 3145 28812
rect 3018 28732 3145 28748
rect 3018 28668 3065 28732
rect 3129 28668 3145 28732
rect 3018 28652 3145 28668
rect 3018 28588 3065 28652
rect 3129 28588 3145 28652
rect 3018 28572 3145 28588
rect -3301 28492 -3174 28508
rect -3301 28428 -3254 28492
rect -3190 28428 -3174 28492
rect -3301 28412 -3174 28428
rect -3301 28288 -3197 28412
rect -3301 28272 -3174 28288
rect -3301 28208 -3254 28272
rect -3190 28208 -3174 28272
rect -3301 28192 -3174 28208
rect -9620 28112 -9493 28128
rect -9620 28048 -9573 28112
rect -9509 28048 -9493 28112
rect -9620 28032 -9493 28048
rect -9620 27968 -9573 28032
rect -9509 27968 -9493 28032
rect -9620 27952 -9493 27968
rect -9620 27888 -9573 27952
rect -9509 27888 -9493 27952
rect -9620 27872 -9493 27888
rect -9620 27808 -9573 27872
rect -9509 27808 -9493 27872
rect -9620 27792 -9493 27808
rect -9620 27728 -9573 27792
rect -9509 27728 -9493 27792
rect -9620 27712 -9493 27728
rect -9620 27648 -9573 27712
rect -9509 27648 -9493 27712
rect -9620 27632 -9493 27648
rect -9620 27568 -9573 27632
rect -9509 27568 -9493 27632
rect -9620 27552 -9493 27568
rect -9620 27488 -9573 27552
rect -9509 27488 -9493 27552
rect -9620 27472 -9493 27488
rect -9620 27408 -9573 27472
rect -9509 27408 -9493 27472
rect -9620 27392 -9493 27408
rect -9620 27328 -9573 27392
rect -9509 27328 -9493 27392
rect -9620 27312 -9493 27328
rect -9620 27248 -9573 27312
rect -9509 27248 -9493 27312
rect -9620 27232 -9493 27248
rect -9620 27168 -9573 27232
rect -9509 27168 -9493 27232
rect -9620 27152 -9493 27168
rect -9620 27088 -9573 27152
rect -9509 27088 -9493 27152
rect -9620 27072 -9493 27088
rect -9620 27008 -9573 27072
rect -9509 27008 -9493 27072
rect -9620 26992 -9493 27008
rect -9620 26928 -9573 26992
rect -9509 26928 -9493 26992
rect -9620 26912 -9493 26928
rect -9620 26848 -9573 26912
rect -9509 26848 -9493 26912
rect -9620 26832 -9493 26848
rect -9620 26768 -9573 26832
rect -9509 26768 -9493 26832
rect -9620 26752 -9493 26768
rect -9620 26688 -9573 26752
rect -9509 26688 -9493 26752
rect -9620 26672 -9493 26688
rect -9620 26608 -9573 26672
rect -9509 26608 -9493 26672
rect -9620 26592 -9493 26608
rect -9620 26528 -9573 26592
rect -9509 26528 -9493 26592
rect -9620 26512 -9493 26528
rect -9620 26448 -9573 26512
rect -9509 26448 -9493 26512
rect -9620 26432 -9493 26448
rect -9620 26368 -9573 26432
rect -9509 26368 -9493 26432
rect -9620 26352 -9493 26368
rect -9620 26288 -9573 26352
rect -9509 26288 -9493 26352
rect -9620 26272 -9493 26288
rect -9620 26208 -9573 26272
rect -9509 26208 -9493 26272
rect -9620 26192 -9493 26208
rect -9620 26128 -9573 26192
rect -9509 26128 -9493 26192
rect -9620 26112 -9493 26128
rect -9620 26048 -9573 26112
rect -9509 26048 -9493 26112
rect -9620 26032 -9493 26048
rect -9620 25968 -9573 26032
rect -9509 25968 -9493 26032
rect -9620 25952 -9493 25968
rect -9620 25888 -9573 25952
rect -9509 25888 -9493 25952
rect -9620 25872 -9493 25888
rect -9620 25808 -9573 25872
rect -9509 25808 -9493 25872
rect -9620 25792 -9493 25808
rect -9620 25728 -9573 25792
rect -9509 25728 -9493 25792
rect -9620 25712 -9493 25728
rect -9620 25648 -9573 25712
rect -9509 25648 -9493 25712
rect -9620 25632 -9493 25648
rect -9620 25568 -9573 25632
rect -9509 25568 -9493 25632
rect -9620 25552 -9493 25568
rect -9620 25488 -9573 25552
rect -9509 25488 -9493 25552
rect -9620 25472 -9493 25488
rect -9620 25408 -9573 25472
rect -9509 25408 -9493 25472
rect -9620 25392 -9493 25408
rect -9620 25328 -9573 25392
rect -9509 25328 -9493 25392
rect -9620 25312 -9493 25328
rect -9620 25248 -9573 25312
rect -9509 25248 -9493 25312
rect -9620 25232 -9493 25248
rect -9620 25168 -9573 25232
rect -9509 25168 -9493 25232
rect -9620 25152 -9493 25168
rect -9620 25088 -9573 25152
rect -9509 25088 -9493 25152
rect -9620 25072 -9493 25088
rect -9620 25008 -9573 25072
rect -9509 25008 -9493 25072
rect -9620 24992 -9493 25008
rect -9620 24928 -9573 24992
rect -9509 24928 -9493 24992
rect -9620 24912 -9493 24928
rect -9620 24848 -9573 24912
rect -9509 24848 -9493 24912
rect -9620 24832 -9493 24848
rect -9620 24768 -9573 24832
rect -9509 24768 -9493 24832
rect -9620 24752 -9493 24768
rect -9620 24688 -9573 24752
rect -9509 24688 -9493 24752
rect -9620 24672 -9493 24688
rect -9620 24608 -9573 24672
rect -9509 24608 -9493 24672
rect -9620 24592 -9493 24608
rect -9620 24528 -9573 24592
rect -9509 24528 -9493 24592
rect -9620 24512 -9493 24528
rect -9620 24448 -9573 24512
rect -9509 24448 -9493 24512
rect -9620 24432 -9493 24448
rect -9620 24368 -9573 24432
rect -9509 24368 -9493 24432
rect -9620 24352 -9493 24368
rect -9620 24288 -9573 24352
rect -9509 24288 -9493 24352
rect -9620 24272 -9493 24288
rect -9620 24208 -9573 24272
rect -9509 24208 -9493 24272
rect -9620 24192 -9493 24208
rect -9620 24128 -9573 24192
rect -9509 24128 -9493 24192
rect -9620 24112 -9493 24128
rect -9620 24048 -9573 24112
rect -9509 24048 -9493 24112
rect -9620 24032 -9493 24048
rect -9620 23968 -9573 24032
rect -9509 23968 -9493 24032
rect -9620 23952 -9493 23968
rect -9620 23888 -9573 23952
rect -9509 23888 -9493 23952
rect -9620 23872 -9493 23888
rect -9620 23808 -9573 23872
rect -9509 23808 -9493 23872
rect -9620 23792 -9493 23808
rect -9620 23728 -9573 23792
rect -9509 23728 -9493 23792
rect -9620 23712 -9493 23728
rect -9620 23648 -9573 23712
rect -9509 23648 -9493 23712
rect -9620 23632 -9493 23648
rect -9620 23568 -9573 23632
rect -9509 23568 -9493 23632
rect -9620 23552 -9493 23568
rect -9620 23488 -9573 23552
rect -9509 23488 -9493 23552
rect -9620 23472 -9493 23488
rect -9620 23408 -9573 23472
rect -9509 23408 -9493 23472
rect -9620 23392 -9493 23408
rect -9620 23328 -9573 23392
rect -9509 23328 -9493 23392
rect -9620 23312 -9493 23328
rect -9620 23248 -9573 23312
rect -9509 23248 -9493 23312
rect -9620 23232 -9493 23248
rect -9620 23168 -9573 23232
rect -9509 23168 -9493 23232
rect -9620 23152 -9493 23168
rect -9620 23088 -9573 23152
rect -9509 23088 -9493 23152
rect -9620 23072 -9493 23088
rect -9620 23008 -9573 23072
rect -9509 23008 -9493 23072
rect -9620 22992 -9493 23008
rect -9620 22928 -9573 22992
rect -9509 22928 -9493 22992
rect -9620 22912 -9493 22928
rect -9620 22848 -9573 22912
rect -9509 22848 -9493 22912
rect -9620 22832 -9493 22848
rect -9620 22768 -9573 22832
rect -9509 22768 -9493 22832
rect -9620 22752 -9493 22768
rect -9620 22688 -9573 22752
rect -9509 22688 -9493 22752
rect -9620 22672 -9493 22688
rect -9620 22608 -9573 22672
rect -9509 22608 -9493 22672
rect -9620 22592 -9493 22608
rect -9620 22528 -9573 22592
rect -9509 22528 -9493 22592
rect -9620 22512 -9493 22528
rect -9620 22448 -9573 22512
rect -9509 22448 -9493 22512
rect -9620 22432 -9493 22448
rect -9620 22368 -9573 22432
rect -9509 22368 -9493 22432
rect -9620 22352 -9493 22368
rect -9620 22288 -9573 22352
rect -9509 22288 -9493 22352
rect -9620 22272 -9493 22288
rect -15939 22192 -15812 22208
rect -15939 22128 -15892 22192
rect -15828 22128 -15812 22192
rect -15939 22112 -15812 22128
rect -15939 21988 -15835 22112
rect -15939 21972 -15812 21988
rect -15939 21908 -15892 21972
rect -15828 21908 -15812 21972
rect -15939 21892 -15812 21908
rect -22258 21812 -22131 21828
rect -22258 21748 -22211 21812
rect -22147 21748 -22131 21812
rect -22258 21732 -22131 21748
rect -22258 21668 -22211 21732
rect -22147 21668 -22131 21732
rect -22258 21652 -22131 21668
rect -22258 21588 -22211 21652
rect -22147 21588 -22131 21652
rect -22258 21572 -22131 21588
rect -22258 21508 -22211 21572
rect -22147 21508 -22131 21572
rect -22258 21492 -22131 21508
rect -22258 21428 -22211 21492
rect -22147 21428 -22131 21492
rect -22258 21412 -22131 21428
rect -22258 21348 -22211 21412
rect -22147 21348 -22131 21412
rect -22258 21332 -22131 21348
rect -22258 21268 -22211 21332
rect -22147 21268 -22131 21332
rect -22258 21252 -22131 21268
rect -22258 21188 -22211 21252
rect -22147 21188 -22131 21252
rect -22258 21172 -22131 21188
rect -22258 21108 -22211 21172
rect -22147 21108 -22131 21172
rect -22258 21092 -22131 21108
rect -22258 21028 -22211 21092
rect -22147 21028 -22131 21092
rect -22258 21012 -22131 21028
rect -22258 20948 -22211 21012
rect -22147 20948 -22131 21012
rect -22258 20932 -22131 20948
rect -22258 20868 -22211 20932
rect -22147 20868 -22131 20932
rect -22258 20852 -22131 20868
rect -22258 20788 -22211 20852
rect -22147 20788 -22131 20852
rect -22258 20772 -22131 20788
rect -22258 20708 -22211 20772
rect -22147 20708 -22131 20772
rect -22258 20692 -22131 20708
rect -22258 20628 -22211 20692
rect -22147 20628 -22131 20692
rect -22258 20612 -22131 20628
rect -22258 20548 -22211 20612
rect -22147 20548 -22131 20612
rect -22258 20532 -22131 20548
rect -22258 20468 -22211 20532
rect -22147 20468 -22131 20532
rect -22258 20452 -22131 20468
rect -22258 20388 -22211 20452
rect -22147 20388 -22131 20452
rect -22258 20372 -22131 20388
rect -22258 20308 -22211 20372
rect -22147 20308 -22131 20372
rect -22258 20292 -22131 20308
rect -22258 20228 -22211 20292
rect -22147 20228 -22131 20292
rect -22258 20212 -22131 20228
rect -22258 20148 -22211 20212
rect -22147 20148 -22131 20212
rect -22258 20132 -22131 20148
rect -22258 20068 -22211 20132
rect -22147 20068 -22131 20132
rect -22258 20052 -22131 20068
rect -22258 19988 -22211 20052
rect -22147 19988 -22131 20052
rect -22258 19972 -22131 19988
rect -22258 19908 -22211 19972
rect -22147 19908 -22131 19972
rect -22258 19892 -22131 19908
rect -22258 19828 -22211 19892
rect -22147 19828 -22131 19892
rect -22258 19812 -22131 19828
rect -22258 19748 -22211 19812
rect -22147 19748 -22131 19812
rect -22258 19732 -22131 19748
rect -22258 19668 -22211 19732
rect -22147 19668 -22131 19732
rect -22258 19652 -22131 19668
rect -22258 19588 -22211 19652
rect -22147 19588 -22131 19652
rect -22258 19572 -22131 19588
rect -22258 19508 -22211 19572
rect -22147 19508 -22131 19572
rect -22258 19492 -22131 19508
rect -22258 19428 -22211 19492
rect -22147 19428 -22131 19492
rect -22258 19412 -22131 19428
rect -22258 19348 -22211 19412
rect -22147 19348 -22131 19412
rect -22258 19332 -22131 19348
rect -22258 19268 -22211 19332
rect -22147 19268 -22131 19332
rect -22258 19252 -22131 19268
rect -22258 19188 -22211 19252
rect -22147 19188 -22131 19252
rect -22258 19172 -22131 19188
rect -22258 19108 -22211 19172
rect -22147 19108 -22131 19172
rect -22258 19092 -22131 19108
rect -22258 19028 -22211 19092
rect -22147 19028 -22131 19092
rect -22258 19012 -22131 19028
rect -22258 18948 -22211 19012
rect -22147 18948 -22131 19012
rect -22258 18932 -22131 18948
rect -22258 18868 -22211 18932
rect -22147 18868 -22131 18932
rect -22258 18852 -22131 18868
rect -22258 18788 -22211 18852
rect -22147 18788 -22131 18852
rect -22258 18772 -22131 18788
rect -22258 18708 -22211 18772
rect -22147 18708 -22131 18772
rect -22258 18692 -22131 18708
rect -22258 18628 -22211 18692
rect -22147 18628 -22131 18692
rect -22258 18612 -22131 18628
rect -22258 18548 -22211 18612
rect -22147 18548 -22131 18612
rect -22258 18532 -22131 18548
rect -22258 18468 -22211 18532
rect -22147 18468 -22131 18532
rect -22258 18452 -22131 18468
rect -22258 18388 -22211 18452
rect -22147 18388 -22131 18452
rect -22258 18372 -22131 18388
rect -22258 18308 -22211 18372
rect -22147 18308 -22131 18372
rect -22258 18292 -22131 18308
rect -22258 18228 -22211 18292
rect -22147 18228 -22131 18292
rect -22258 18212 -22131 18228
rect -22258 18148 -22211 18212
rect -22147 18148 -22131 18212
rect -22258 18132 -22131 18148
rect -22258 18068 -22211 18132
rect -22147 18068 -22131 18132
rect -22258 18052 -22131 18068
rect -22258 17988 -22211 18052
rect -22147 17988 -22131 18052
rect -22258 17972 -22131 17988
rect -22258 17908 -22211 17972
rect -22147 17908 -22131 17972
rect -22258 17892 -22131 17908
rect -22258 17828 -22211 17892
rect -22147 17828 -22131 17892
rect -22258 17812 -22131 17828
rect -22258 17748 -22211 17812
rect -22147 17748 -22131 17812
rect -22258 17732 -22131 17748
rect -22258 17668 -22211 17732
rect -22147 17668 -22131 17732
rect -22258 17652 -22131 17668
rect -22258 17588 -22211 17652
rect -22147 17588 -22131 17652
rect -22258 17572 -22131 17588
rect -22258 17508 -22211 17572
rect -22147 17508 -22131 17572
rect -22258 17492 -22131 17508
rect -22258 17428 -22211 17492
rect -22147 17428 -22131 17492
rect -22258 17412 -22131 17428
rect -22258 17348 -22211 17412
rect -22147 17348 -22131 17412
rect -22258 17332 -22131 17348
rect -22258 17268 -22211 17332
rect -22147 17268 -22131 17332
rect -22258 17252 -22131 17268
rect -22258 17188 -22211 17252
rect -22147 17188 -22131 17252
rect -22258 17172 -22131 17188
rect -22258 17108 -22211 17172
rect -22147 17108 -22131 17172
rect -22258 17092 -22131 17108
rect -22258 17028 -22211 17092
rect -22147 17028 -22131 17092
rect -22258 17012 -22131 17028
rect -22258 16948 -22211 17012
rect -22147 16948 -22131 17012
rect -22258 16932 -22131 16948
rect -22258 16868 -22211 16932
rect -22147 16868 -22131 16932
rect -22258 16852 -22131 16868
rect -22258 16788 -22211 16852
rect -22147 16788 -22131 16852
rect -22258 16772 -22131 16788
rect -22258 16708 -22211 16772
rect -22147 16708 -22131 16772
rect -22258 16692 -22131 16708
rect -22258 16628 -22211 16692
rect -22147 16628 -22131 16692
rect -22258 16612 -22131 16628
rect -22258 16548 -22211 16612
rect -22147 16548 -22131 16612
rect -22258 16532 -22131 16548
rect -22258 16468 -22211 16532
rect -22147 16468 -22131 16532
rect -22258 16452 -22131 16468
rect -22258 16388 -22211 16452
rect -22147 16388 -22131 16452
rect -22258 16372 -22131 16388
rect -22258 16308 -22211 16372
rect -22147 16308 -22131 16372
rect -22258 16292 -22131 16308
rect -22258 16228 -22211 16292
rect -22147 16228 -22131 16292
rect -22258 16212 -22131 16228
rect -22258 16148 -22211 16212
rect -22147 16148 -22131 16212
rect -22258 16132 -22131 16148
rect -22258 16068 -22211 16132
rect -22147 16068 -22131 16132
rect -22258 16052 -22131 16068
rect -22258 15988 -22211 16052
rect -22147 15988 -22131 16052
rect -22258 15972 -22131 15988
rect -28577 15892 -28450 15908
rect -28577 15828 -28530 15892
rect -28466 15828 -28450 15892
rect -28577 15812 -28450 15828
rect -28577 15688 -28473 15812
rect -28577 15672 -28450 15688
rect -28577 15608 -28530 15672
rect -28466 15608 -28450 15672
rect -28577 15592 -28450 15608
rect -34896 15512 -34769 15528
rect -34896 15448 -34849 15512
rect -34785 15448 -34769 15512
rect -34896 15432 -34769 15448
rect -34896 15368 -34849 15432
rect -34785 15368 -34769 15432
rect -34896 15352 -34769 15368
rect -34896 15288 -34849 15352
rect -34785 15288 -34769 15352
rect -34896 15272 -34769 15288
rect -34896 15208 -34849 15272
rect -34785 15208 -34769 15272
rect -34896 15192 -34769 15208
rect -34896 15128 -34849 15192
rect -34785 15128 -34769 15192
rect -34896 15112 -34769 15128
rect -34896 15048 -34849 15112
rect -34785 15048 -34769 15112
rect -34896 15032 -34769 15048
rect -34896 14968 -34849 15032
rect -34785 14968 -34769 15032
rect -34896 14952 -34769 14968
rect -34896 14888 -34849 14952
rect -34785 14888 -34769 14952
rect -34896 14872 -34769 14888
rect -34896 14808 -34849 14872
rect -34785 14808 -34769 14872
rect -34896 14792 -34769 14808
rect -34896 14728 -34849 14792
rect -34785 14728 -34769 14792
rect -34896 14712 -34769 14728
rect -34896 14648 -34849 14712
rect -34785 14648 -34769 14712
rect -34896 14632 -34769 14648
rect -34896 14568 -34849 14632
rect -34785 14568 -34769 14632
rect -34896 14552 -34769 14568
rect -34896 14488 -34849 14552
rect -34785 14488 -34769 14552
rect -34896 14472 -34769 14488
rect -34896 14408 -34849 14472
rect -34785 14408 -34769 14472
rect -34896 14392 -34769 14408
rect -34896 14328 -34849 14392
rect -34785 14328 -34769 14392
rect -34896 14312 -34769 14328
rect -34896 14248 -34849 14312
rect -34785 14248 -34769 14312
rect -34896 14232 -34769 14248
rect -34896 14168 -34849 14232
rect -34785 14168 -34769 14232
rect -34896 14152 -34769 14168
rect -34896 14088 -34849 14152
rect -34785 14088 -34769 14152
rect -34896 14072 -34769 14088
rect -34896 14008 -34849 14072
rect -34785 14008 -34769 14072
rect -34896 13992 -34769 14008
rect -34896 13928 -34849 13992
rect -34785 13928 -34769 13992
rect -34896 13912 -34769 13928
rect -34896 13848 -34849 13912
rect -34785 13848 -34769 13912
rect -34896 13832 -34769 13848
rect -34896 13768 -34849 13832
rect -34785 13768 -34769 13832
rect -34896 13752 -34769 13768
rect -34896 13688 -34849 13752
rect -34785 13688 -34769 13752
rect -34896 13672 -34769 13688
rect -34896 13608 -34849 13672
rect -34785 13608 -34769 13672
rect -34896 13592 -34769 13608
rect -34896 13528 -34849 13592
rect -34785 13528 -34769 13592
rect -34896 13512 -34769 13528
rect -34896 13448 -34849 13512
rect -34785 13448 -34769 13512
rect -34896 13432 -34769 13448
rect -34896 13368 -34849 13432
rect -34785 13368 -34769 13432
rect -34896 13352 -34769 13368
rect -34896 13288 -34849 13352
rect -34785 13288 -34769 13352
rect -34896 13272 -34769 13288
rect -34896 13208 -34849 13272
rect -34785 13208 -34769 13272
rect -34896 13192 -34769 13208
rect -34896 13128 -34849 13192
rect -34785 13128 -34769 13192
rect -34896 13112 -34769 13128
rect -34896 13048 -34849 13112
rect -34785 13048 -34769 13112
rect -34896 13032 -34769 13048
rect -34896 12968 -34849 13032
rect -34785 12968 -34769 13032
rect -34896 12952 -34769 12968
rect -34896 12888 -34849 12952
rect -34785 12888 -34769 12952
rect -34896 12872 -34769 12888
rect -34896 12808 -34849 12872
rect -34785 12808 -34769 12872
rect -34896 12792 -34769 12808
rect -34896 12728 -34849 12792
rect -34785 12728 -34769 12792
rect -34896 12712 -34769 12728
rect -34896 12648 -34849 12712
rect -34785 12648 -34769 12712
rect -34896 12632 -34769 12648
rect -34896 12568 -34849 12632
rect -34785 12568 -34769 12632
rect -34896 12552 -34769 12568
rect -34896 12488 -34849 12552
rect -34785 12488 -34769 12552
rect -34896 12472 -34769 12488
rect -34896 12408 -34849 12472
rect -34785 12408 -34769 12472
rect -34896 12392 -34769 12408
rect -34896 12328 -34849 12392
rect -34785 12328 -34769 12392
rect -34896 12312 -34769 12328
rect -34896 12248 -34849 12312
rect -34785 12248 -34769 12312
rect -34896 12232 -34769 12248
rect -34896 12168 -34849 12232
rect -34785 12168 -34769 12232
rect -34896 12152 -34769 12168
rect -34896 12088 -34849 12152
rect -34785 12088 -34769 12152
rect -34896 12072 -34769 12088
rect -34896 12008 -34849 12072
rect -34785 12008 -34769 12072
rect -34896 11992 -34769 12008
rect -34896 11928 -34849 11992
rect -34785 11928 -34769 11992
rect -34896 11912 -34769 11928
rect -34896 11848 -34849 11912
rect -34785 11848 -34769 11912
rect -34896 11832 -34769 11848
rect -34896 11768 -34849 11832
rect -34785 11768 -34769 11832
rect -34896 11752 -34769 11768
rect -34896 11688 -34849 11752
rect -34785 11688 -34769 11752
rect -34896 11672 -34769 11688
rect -34896 11608 -34849 11672
rect -34785 11608 -34769 11672
rect -34896 11592 -34769 11608
rect -34896 11528 -34849 11592
rect -34785 11528 -34769 11592
rect -34896 11512 -34769 11528
rect -34896 11448 -34849 11512
rect -34785 11448 -34769 11512
rect -34896 11432 -34769 11448
rect -34896 11368 -34849 11432
rect -34785 11368 -34769 11432
rect -34896 11352 -34769 11368
rect -34896 11288 -34849 11352
rect -34785 11288 -34769 11352
rect -34896 11272 -34769 11288
rect -34896 11208 -34849 11272
rect -34785 11208 -34769 11272
rect -34896 11192 -34769 11208
rect -34896 11128 -34849 11192
rect -34785 11128 -34769 11192
rect -34896 11112 -34769 11128
rect -34896 11048 -34849 11112
rect -34785 11048 -34769 11112
rect -34896 11032 -34769 11048
rect -34896 10968 -34849 11032
rect -34785 10968 -34769 11032
rect -34896 10952 -34769 10968
rect -34896 10888 -34849 10952
rect -34785 10888 -34769 10952
rect -34896 10872 -34769 10888
rect -34896 10808 -34849 10872
rect -34785 10808 -34769 10872
rect -34896 10792 -34769 10808
rect -34896 10728 -34849 10792
rect -34785 10728 -34769 10792
rect -34896 10712 -34769 10728
rect -34896 10648 -34849 10712
rect -34785 10648 -34769 10712
rect -34896 10632 -34769 10648
rect -34896 10568 -34849 10632
rect -34785 10568 -34769 10632
rect -34896 10552 -34769 10568
rect -34896 10488 -34849 10552
rect -34785 10488 -34769 10552
rect -34896 10472 -34769 10488
rect -34896 10408 -34849 10472
rect -34785 10408 -34769 10472
rect -34896 10392 -34769 10408
rect -34896 10328 -34849 10392
rect -34785 10328 -34769 10392
rect -34896 10312 -34769 10328
rect -34896 10248 -34849 10312
rect -34785 10248 -34769 10312
rect -34896 10232 -34769 10248
rect -34896 10168 -34849 10232
rect -34785 10168 -34769 10232
rect -34896 10152 -34769 10168
rect -34896 10088 -34849 10152
rect -34785 10088 -34769 10152
rect -34896 10072 -34769 10088
rect -34896 10008 -34849 10072
rect -34785 10008 -34769 10072
rect -34896 9992 -34769 10008
rect -34896 9928 -34849 9992
rect -34785 9928 -34769 9992
rect -34896 9912 -34769 9928
rect -34896 9848 -34849 9912
rect -34785 9848 -34769 9912
rect -34896 9832 -34769 9848
rect -34896 9768 -34849 9832
rect -34785 9768 -34769 9832
rect -34896 9752 -34769 9768
rect -34896 9688 -34849 9752
rect -34785 9688 -34769 9752
rect -34896 9672 -34769 9688
rect -41215 9592 -41088 9608
rect -41215 9528 -41168 9592
rect -41104 9528 -41088 9592
rect -41215 9512 -41088 9528
rect -41215 9388 -41111 9512
rect -41215 9372 -41088 9388
rect -41215 9308 -41168 9372
rect -41104 9308 -41088 9372
rect -41215 9292 -41088 9308
rect -47244 9252 -41322 9261
rect -47244 3348 -47235 9252
rect -41331 3348 -41322 9252
rect -47244 3339 -41322 3348
rect -41215 9228 -41168 9292
rect -41104 9228 -41088 9292
rect -38016 9261 -37912 9639
rect -34896 9608 -34849 9672
rect -34785 9608 -34769 9672
rect -34606 15552 -28684 15561
rect -34606 9648 -34597 15552
rect -28693 9648 -28684 15552
rect -34606 9639 -28684 9648
rect -28577 15528 -28530 15592
rect -28466 15528 -28450 15592
rect -25378 15561 -25274 15939
rect -22258 15908 -22211 15972
rect -22147 15908 -22131 15972
rect -21968 21852 -16046 21861
rect -21968 15948 -21959 21852
rect -16055 15948 -16046 21852
rect -21968 15939 -16046 15948
rect -15939 21828 -15892 21892
rect -15828 21828 -15812 21892
rect -12740 21861 -12636 22239
rect -9620 22208 -9573 22272
rect -9509 22208 -9493 22272
rect -9330 28152 -3408 28161
rect -9330 22248 -9321 28152
rect -3417 22248 -3408 28152
rect -9330 22239 -3408 22248
rect -3301 28128 -3254 28192
rect -3190 28128 -3174 28192
rect -102 28161 2 28539
rect 3018 28508 3065 28572
rect 3129 28508 3145 28572
rect 3308 34452 9230 34461
rect 3308 28548 3317 34452
rect 9221 28548 9230 34452
rect 3308 28539 9230 28548
rect 9337 34428 9384 34492
rect 9448 34428 9464 34492
rect 12536 34461 12640 34839
rect 15656 34808 15703 34872
rect 15767 34808 15783 34872
rect 15946 40752 21868 40761
rect 15946 34848 15955 40752
rect 21859 34848 21868 40752
rect 15946 34839 21868 34848
rect 21975 40728 22022 40792
rect 22086 40728 22102 40792
rect 25174 40761 25278 41139
rect 28294 41108 28341 41172
rect 28405 41108 28421 41172
rect 28584 47052 34506 47061
rect 28584 41148 28593 47052
rect 34497 41148 34506 47052
rect 28584 41139 34506 41148
rect 34613 47028 34660 47092
rect 34724 47028 34740 47092
rect 37812 47061 37916 47250
rect 40932 47188 41036 47250
rect 40932 47172 41059 47188
rect 40932 47108 40979 47172
rect 41043 47108 41059 47172
rect 40932 47092 41059 47108
rect 34613 47012 34740 47028
rect 34613 46948 34660 47012
rect 34724 46948 34740 47012
rect 34613 46932 34740 46948
rect 34613 46868 34660 46932
rect 34724 46868 34740 46932
rect 34613 46852 34740 46868
rect 34613 46788 34660 46852
rect 34724 46788 34740 46852
rect 34613 46772 34740 46788
rect 34613 46708 34660 46772
rect 34724 46708 34740 46772
rect 34613 46692 34740 46708
rect 34613 46628 34660 46692
rect 34724 46628 34740 46692
rect 34613 46612 34740 46628
rect 34613 46548 34660 46612
rect 34724 46548 34740 46612
rect 34613 46532 34740 46548
rect 34613 46468 34660 46532
rect 34724 46468 34740 46532
rect 34613 46452 34740 46468
rect 34613 46388 34660 46452
rect 34724 46388 34740 46452
rect 34613 46372 34740 46388
rect 34613 46308 34660 46372
rect 34724 46308 34740 46372
rect 34613 46292 34740 46308
rect 34613 46228 34660 46292
rect 34724 46228 34740 46292
rect 34613 46212 34740 46228
rect 34613 46148 34660 46212
rect 34724 46148 34740 46212
rect 34613 46132 34740 46148
rect 34613 46068 34660 46132
rect 34724 46068 34740 46132
rect 34613 46052 34740 46068
rect 34613 45988 34660 46052
rect 34724 45988 34740 46052
rect 34613 45972 34740 45988
rect 34613 45908 34660 45972
rect 34724 45908 34740 45972
rect 34613 45892 34740 45908
rect 34613 45828 34660 45892
rect 34724 45828 34740 45892
rect 34613 45812 34740 45828
rect 34613 45748 34660 45812
rect 34724 45748 34740 45812
rect 34613 45732 34740 45748
rect 34613 45668 34660 45732
rect 34724 45668 34740 45732
rect 34613 45652 34740 45668
rect 34613 45588 34660 45652
rect 34724 45588 34740 45652
rect 34613 45572 34740 45588
rect 34613 45508 34660 45572
rect 34724 45508 34740 45572
rect 34613 45492 34740 45508
rect 34613 45428 34660 45492
rect 34724 45428 34740 45492
rect 34613 45412 34740 45428
rect 34613 45348 34660 45412
rect 34724 45348 34740 45412
rect 34613 45332 34740 45348
rect 34613 45268 34660 45332
rect 34724 45268 34740 45332
rect 34613 45252 34740 45268
rect 34613 45188 34660 45252
rect 34724 45188 34740 45252
rect 34613 45172 34740 45188
rect 34613 45108 34660 45172
rect 34724 45108 34740 45172
rect 34613 45092 34740 45108
rect 34613 45028 34660 45092
rect 34724 45028 34740 45092
rect 34613 45012 34740 45028
rect 34613 44948 34660 45012
rect 34724 44948 34740 45012
rect 34613 44932 34740 44948
rect 34613 44868 34660 44932
rect 34724 44868 34740 44932
rect 34613 44852 34740 44868
rect 34613 44788 34660 44852
rect 34724 44788 34740 44852
rect 34613 44772 34740 44788
rect 34613 44708 34660 44772
rect 34724 44708 34740 44772
rect 34613 44692 34740 44708
rect 34613 44628 34660 44692
rect 34724 44628 34740 44692
rect 34613 44612 34740 44628
rect 34613 44548 34660 44612
rect 34724 44548 34740 44612
rect 34613 44532 34740 44548
rect 34613 44468 34660 44532
rect 34724 44468 34740 44532
rect 34613 44452 34740 44468
rect 34613 44388 34660 44452
rect 34724 44388 34740 44452
rect 34613 44372 34740 44388
rect 34613 44308 34660 44372
rect 34724 44308 34740 44372
rect 34613 44292 34740 44308
rect 34613 44228 34660 44292
rect 34724 44228 34740 44292
rect 34613 44212 34740 44228
rect 34613 44148 34660 44212
rect 34724 44148 34740 44212
rect 34613 44132 34740 44148
rect 34613 44068 34660 44132
rect 34724 44068 34740 44132
rect 34613 44052 34740 44068
rect 34613 43988 34660 44052
rect 34724 43988 34740 44052
rect 34613 43972 34740 43988
rect 34613 43908 34660 43972
rect 34724 43908 34740 43972
rect 34613 43892 34740 43908
rect 34613 43828 34660 43892
rect 34724 43828 34740 43892
rect 34613 43812 34740 43828
rect 34613 43748 34660 43812
rect 34724 43748 34740 43812
rect 34613 43732 34740 43748
rect 34613 43668 34660 43732
rect 34724 43668 34740 43732
rect 34613 43652 34740 43668
rect 34613 43588 34660 43652
rect 34724 43588 34740 43652
rect 34613 43572 34740 43588
rect 34613 43508 34660 43572
rect 34724 43508 34740 43572
rect 34613 43492 34740 43508
rect 34613 43428 34660 43492
rect 34724 43428 34740 43492
rect 34613 43412 34740 43428
rect 34613 43348 34660 43412
rect 34724 43348 34740 43412
rect 34613 43332 34740 43348
rect 34613 43268 34660 43332
rect 34724 43268 34740 43332
rect 34613 43252 34740 43268
rect 34613 43188 34660 43252
rect 34724 43188 34740 43252
rect 34613 43172 34740 43188
rect 34613 43108 34660 43172
rect 34724 43108 34740 43172
rect 34613 43092 34740 43108
rect 34613 43028 34660 43092
rect 34724 43028 34740 43092
rect 34613 43012 34740 43028
rect 34613 42948 34660 43012
rect 34724 42948 34740 43012
rect 34613 42932 34740 42948
rect 34613 42868 34660 42932
rect 34724 42868 34740 42932
rect 34613 42852 34740 42868
rect 34613 42788 34660 42852
rect 34724 42788 34740 42852
rect 34613 42772 34740 42788
rect 34613 42708 34660 42772
rect 34724 42708 34740 42772
rect 34613 42692 34740 42708
rect 34613 42628 34660 42692
rect 34724 42628 34740 42692
rect 34613 42612 34740 42628
rect 34613 42548 34660 42612
rect 34724 42548 34740 42612
rect 34613 42532 34740 42548
rect 34613 42468 34660 42532
rect 34724 42468 34740 42532
rect 34613 42452 34740 42468
rect 34613 42388 34660 42452
rect 34724 42388 34740 42452
rect 34613 42372 34740 42388
rect 34613 42308 34660 42372
rect 34724 42308 34740 42372
rect 34613 42292 34740 42308
rect 34613 42228 34660 42292
rect 34724 42228 34740 42292
rect 34613 42212 34740 42228
rect 34613 42148 34660 42212
rect 34724 42148 34740 42212
rect 34613 42132 34740 42148
rect 34613 42068 34660 42132
rect 34724 42068 34740 42132
rect 34613 42052 34740 42068
rect 34613 41988 34660 42052
rect 34724 41988 34740 42052
rect 34613 41972 34740 41988
rect 34613 41908 34660 41972
rect 34724 41908 34740 41972
rect 34613 41892 34740 41908
rect 34613 41828 34660 41892
rect 34724 41828 34740 41892
rect 34613 41812 34740 41828
rect 34613 41748 34660 41812
rect 34724 41748 34740 41812
rect 34613 41732 34740 41748
rect 34613 41668 34660 41732
rect 34724 41668 34740 41732
rect 34613 41652 34740 41668
rect 34613 41588 34660 41652
rect 34724 41588 34740 41652
rect 34613 41572 34740 41588
rect 34613 41508 34660 41572
rect 34724 41508 34740 41572
rect 34613 41492 34740 41508
rect 34613 41428 34660 41492
rect 34724 41428 34740 41492
rect 34613 41412 34740 41428
rect 34613 41348 34660 41412
rect 34724 41348 34740 41412
rect 34613 41332 34740 41348
rect 34613 41268 34660 41332
rect 34724 41268 34740 41332
rect 34613 41252 34740 41268
rect 34613 41188 34660 41252
rect 34724 41188 34740 41252
rect 34613 41172 34740 41188
rect 28294 41092 28421 41108
rect 28294 41028 28341 41092
rect 28405 41028 28421 41092
rect 28294 41012 28421 41028
rect 28294 40888 28398 41012
rect 28294 40872 28421 40888
rect 28294 40808 28341 40872
rect 28405 40808 28421 40872
rect 28294 40792 28421 40808
rect 21975 40712 22102 40728
rect 21975 40648 22022 40712
rect 22086 40648 22102 40712
rect 21975 40632 22102 40648
rect 21975 40568 22022 40632
rect 22086 40568 22102 40632
rect 21975 40552 22102 40568
rect 21975 40488 22022 40552
rect 22086 40488 22102 40552
rect 21975 40472 22102 40488
rect 21975 40408 22022 40472
rect 22086 40408 22102 40472
rect 21975 40392 22102 40408
rect 21975 40328 22022 40392
rect 22086 40328 22102 40392
rect 21975 40312 22102 40328
rect 21975 40248 22022 40312
rect 22086 40248 22102 40312
rect 21975 40232 22102 40248
rect 21975 40168 22022 40232
rect 22086 40168 22102 40232
rect 21975 40152 22102 40168
rect 21975 40088 22022 40152
rect 22086 40088 22102 40152
rect 21975 40072 22102 40088
rect 21975 40008 22022 40072
rect 22086 40008 22102 40072
rect 21975 39992 22102 40008
rect 21975 39928 22022 39992
rect 22086 39928 22102 39992
rect 21975 39912 22102 39928
rect 21975 39848 22022 39912
rect 22086 39848 22102 39912
rect 21975 39832 22102 39848
rect 21975 39768 22022 39832
rect 22086 39768 22102 39832
rect 21975 39752 22102 39768
rect 21975 39688 22022 39752
rect 22086 39688 22102 39752
rect 21975 39672 22102 39688
rect 21975 39608 22022 39672
rect 22086 39608 22102 39672
rect 21975 39592 22102 39608
rect 21975 39528 22022 39592
rect 22086 39528 22102 39592
rect 21975 39512 22102 39528
rect 21975 39448 22022 39512
rect 22086 39448 22102 39512
rect 21975 39432 22102 39448
rect 21975 39368 22022 39432
rect 22086 39368 22102 39432
rect 21975 39352 22102 39368
rect 21975 39288 22022 39352
rect 22086 39288 22102 39352
rect 21975 39272 22102 39288
rect 21975 39208 22022 39272
rect 22086 39208 22102 39272
rect 21975 39192 22102 39208
rect 21975 39128 22022 39192
rect 22086 39128 22102 39192
rect 21975 39112 22102 39128
rect 21975 39048 22022 39112
rect 22086 39048 22102 39112
rect 21975 39032 22102 39048
rect 21975 38968 22022 39032
rect 22086 38968 22102 39032
rect 21975 38952 22102 38968
rect 21975 38888 22022 38952
rect 22086 38888 22102 38952
rect 21975 38872 22102 38888
rect 21975 38808 22022 38872
rect 22086 38808 22102 38872
rect 21975 38792 22102 38808
rect 21975 38728 22022 38792
rect 22086 38728 22102 38792
rect 21975 38712 22102 38728
rect 21975 38648 22022 38712
rect 22086 38648 22102 38712
rect 21975 38632 22102 38648
rect 21975 38568 22022 38632
rect 22086 38568 22102 38632
rect 21975 38552 22102 38568
rect 21975 38488 22022 38552
rect 22086 38488 22102 38552
rect 21975 38472 22102 38488
rect 21975 38408 22022 38472
rect 22086 38408 22102 38472
rect 21975 38392 22102 38408
rect 21975 38328 22022 38392
rect 22086 38328 22102 38392
rect 21975 38312 22102 38328
rect 21975 38248 22022 38312
rect 22086 38248 22102 38312
rect 21975 38232 22102 38248
rect 21975 38168 22022 38232
rect 22086 38168 22102 38232
rect 21975 38152 22102 38168
rect 21975 38088 22022 38152
rect 22086 38088 22102 38152
rect 21975 38072 22102 38088
rect 21975 38008 22022 38072
rect 22086 38008 22102 38072
rect 21975 37992 22102 38008
rect 21975 37928 22022 37992
rect 22086 37928 22102 37992
rect 21975 37912 22102 37928
rect 21975 37848 22022 37912
rect 22086 37848 22102 37912
rect 21975 37832 22102 37848
rect 21975 37768 22022 37832
rect 22086 37768 22102 37832
rect 21975 37752 22102 37768
rect 21975 37688 22022 37752
rect 22086 37688 22102 37752
rect 21975 37672 22102 37688
rect 21975 37608 22022 37672
rect 22086 37608 22102 37672
rect 21975 37592 22102 37608
rect 21975 37528 22022 37592
rect 22086 37528 22102 37592
rect 21975 37512 22102 37528
rect 21975 37448 22022 37512
rect 22086 37448 22102 37512
rect 21975 37432 22102 37448
rect 21975 37368 22022 37432
rect 22086 37368 22102 37432
rect 21975 37352 22102 37368
rect 21975 37288 22022 37352
rect 22086 37288 22102 37352
rect 21975 37272 22102 37288
rect 21975 37208 22022 37272
rect 22086 37208 22102 37272
rect 21975 37192 22102 37208
rect 21975 37128 22022 37192
rect 22086 37128 22102 37192
rect 21975 37112 22102 37128
rect 21975 37048 22022 37112
rect 22086 37048 22102 37112
rect 21975 37032 22102 37048
rect 21975 36968 22022 37032
rect 22086 36968 22102 37032
rect 21975 36952 22102 36968
rect 21975 36888 22022 36952
rect 22086 36888 22102 36952
rect 21975 36872 22102 36888
rect 21975 36808 22022 36872
rect 22086 36808 22102 36872
rect 21975 36792 22102 36808
rect 21975 36728 22022 36792
rect 22086 36728 22102 36792
rect 21975 36712 22102 36728
rect 21975 36648 22022 36712
rect 22086 36648 22102 36712
rect 21975 36632 22102 36648
rect 21975 36568 22022 36632
rect 22086 36568 22102 36632
rect 21975 36552 22102 36568
rect 21975 36488 22022 36552
rect 22086 36488 22102 36552
rect 21975 36472 22102 36488
rect 21975 36408 22022 36472
rect 22086 36408 22102 36472
rect 21975 36392 22102 36408
rect 21975 36328 22022 36392
rect 22086 36328 22102 36392
rect 21975 36312 22102 36328
rect 21975 36248 22022 36312
rect 22086 36248 22102 36312
rect 21975 36232 22102 36248
rect 21975 36168 22022 36232
rect 22086 36168 22102 36232
rect 21975 36152 22102 36168
rect 21975 36088 22022 36152
rect 22086 36088 22102 36152
rect 21975 36072 22102 36088
rect 21975 36008 22022 36072
rect 22086 36008 22102 36072
rect 21975 35992 22102 36008
rect 21975 35928 22022 35992
rect 22086 35928 22102 35992
rect 21975 35912 22102 35928
rect 21975 35848 22022 35912
rect 22086 35848 22102 35912
rect 21975 35832 22102 35848
rect 21975 35768 22022 35832
rect 22086 35768 22102 35832
rect 21975 35752 22102 35768
rect 21975 35688 22022 35752
rect 22086 35688 22102 35752
rect 21975 35672 22102 35688
rect 21975 35608 22022 35672
rect 22086 35608 22102 35672
rect 21975 35592 22102 35608
rect 21975 35528 22022 35592
rect 22086 35528 22102 35592
rect 21975 35512 22102 35528
rect 21975 35448 22022 35512
rect 22086 35448 22102 35512
rect 21975 35432 22102 35448
rect 21975 35368 22022 35432
rect 22086 35368 22102 35432
rect 21975 35352 22102 35368
rect 21975 35288 22022 35352
rect 22086 35288 22102 35352
rect 21975 35272 22102 35288
rect 21975 35208 22022 35272
rect 22086 35208 22102 35272
rect 21975 35192 22102 35208
rect 21975 35128 22022 35192
rect 22086 35128 22102 35192
rect 21975 35112 22102 35128
rect 21975 35048 22022 35112
rect 22086 35048 22102 35112
rect 21975 35032 22102 35048
rect 21975 34968 22022 35032
rect 22086 34968 22102 35032
rect 21975 34952 22102 34968
rect 21975 34888 22022 34952
rect 22086 34888 22102 34952
rect 21975 34872 22102 34888
rect 15656 34792 15783 34808
rect 15656 34728 15703 34792
rect 15767 34728 15783 34792
rect 15656 34712 15783 34728
rect 15656 34588 15760 34712
rect 15656 34572 15783 34588
rect 15656 34508 15703 34572
rect 15767 34508 15783 34572
rect 15656 34492 15783 34508
rect 9337 34412 9464 34428
rect 9337 34348 9384 34412
rect 9448 34348 9464 34412
rect 9337 34332 9464 34348
rect 9337 34268 9384 34332
rect 9448 34268 9464 34332
rect 9337 34252 9464 34268
rect 9337 34188 9384 34252
rect 9448 34188 9464 34252
rect 9337 34172 9464 34188
rect 9337 34108 9384 34172
rect 9448 34108 9464 34172
rect 9337 34092 9464 34108
rect 9337 34028 9384 34092
rect 9448 34028 9464 34092
rect 9337 34012 9464 34028
rect 9337 33948 9384 34012
rect 9448 33948 9464 34012
rect 9337 33932 9464 33948
rect 9337 33868 9384 33932
rect 9448 33868 9464 33932
rect 9337 33852 9464 33868
rect 9337 33788 9384 33852
rect 9448 33788 9464 33852
rect 9337 33772 9464 33788
rect 9337 33708 9384 33772
rect 9448 33708 9464 33772
rect 9337 33692 9464 33708
rect 9337 33628 9384 33692
rect 9448 33628 9464 33692
rect 9337 33612 9464 33628
rect 9337 33548 9384 33612
rect 9448 33548 9464 33612
rect 9337 33532 9464 33548
rect 9337 33468 9384 33532
rect 9448 33468 9464 33532
rect 9337 33452 9464 33468
rect 9337 33388 9384 33452
rect 9448 33388 9464 33452
rect 9337 33372 9464 33388
rect 9337 33308 9384 33372
rect 9448 33308 9464 33372
rect 9337 33292 9464 33308
rect 9337 33228 9384 33292
rect 9448 33228 9464 33292
rect 9337 33212 9464 33228
rect 9337 33148 9384 33212
rect 9448 33148 9464 33212
rect 9337 33132 9464 33148
rect 9337 33068 9384 33132
rect 9448 33068 9464 33132
rect 9337 33052 9464 33068
rect 9337 32988 9384 33052
rect 9448 32988 9464 33052
rect 9337 32972 9464 32988
rect 9337 32908 9384 32972
rect 9448 32908 9464 32972
rect 9337 32892 9464 32908
rect 9337 32828 9384 32892
rect 9448 32828 9464 32892
rect 9337 32812 9464 32828
rect 9337 32748 9384 32812
rect 9448 32748 9464 32812
rect 9337 32732 9464 32748
rect 9337 32668 9384 32732
rect 9448 32668 9464 32732
rect 9337 32652 9464 32668
rect 9337 32588 9384 32652
rect 9448 32588 9464 32652
rect 9337 32572 9464 32588
rect 9337 32508 9384 32572
rect 9448 32508 9464 32572
rect 9337 32492 9464 32508
rect 9337 32428 9384 32492
rect 9448 32428 9464 32492
rect 9337 32412 9464 32428
rect 9337 32348 9384 32412
rect 9448 32348 9464 32412
rect 9337 32332 9464 32348
rect 9337 32268 9384 32332
rect 9448 32268 9464 32332
rect 9337 32252 9464 32268
rect 9337 32188 9384 32252
rect 9448 32188 9464 32252
rect 9337 32172 9464 32188
rect 9337 32108 9384 32172
rect 9448 32108 9464 32172
rect 9337 32092 9464 32108
rect 9337 32028 9384 32092
rect 9448 32028 9464 32092
rect 9337 32012 9464 32028
rect 9337 31948 9384 32012
rect 9448 31948 9464 32012
rect 9337 31932 9464 31948
rect 9337 31868 9384 31932
rect 9448 31868 9464 31932
rect 9337 31852 9464 31868
rect 9337 31788 9384 31852
rect 9448 31788 9464 31852
rect 9337 31772 9464 31788
rect 9337 31708 9384 31772
rect 9448 31708 9464 31772
rect 9337 31692 9464 31708
rect 9337 31628 9384 31692
rect 9448 31628 9464 31692
rect 9337 31612 9464 31628
rect 9337 31548 9384 31612
rect 9448 31548 9464 31612
rect 9337 31532 9464 31548
rect 9337 31468 9384 31532
rect 9448 31468 9464 31532
rect 9337 31452 9464 31468
rect 9337 31388 9384 31452
rect 9448 31388 9464 31452
rect 9337 31372 9464 31388
rect 9337 31308 9384 31372
rect 9448 31308 9464 31372
rect 9337 31292 9464 31308
rect 9337 31228 9384 31292
rect 9448 31228 9464 31292
rect 9337 31212 9464 31228
rect 9337 31148 9384 31212
rect 9448 31148 9464 31212
rect 9337 31132 9464 31148
rect 9337 31068 9384 31132
rect 9448 31068 9464 31132
rect 9337 31052 9464 31068
rect 9337 30988 9384 31052
rect 9448 30988 9464 31052
rect 9337 30972 9464 30988
rect 9337 30908 9384 30972
rect 9448 30908 9464 30972
rect 9337 30892 9464 30908
rect 9337 30828 9384 30892
rect 9448 30828 9464 30892
rect 9337 30812 9464 30828
rect 9337 30748 9384 30812
rect 9448 30748 9464 30812
rect 9337 30732 9464 30748
rect 9337 30668 9384 30732
rect 9448 30668 9464 30732
rect 9337 30652 9464 30668
rect 9337 30588 9384 30652
rect 9448 30588 9464 30652
rect 9337 30572 9464 30588
rect 9337 30508 9384 30572
rect 9448 30508 9464 30572
rect 9337 30492 9464 30508
rect 9337 30428 9384 30492
rect 9448 30428 9464 30492
rect 9337 30412 9464 30428
rect 9337 30348 9384 30412
rect 9448 30348 9464 30412
rect 9337 30332 9464 30348
rect 9337 30268 9384 30332
rect 9448 30268 9464 30332
rect 9337 30252 9464 30268
rect 9337 30188 9384 30252
rect 9448 30188 9464 30252
rect 9337 30172 9464 30188
rect 9337 30108 9384 30172
rect 9448 30108 9464 30172
rect 9337 30092 9464 30108
rect 9337 30028 9384 30092
rect 9448 30028 9464 30092
rect 9337 30012 9464 30028
rect 9337 29948 9384 30012
rect 9448 29948 9464 30012
rect 9337 29932 9464 29948
rect 9337 29868 9384 29932
rect 9448 29868 9464 29932
rect 9337 29852 9464 29868
rect 9337 29788 9384 29852
rect 9448 29788 9464 29852
rect 9337 29772 9464 29788
rect 9337 29708 9384 29772
rect 9448 29708 9464 29772
rect 9337 29692 9464 29708
rect 9337 29628 9384 29692
rect 9448 29628 9464 29692
rect 9337 29612 9464 29628
rect 9337 29548 9384 29612
rect 9448 29548 9464 29612
rect 9337 29532 9464 29548
rect 9337 29468 9384 29532
rect 9448 29468 9464 29532
rect 9337 29452 9464 29468
rect 9337 29388 9384 29452
rect 9448 29388 9464 29452
rect 9337 29372 9464 29388
rect 9337 29308 9384 29372
rect 9448 29308 9464 29372
rect 9337 29292 9464 29308
rect 9337 29228 9384 29292
rect 9448 29228 9464 29292
rect 9337 29212 9464 29228
rect 9337 29148 9384 29212
rect 9448 29148 9464 29212
rect 9337 29132 9464 29148
rect 9337 29068 9384 29132
rect 9448 29068 9464 29132
rect 9337 29052 9464 29068
rect 9337 28988 9384 29052
rect 9448 28988 9464 29052
rect 9337 28972 9464 28988
rect 9337 28908 9384 28972
rect 9448 28908 9464 28972
rect 9337 28892 9464 28908
rect 9337 28828 9384 28892
rect 9448 28828 9464 28892
rect 9337 28812 9464 28828
rect 9337 28748 9384 28812
rect 9448 28748 9464 28812
rect 9337 28732 9464 28748
rect 9337 28668 9384 28732
rect 9448 28668 9464 28732
rect 9337 28652 9464 28668
rect 9337 28588 9384 28652
rect 9448 28588 9464 28652
rect 9337 28572 9464 28588
rect 3018 28492 3145 28508
rect 3018 28428 3065 28492
rect 3129 28428 3145 28492
rect 3018 28412 3145 28428
rect 3018 28288 3122 28412
rect 3018 28272 3145 28288
rect 3018 28208 3065 28272
rect 3129 28208 3145 28272
rect 3018 28192 3145 28208
rect -3301 28112 -3174 28128
rect -3301 28048 -3254 28112
rect -3190 28048 -3174 28112
rect -3301 28032 -3174 28048
rect -3301 27968 -3254 28032
rect -3190 27968 -3174 28032
rect -3301 27952 -3174 27968
rect -3301 27888 -3254 27952
rect -3190 27888 -3174 27952
rect -3301 27872 -3174 27888
rect -3301 27808 -3254 27872
rect -3190 27808 -3174 27872
rect -3301 27792 -3174 27808
rect -3301 27728 -3254 27792
rect -3190 27728 -3174 27792
rect -3301 27712 -3174 27728
rect -3301 27648 -3254 27712
rect -3190 27648 -3174 27712
rect -3301 27632 -3174 27648
rect -3301 27568 -3254 27632
rect -3190 27568 -3174 27632
rect -3301 27552 -3174 27568
rect -3301 27488 -3254 27552
rect -3190 27488 -3174 27552
rect -3301 27472 -3174 27488
rect -3301 27408 -3254 27472
rect -3190 27408 -3174 27472
rect -3301 27392 -3174 27408
rect -3301 27328 -3254 27392
rect -3190 27328 -3174 27392
rect -3301 27312 -3174 27328
rect -3301 27248 -3254 27312
rect -3190 27248 -3174 27312
rect -3301 27232 -3174 27248
rect -3301 27168 -3254 27232
rect -3190 27168 -3174 27232
rect -3301 27152 -3174 27168
rect -3301 27088 -3254 27152
rect -3190 27088 -3174 27152
rect -3301 27072 -3174 27088
rect -3301 27008 -3254 27072
rect -3190 27008 -3174 27072
rect -3301 26992 -3174 27008
rect -3301 26928 -3254 26992
rect -3190 26928 -3174 26992
rect -3301 26912 -3174 26928
rect -3301 26848 -3254 26912
rect -3190 26848 -3174 26912
rect -3301 26832 -3174 26848
rect -3301 26768 -3254 26832
rect -3190 26768 -3174 26832
rect -3301 26752 -3174 26768
rect -3301 26688 -3254 26752
rect -3190 26688 -3174 26752
rect -3301 26672 -3174 26688
rect -3301 26608 -3254 26672
rect -3190 26608 -3174 26672
rect -3301 26592 -3174 26608
rect -3301 26528 -3254 26592
rect -3190 26528 -3174 26592
rect -3301 26512 -3174 26528
rect -3301 26448 -3254 26512
rect -3190 26448 -3174 26512
rect -3301 26432 -3174 26448
rect -3301 26368 -3254 26432
rect -3190 26368 -3174 26432
rect -3301 26352 -3174 26368
rect -3301 26288 -3254 26352
rect -3190 26288 -3174 26352
rect -3301 26272 -3174 26288
rect -3301 26208 -3254 26272
rect -3190 26208 -3174 26272
rect -3301 26192 -3174 26208
rect -3301 26128 -3254 26192
rect -3190 26128 -3174 26192
rect -3301 26112 -3174 26128
rect -3301 26048 -3254 26112
rect -3190 26048 -3174 26112
rect -3301 26032 -3174 26048
rect -3301 25968 -3254 26032
rect -3190 25968 -3174 26032
rect -3301 25952 -3174 25968
rect -3301 25888 -3254 25952
rect -3190 25888 -3174 25952
rect -3301 25872 -3174 25888
rect -3301 25808 -3254 25872
rect -3190 25808 -3174 25872
rect -3301 25792 -3174 25808
rect -3301 25728 -3254 25792
rect -3190 25728 -3174 25792
rect -3301 25712 -3174 25728
rect -3301 25648 -3254 25712
rect -3190 25648 -3174 25712
rect -3301 25632 -3174 25648
rect -3301 25568 -3254 25632
rect -3190 25568 -3174 25632
rect -3301 25552 -3174 25568
rect -3301 25488 -3254 25552
rect -3190 25488 -3174 25552
rect -3301 25472 -3174 25488
rect -3301 25408 -3254 25472
rect -3190 25408 -3174 25472
rect -3301 25392 -3174 25408
rect -3301 25328 -3254 25392
rect -3190 25328 -3174 25392
rect -3301 25312 -3174 25328
rect -3301 25248 -3254 25312
rect -3190 25248 -3174 25312
rect -3301 25232 -3174 25248
rect -3301 25168 -3254 25232
rect -3190 25168 -3174 25232
rect -3301 25152 -3174 25168
rect -3301 25088 -3254 25152
rect -3190 25088 -3174 25152
rect -3301 25072 -3174 25088
rect -3301 25008 -3254 25072
rect -3190 25008 -3174 25072
rect -3301 24992 -3174 25008
rect -3301 24928 -3254 24992
rect -3190 24928 -3174 24992
rect -3301 24912 -3174 24928
rect -3301 24848 -3254 24912
rect -3190 24848 -3174 24912
rect -3301 24832 -3174 24848
rect -3301 24768 -3254 24832
rect -3190 24768 -3174 24832
rect -3301 24752 -3174 24768
rect -3301 24688 -3254 24752
rect -3190 24688 -3174 24752
rect -3301 24672 -3174 24688
rect -3301 24608 -3254 24672
rect -3190 24608 -3174 24672
rect -3301 24592 -3174 24608
rect -3301 24528 -3254 24592
rect -3190 24528 -3174 24592
rect -3301 24512 -3174 24528
rect -3301 24448 -3254 24512
rect -3190 24448 -3174 24512
rect -3301 24432 -3174 24448
rect -3301 24368 -3254 24432
rect -3190 24368 -3174 24432
rect -3301 24352 -3174 24368
rect -3301 24288 -3254 24352
rect -3190 24288 -3174 24352
rect -3301 24272 -3174 24288
rect -3301 24208 -3254 24272
rect -3190 24208 -3174 24272
rect -3301 24192 -3174 24208
rect -3301 24128 -3254 24192
rect -3190 24128 -3174 24192
rect -3301 24112 -3174 24128
rect -3301 24048 -3254 24112
rect -3190 24048 -3174 24112
rect -3301 24032 -3174 24048
rect -3301 23968 -3254 24032
rect -3190 23968 -3174 24032
rect -3301 23952 -3174 23968
rect -3301 23888 -3254 23952
rect -3190 23888 -3174 23952
rect -3301 23872 -3174 23888
rect -3301 23808 -3254 23872
rect -3190 23808 -3174 23872
rect -3301 23792 -3174 23808
rect -3301 23728 -3254 23792
rect -3190 23728 -3174 23792
rect -3301 23712 -3174 23728
rect -3301 23648 -3254 23712
rect -3190 23648 -3174 23712
rect -3301 23632 -3174 23648
rect -3301 23568 -3254 23632
rect -3190 23568 -3174 23632
rect -3301 23552 -3174 23568
rect -3301 23488 -3254 23552
rect -3190 23488 -3174 23552
rect -3301 23472 -3174 23488
rect -3301 23408 -3254 23472
rect -3190 23408 -3174 23472
rect -3301 23392 -3174 23408
rect -3301 23328 -3254 23392
rect -3190 23328 -3174 23392
rect -3301 23312 -3174 23328
rect -3301 23248 -3254 23312
rect -3190 23248 -3174 23312
rect -3301 23232 -3174 23248
rect -3301 23168 -3254 23232
rect -3190 23168 -3174 23232
rect -3301 23152 -3174 23168
rect -3301 23088 -3254 23152
rect -3190 23088 -3174 23152
rect -3301 23072 -3174 23088
rect -3301 23008 -3254 23072
rect -3190 23008 -3174 23072
rect -3301 22992 -3174 23008
rect -3301 22928 -3254 22992
rect -3190 22928 -3174 22992
rect -3301 22912 -3174 22928
rect -3301 22848 -3254 22912
rect -3190 22848 -3174 22912
rect -3301 22832 -3174 22848
rect -3301 22768 -3254 22832
rect -3190 22768 -3174 22832
rect -3301 22752 -3174 22768
rect -3301 22688 -3254 22752
rect -3190 22688 -3174 22752
rect -3301 22672 -3174 22688
rect -3301 22608 -3254 22672
rect -3190 22608 -3174 22672
rect -3301 22592 -3174 22608
rect -3301 22528 -3254 22592
rect -3190 22528 -3174 22592
rect -3301 22512 -3174 22528
rect -3301 22448 -3254 22512
rect -3190 22448 -3174 22512
rect -3301 22432 -3174 22448
rect -3301 22368 -3254 22432
rect -3190 22368 -3174 22432
rect -3301 22352 -3174 22368
rect -3301 22288 -3254 22352
rect -3190 22288 -3174 22352
rect -3301 22272 -3174 22288
rect -9620 22192 -9493 22208
rect -9620 22128 -9573 22192
rect -9509 22128 -9493 22192
rect -9620 22112 -9493 22128
rect -9620 21988 -9516 22112
rect -9620 21972 -9493 21988
rect -9620 21908 -9573 21972
rect -9509 21908 -9493 21972
rect -9620 21892 -9493 21908
rect -15939 21812 -15812 21828
rect -15939 21748 -15892 21812
rect -15828 21748 -15812 21812
rect -15939 21732 -15812 21748
rect -15939 21668 -15892 21732
rect -15828 21668 -15812 21732
rect -15939 21652 -15812 21668
rect -15939 21588 -15892 21652
rect -15828 21588 -15812 21652
rect -15939 21572 -15812 21588
rect -15939 21508 -15892 21572
rect -15828 21508 -15812 21572
rect -15939 21492 -15812 21508
rect -15939 21428 -15892 21492
rect -15828 21428 -15812 21492
rect -15939 21412 -15812 21428
rect -15939 21348 -15892 21412
rect -15828 21348 -15812 21412
rect -15939 21332 -15812 21348
rect -15939 21268 -15892 21332
rect -15828 21268 -15812 21332
rect -15939 21252 -15812 21268
rect -15939 21188 -15892 21252
rect -15828 21188 -15812 21252
rect -15939 21172 -15812 21188
rect -15939 21108 -15892 21172
rect -15828 21108 -15812 21172
rect -15939 21092 -15812 21108
rect -15939 21028 -15892 21092
rect -15828 21028 -15812 21092
rect -15939 21012 -15812 21028
rect -15939 20948 -15892 21012
rect -15828 20948 -15812 21012
rect -15939 20932 -15812 20948
rect -15939 20868 -15892 20932
rect -15828 20868 -15812 20932
rect -15939 20852 -15812 20868
rect -15939 20788 -15892 20852
rect -15828 20788 -15812 20852
rect -15939 20772 -15812 20788
rect -15939 20708 -15892 20772
rect -15828 20708 -15812 20772
rect -15939 20692 -15812 20708
rect -15939 20628 -15892 20692
rect -15828 20628 -15812 20692
rect -15939 20612 -15812 20628
rect -15939 20548 -15892 20612
rect -15828 20548 -15812 20612
rect -15939 20532 -15812 20548
rect -15939 20468 -15892 20532
rect -15828 20468 -15812 20532
rect -15939 20452 -15812 20468
rect -15939 20388 -15892 20452
rect -15828 20388 -15812 20452
rect -15939 20372 -15812 20388
rect -15939 20308 -15892 20372
rect -15828 20308 -15812 20372
rect -15939 20292 -15812 20308
rect -15939 20228 -15892 20292
rect -15828 20228 -15812 20292
rect -15939 20212 -15812 20228
rect -15939 20148 -15892 20212
rect -15828 20148 -15812 20212
rect -15939 20132 -15812 20148
rect -15939 20068 -15892 20132
rect -15828 20068 -15812 20132
rect -15939 20052 -15812 20068
rect -15939 19988 -15892 20052
rect -15828 19988 -15812 20052
rect -15939 19972 -15812 19988
rect -15939 19908 -15892 19972
rect -15828 19908 -15812 19972
rect -15939 19892 -15812 19908
rect -15939 19828 -15892 19892
rect -15828 19828 -15812 19892
rect -15939 19812 -15812 19828
rect -15939 19748 -15892 19812
rect -15828 19748 -15812 19812
rect -15939 19732 -15812 19748
rect -15939 19668 -15892 19732
rect -15828 19668 -15812 19732
rect -15939 19652 -15812 19668
rect -15939 19588 -15892 19652
rect -15828 19588 -15812 19652
rect -15939 19572 -15812 19588
rect -15939 19508 -15892 19572
rect -15828 19508 -15812 19572
rect -15939 19492 -15812 19508
rect -15939 19428 -15892 19492
rect -15828 19428 -15812 19492
rect -15939 19412 -15812 19428
rect -15939 19348 -15892 19412
rect -15828 19348 -15812 19412
rect -15939 19332 -15812 19348
rect -15939 19268 -15892 19332
rect -15828 19268 -15812 19332
rect -15939 19252 -15812 19268
rect -15939 19188 -15892 19252
rect -15828 19188 -15812 19252
rect -15939 19172 -15812 19188
rect -15939 19108 -15892 19172
rect -15828 19108 -15812 19172
rect -15939 19092 -15812 19108
rect -15939 19028 -15892 19092
rect -15828 19028 -15812 19092
rect -15939 19012 -15812 19028
rect -15939 18948 -15892 19012
rect -15828 18948 -15812 19012
rect -15939 18932 -15812 18948
rect -15939 18868 -15892 18932
rect -15828 18868 -15812 18932
rect -15939 18852 -15812 18868
rect -15939 18788 -15892 18852
rect -15828 18788 -15812 18852
rect -15939 18772 -15812 18788
rect -15939 18708 -15892 18772
rect -15828 18708 -15812 18772
rect -15939 18692 -15812 18708
rect -15939 18628 -15892 18692
rect -15828 18628 -15812 18692
rect -15939 18612 -15812 18628
rect -15939 18548 -15892 18612
rect -15828 18548 -15812 18612
rect -15939 18532 -15812 18548
rect -15939 18468 -15892 18532
rect -15828 18468 -15812 18532
rect -15939 18452 -15812 18468
rect -15939 18388 -15892 18452
rect -15828 18388 -15812 18452
rect -15939 18372 -15812 18388
rect -15939 18308 -15892 18372
rect -15828 18308 -15812 18372
rect -15939 18292 -15812 18308
rect -15939 18228 -15892 18292
rect -15828 18228 -15812 18292
rect -15939 18212 -15812 18228
rect -15939 18148 -15892 18212
rect -15828 18148 -15812 18212
rect -15939 18132 -15812 18148
rect -15939 18068 -15892 18132
rect -15828 18068 -15812 18132
rect -15939 18052 -15812 18068
rect -15939 17988 -15892 18052
rect -15828 17988 -15812 18052
rect -15939 17972 -15812 17988
rect -15939 17908 -15892 17972
rect -15828 17908 -15812 17972
rect -15939 17892 -15812 17908
rect -15939 17828 -15892 17892
rect -15828 17828 -15812 17892
rect -15939 17812 -15812 17828
rect -15939 17748 -15892 17812
rect -15828 17748 -15812 17812
rect -15939 17732 -15812 17748
rect -15939 17668 -15892 17732
rect -15828 17668 -15812 17732
rect -15939 17652 -15812 17668
rect -15939 17588 -15892 17652
rect -15828 17588 -15812 17652
rect -15939 17572 -15812 17588
rect -15939 17508 -15892 17572
rect -15828 17508 -15812 17572
rect -15939 17492 -15812 17508
rect -15939 17428 -15892 17492
rect -15828 17428 -15812 17492
rect -15939 17412 -15812 17428
rect -15939 17348 -15892 17412
rect -15828 17348 -15812 17412
rect -15939 17332 -15812 17348
rect -15939 17268 -15892 17332
rect -15828 17268 -15812 17332
rect -15939 17252 -15812 17268
rect -15939 17188 -15892 17252
rect -15828 17188 -15812 17252
rect -15939 17172 -15812 17188
rect -15939 17108 -15892 17172
rect -15828 17108 -15812 17172
rect -15939 17092 -15812 17108
rect -15939 17028 -15892 17092
rect -15828 17028 -15812 17092
rect -15939 17012 -15812 17028
rect -15939 16948 -15892 17012
rect -15828 16948 -15812 17012
rect -15939 16932 -15812 16948
rect -15939 16868 -15892 16932
rect -15828 16868 -15812 16932
rect -15939 16852 -15812 16868
rect -15939 16788 -15892 16852
rect -15828 16788 -15812 16852
rect -15939 16772 -15812 16788
rect -15939 16708 -15892 16772
rect -15828 16708 -15812 16772
rect -15939 16692 -15812 16708
rect -15939 16628 -15892 16692
rect -15828 16628 -15812 16692
rect -15939 16612 -15812 16628
rect -15939 16548 -15892 16612
rect -15828 16548 -15812 16612
rect -15939 16532 -15812 16548
rect -15939 16468 -15892 16532
rect -15828 16468 -15812 16532
rect -15939 16452 -15812 16468
rect -15939 16388 -15892 16452
rect -15828 16388 -15812 16452
rect -15939 16372 -15812 16388
rect -15939 16308 -15892 16372
rect -15828 16308 -15812 16372
rect -15939 16292 -15812 16308
rect -15939 16228 -15892 16292
rect -15828 16228 -15812 16292
rect -15939 16212 -15812 16228
rect -15939 16148 -15892 16212
rect -15828 16148 -15812 16212
rect -15939 16132 -15812 16148
rect -15939 16068 -15892 16132
rect -15828 16068 -15812 16132
rect -15939 16052 -15812 16068
rect -15939 15988 -15892 16052
rect -15828 15988 -15812 16052
rect -15939 15972 -15812 15988
rect -22258 15892 -22131 15908
rect -22258 15828 -22211 15892
rect -22147 15828 -22131 15892
rect -22258 15812 -22131 15828
rect -22258 15688 -22154 15812
rect -22258 15672 -22131 15688
rect -22258 15608 -22211 15672
rect -22147 15608 -22131 15672
rect -22258 15592 -22131 15608
rect -28577 15512 -28450 15528
rect -28577 15448 -28530 15512
rect -28466 15448 -28450 15512
rect -28577 15432 -28450 15448
rect -28577 15368 -28530 15432
rect -28466 15368 -28450 15432
rect -28577 15352 -28450 15368
rect -28577 15288 -28530 15352
rect -28466 15288 -28450 15352
rect -28577 15272 -28450 15288
rect -28577 15208 -28530 15272
rect -28466 15208 -28450 15272
rect -28577 15192 -28450 15208
rect -28577 15128 -28530 15192
rect -28466 15128 -28450 15192
rect -28577 15112 -28450 15128
rect -28577 15048 -28530 15112
rect -28466 15048 -28450 15112
rect -28577 15032 -28450 15048
rect -28577 14968 -28530 15032
rect -28466 14968 -28450 15032
rect -28577 14952 -28450 14968
rect -28577 14888 -28530 14952
rect -28466 14888 -28450 14952
rect -28577 14872 -28450 14888
rect -28577 14808 -28530 14872
rect -28466 14808 -28450 14872
rect -28577 14792 -28450 14808
rect -28577 14728 -28530 14792
rect -28466 14728 -28450 14792
rect -28577 14712 -28450 14728
rect -28577 14648 -28530 14712
rect -28466 14648 -28450 14712
rect -28577 14632 -28450 14648
rect -28577 14568 -28530 14632
rect -28466 14568 -28450 14632
rect -28577 14552 -28450 14568
rect -28577 14488 -28530 14552
rect -28466 14488 -28450 14552
rect -28577 14472 -28450 14488
rect -28577 14408 -28530 14472
rect -28466 14408 -28450 14472
rect -28577 14392 -28450 14408
rect -28577 14328 -28530 14392
rect -28466 14328 -28450 14392
rect -28577 14312 -28450 14328
rect -28577 14248 -28530 14312
rect -28466 14248 -28450 14312
rect -28577 14232 -28450 14248
rect -28577 14168 -28530 14232
rect -28466 14168 -28450 14232
rect -28577 14152 -28450 14168
rect -28577 14088 -28530 14152
rect -28466 14088 -28450 14152
rect -28577 14072 -28450 14088
rect -28577 14008 -28530 14072
rect -28466 14008 -28450 14072
rect -28577 13992 -28450 14008
rect -28577 13928 -28530 13992
rect -28466 13928 -28450 13992
rect -28577 13912 -28450 13928
rect -28577 13848 -28530 13912
rect -28466 13848 -28450 13912
rect -28577 13832 -28450 13848
rect -28577 13768 -28530 13832
rect -28466 13768 -28450 13832
rect -28577 13752 -28450 13768
rect -28577 13688 -28530 13752
rect -28466 13688 -28450 13752
rect -28577 13672 -28450 13688
rect -28577 13608 -28530 13672
rect -28466 13608 -28450 13672
rect -28577 13592 -28450 13608
rect -28577 13528 -28530 13592
rect -28466 13528 -28450 13592
rect -28577 13512 -28450 13528
rect -28577 13448 -28530 13512
rect -28466 13448 -28450 13512
rect -28577 13432 -28450 13448
rect -28577 13368 -28530 13432
rect -28466 13368 -28450 13432
rect -28577 13352 -28450 13368
rect -28577 13288 -28530 13352
rect -28466 13288 -28450 13352
rect -28577 13272 -28450 13288
rect -28577 13208 -28530 13272
rect -28466 13208 -28450 13272
rect -28577 13192 -28450 13208
rect -28577 13128 -28530 13192
rect -28466 13128 -28450 13192
rect -28577 13112 -28450 13128
rect -28577 13048 -28530 13112
rect -28466 13048 -28450 13112
rect -28577 13032 -28450 13048
rect -28577 12968 -28530 13032
rect -28466 12968 -28450 13032
rect -28577 12952 -28450 12968
rect -28577 12888 -28530 12952
rect -28466 12888 -28450 12952
rect -28577 12872 -28450 12888
rect -28577 12808 -28530 12872
rect -28466 12808 -28450 12872
rect -28577 12792 -28450 12808
rect -28577 12728 -28530 12792
rect -28466 12728 -28450 12792
rect -28577 12712 -28450 12728
rect -28577 12648 -28530 12712
rect -28466 12648 -28450 12712
rect -28577 12632 -28450 12648
rect -28577 12568 -28530 12632
rect -28466 12568 -28450 12632
rect -28577 12552 -28450 12568
rect -28577 12488 -28530 12552
rect -28466 12488 -28450 12552
rect -28577 12472 -28450 12488
rect -28577 12408 -28530 12472
rect -28466 12408 -28450 12472
rect -28577 12392 -28450 12408
rect -28577 12328 -28530 12392
rect -28466 12328 -28450 12392
rect -28577 12312 -28450 12328
rect -28577 12248 -28530 12312
rect -28466 12248 -28450 12312
rect -28577 12232 -28450 12248
rect -28577 12168 -28530 12232
rect -28466 12168 -28450 12232
rect -28577 12152 -28450 12168
rect -28577 12088 -28530 12152
rect -28466 12088 -28450 12152
rect -28577 12072 -28450 12088
rect -28577 12008 -28530 12072
rect -28466 12008 -28450 12072
rect -28577 11992 -28450 12008
rect -28577 11928 -28530 11992
rect -28466 11928 -28450 11992
rect -28577 11912 -28450 11928
rect -28577 11848 -28530 11912
rect -28466 11848 -28450 11912
rect -28577 11832 -28450 11848
rect -28577 11768 -28530 11832
rect -28466 11768 -28450 11832
rect -28577 11752 -28450 11768
rect -28577 11688 -28530 11752
rect -28466 11688 -28450 11752
rect -28577 11672 -28450 11688
rect -28577 11608 -28530 11672
rect -28466 11608 -28450 11672
rect -28577 11592 -28450 11608
rect -28577 11528 -28530 11592
rect -28466 11528 -28450 11592
rect -28577 11512 -28450 11528
rect -28577 11448 -28530 11512
rect -28466 11448 -28450 11512
rect -28577 11432 -28450 11448
rect -28577 11368 -28530 11432
rect -28466 11368 -28450 11432
rect -28577 11352 -28450 11368
rect -28577 11288 -28530 11352
rect -28466 11288 -28450 11352
rect -28577 11272 -28450 11288
rect -28577 11208 -28530 11272
rect -28466 11208 -28450 11272
rect -28577 11192 -28450 11208
rect -28577 11128 -28530 11192
rect -28466 11128 -28450 11192
rect -28577 11112 -28450 11128
rect -28577 11048 -28530 11112
rect -28466 11048 -28450 11112
rect -28577 11032 -28450 11048
rect -28577 10968 -28530 11032
rect -28466 10968 -28450 11032
rect -28577 10952 -28450 10968
rect -28577 10888 -28530 10952
rect -28466 10888 -28450 10952
rect -28577 10872 -28450 10888
rect -28577 10808 -28530 10872
rect -28466 10808 -28450 10872
rect -28577 10792 -28450 10808
rect -28577 10728 -28530 10792
rect -28466 10728 -28450 10792
rect -28577 10712 -28450 10728
rect -28577 10648 -28530 10712
rect -28466 10648 -28450 10712
rect -28577 10632 -28450 10648
rect -28577 10568 -28530 10632
rect -28466 10568 -28450 10632
rect -28577 10552 -28450 10568
rect -28577 10488 -28530 10552
rect -28466 10488 -28450 10552
rect -28577 10472 -28450 10488
rect -28577 10408 -28530 10472
rect -28466 10408 -28450 10472
rect -28577 10392 -28450 10408
rect -28577 10328 -28530 10392
rect -28466 10328 -28450 10392
rect -28577 10312 -28450 10328
rect -28577 10248 -28530 10312
rect -28466 10248 -28450 10312
rect -28577 10232 -28450 10248
rect -28577 10168 -28530 10232
rect -28466 10168 -28450 10232
rect -28577 10152 -28450 10168
rect -28577 10088 -28530 10152
rect -28466 10088 -28450 10152
rect -28577 10072 -28450 10088
rect -28577 10008 -28530 10072
rect -28466 10008 -28450 10072
rect -28577 9992 -28450 10008
rect -28577 9928 -28530 9992
rect -28466 9928 -28450 9992
rect -28577 9912 -28450 9928
rect -28577 9848 -28530 9912
rect -28466 9848 -28450 9912
rect -28577 9832 -28450 9848
rect -28577 9768 -28530 9832
rect -28466 9768 -28450 9832
rect -28577 9752 -28450 9768
rect -28577 9688 -28530 9752
rect -28466 9688 -28450 9752
rect -28577 9672 -28450 9688
rect -34896 9592 -34769 9608
rect -34896 9528 -34849 9592
rect -34785 9528 -34769 9592
rect -34896 9512 -34769 9528
rect -34896 9388 -34792 9512
rect -34896 9372 -34769 9388
rect -34896 9308 -34849 9372
rect -34785 9308 -34769 9372
rect -34896 9292 -34769 9308
rect -41215 9212 -41088 9228
rect -41215 9148 -41168 9212
rect -41104 9148 -41088 9212
rect -41215 9132 -41088 9148
rect -41215 9068 -41168 9132
rect -41104 9068 -41088 9132
rect -41215 9052 -41088 9068
rect -41215 8988 -41168 9052
rect -41104 8988 -41088 9052
rect -41215 8972 -41088 8988
rect -41215 8908 -41168 8972
rect -41104 8908 -41088 8972
rect -41215 8892 -41088 8908
rect -41215 8828 -41168 8892
rect -41104 8828 -41088 8892
rect -41215 8812 -41088 8828
rect -41215 8748 -41168 8812
rect -41104 8748 -41088 8812
rect -41215 8732 -41088 8748
rect -41215 8668 -41168 8732
rect -41104 8668 -41088 8732
rect -41215 8652 -41088 8668
rect -41215 8588 -41168 8652
rect -41104 8588 -41088 8652
rect -41215 8572 -41088 8588
rect -41215 8508 -41168 8572
rect -41104 8508 -41088 8572
rect -41215 8492 -41088 8508
rect -41215 8428 -41168 8492
rect -41104 8428 -41088 8492
rect -41215 8412 -41088 8428
rect -41215 8348 -41168 8412
rect -41104 8348 -41088 8412
rect -41215 8332 -41088 8348
rect -41215 8268 -41168 8332
rect -41104 8268 -41088 8332
rect -41215 8252 -41088 8268
rect -41215 8188 -41168 8252
rect -41104 8188 -41088 8252
rect -41215 8172 -41088 8188
rect -41215 8108 -41168 8172
rect -41104 8108 -41088 8172
rect -41215 8092 -41088 8108
rect -41215 8028 -41168 8092
rect -41104 8028 -41088 8092
rect -41215 8012 -41088 8028
rect -41215 7948 -41168 8012
rect -41104 7948 -41088 8012
rect -41215 7932 -41088 7948
rect -41215 7868 -41168 7932
rect -41104 7868 -41088 7932
rect -41215 7852 -41088 7868
rect -41215 7788 -41168 7852
rect -41104 7788 -41088 7852
rect -41215 7772 -41088 7788
rect -41215 7708 -41168 7772
rect -41104 7708 -41088 7772
rect -41215 7692 -41088 7708
rect -41215 7628 -41168 7692
rect -41104 7628 -41088 7692
rect -41215 7612 -41088 7628
rect -41215 7548 -41168 7612
rect -41104 7548 -41088 7612
rect -41215 7532 -41088 7548
rect -41215 7468 -41168 7532
rect -41104 7468 -41088 7532
rect -41215 7452 -41088 7468
rect -41215 7388 -41168 7452
rect -41104 7388 -41088 7452
rect -41215 7372 -41088 7388
rect -41215 7308 -41168 7372
rect -41104 7308 -41088 7372
rect -41215 7292 -41088 7308
rect -41215 7228 -41168 7292
rect -41104 7228 -41088 7292
rect -41215 7212 -41088 7228
rect -41215 7148 -41168 7212
rect -41104 7148 -41088 7212
rect -41215 7132 -41088 7148
rect -41215 7068 -41168 7132
rect -41104 7068 -41088 7132
rect -41215 7052 -41088 7068
rect -41215 6988 -41168 7052
rect -41104 6988 -41088 7052
rect -41215 6972 -41088 6988
rect -41215 6908 -41168 6972
rect -41104 6908 -41088 6972
rect -41215 6892 -41088 6908
rect -41215 6828 -41168 6892
rect -41104 6828 -41088 6892
rect -41215 6812 -41088 6828
rect -41215 6748 -41168 6812
rect -41104 6748 -41088 6812
rect -41215 6732 -41088 6748
rect -41215 6668 -41168 6732
rect -41104 6668 -41088 6732
rect -41215 6652 -41088 6668
rect -41215 6588 -41168 6652
rect -41104 6588 -41088 6652
rect -41215 6572 -41088 6588
rect -41215 6508 -41168 6572
rect -41104 6508 -41088 6572
rect -41215 6492 -41088 6508
rect -41215 6428 -41168 6492
rect -41104 6428 -41088 6492
rect -41215 6412 -41088 6428
rect -41215 6348 -41168 6412
rect -41104 6348 -41088 6412
rect -41215 6332 -41088 6348
rect -41215 6268 -41168 6332
rect -41104 6268 -41088 6332
rect -41215 6252 -41088 6268
rect -41215 6188 -41168 6252
rect -41104 6188 -41088 6252
rect -41215 6172 -41088 6188
rect -41215 6108 -41168 6172
rect -41104 6108 -41088 6172
rect -41215 6092 -41088 6108
rect -41215 6028 -41168 6092
rect -41104 6028 -41088 6092
rect -41215 6012 -41088 6028
rect -41215 5948 -41168 6012
rect -41104 5948 -41088 6012
rect -41215 5932 -41088 5948
rect -41215 5868 -41168 5932
rect -41104 5868 -41088 5932
rect -41215 5852 -41088 5868
rect -41215 5788 -41168 5852
rect -41104 5788 -41088 5852
rect -41215 5772 -41088 5788
rect -41215 5708 -41168 5772
rect -41104 5708 -41088 5772
rect -41215 5692 -41088 5708
rect -41215 5628 -41168 5692
rect -41104 5628 -41088 5692
rect -41215 5612 -41088 5628
rect -41215 5548 -41168 5612
rect -41104 5548 -41088 5612
rect -41215 5532 -41088 5548
rect -41215 5468 -41168 5532
rect -41104 5468 -41088 5532
rect -41215 5452 -41088 5468
rect -41215 5388 -41168 5452
rect -41104 5388 -41088 5452
rect -41215 5372 -41088 5388
rect -41215 5308 -41168 5372
rect -41104 5308 -41088 5372
rect -41215 5292 -41088 5308
rect -41215 5228 -41168 5292
rect -41104 5228 -41088 5292
rect -41215 5212 -41088 5228
rect -41215 5148 -41168 5212
rect -41104 5148 -41088 5212
rect -41215 5132 -41088 5148
rect -41215 5068 -41168 5132
rect -41104 5068 -41088 5132
rect -41215 5052 -41088 5068
rect -41215 4988 -41168 5052
rect -41104 4988 -41088 5052
rect -41215 4972 -41088 4988
rect -41215 4908 -41168 4972
rect -41104 4908 -41088 4972
rect -41215 4892 -41088 4908
rect -41215 4828 -41168 4892
rect -41104 4828 -41088 4892
rect -41215 4812 -41088 4828
rect -41215 4748 -41168 4812
rect -41104 4748 -41088 4812
rect -41215 4732 -41088 4748
rect -41215 4668 -41168 4732
rect -41104 4668 -41088 4732
rect -41215 4652 -41088 4668
rect -41215 4588 -41168 4652
rect -41104 4588 -41088 4652
rect -41215 4572 -41088 4588
rect -41215 4508 -41168 4572
rect -41104 4508 -41088 4572
rect -41215 4492 -41088 4508
rect -41215 4428 -41168 4492
rect -41104 4428 -41088 4492
rect -41215 4412 -41088 4428
rect -41215 4348 -41168 4412
rect -41104 4348 -41088 4412
rect -41215 4332 -41088 4348
rect -41215 4268 -41168 4332
rect -41104 4268 -41088 4332
rect -41215 4252 -41088 4268
rect -41215 4188 -41168 4252
rect -41104 4188 -41088 4252
rect -41215 4172 -41088 4188
rect -41215 4108 -41168 4172
rect -41104 4108 -41088 4172
rect -41215 4092 -41088 4108
rect -41215 4028 -41168 4092
rect -41104 4028 -41088 4092
rect -41215 4012 -41088 4028
rect -41215 3948 -41168 4012
rect -41104 3948 -41088 4012
rect -41215 3932 -41088 3948
rect -41215 3868 -41168 3932
rect -41104 3868 -41088 3932
rect -41215 3852 -41088 3868
rect -41215 3788 -41168 3852
rect -41104 3788 -41088 3852
rect -41215 3772 -41088 3788
rect -41215 3708 -41168 3772
rect -41104 3708 -41088 3772
rect -41215 3692 -41088 3708
rect -41215 3628 -41168 3692
rect -41104 3628 -41088 3692
rect -41215 3612 -41088 3628
rect -41215 3548 -41168 3612
rect -41104 3548 -41088 3612
rect -41215 3532 -41088 3548
rect -41215 3468 -41168 3532
rect -41104 3468 -41088 3532
rect -41215 3452 -41088 3468
rect -41215 3388 -41168 3452
rect -41104 3388 -41088 3452
rect -41215 3372 -41088 3388
rect -44335 2961 -44231 3339
rect -41215 3308 -41168 3372
rect -41104 3308 -41088 3372
rect -40925 9252 -35003 9261
rect -40925 3348 -40916 9252
rect -35012 3348 -35003 9252
rect -40925 3339 -35003 3348
rect -34896 9228 -34849 9292
rect -34785 9228 -34769 9292
rect -31697 9261 -31593 9639
rect -28577 9608 -28530 9672
rect -28466 9608 -28450 9672
rect -28287 15552 -22365 15561
rect -28287 9648 -28278 15552
rect -22374 9648 -22365 15552
rect -28287 9639 -22365 9648
rect -22258 15528 -22211 15592
rect -22147 15528 -22131 15592
rect -19059 15561 -18955 15939
rect -15939 15908 -15892 15972
rect -15828 15908 -15812 15972
rect -15649 21852 -9727 21861
rect -15649 15948 -15640 21852
rect -9736 15948 -9727 21852
rect -15649 15939 -9727 15948
rect -9620 21828 -9573 21892
rect -9509 21828 -9493 21892
rect -6421 21861 -6317 22239
rect -3301 22208 -3254 22272
rect -3190 22208 -3174 22272
rect -3011 28152 2911 28161
rect -3011 22248 -3002 28152
rect 2902 22248 2911 28152
rect -3011 22239 2911 22248
rect 3018 28128 3065 28192
rect 3129 28128 3145 28192
rect 6217 28161 6321 28539
rect 9337 28508 9384 28572
rect 9448 28508 9464 28572
rect 9627 34452 15549 34461
rect 9627 28548 9636 34452
rect 15540 28548 15549 34452
rect 9627 28539 15549 28548
rect 15656 34428 15703 34492
rect 15767 34428 15783 34492
rect 18855 34461 18959 34839
rect 21975 34808 22022 34872
rect 22086 34808 22102 34872
rect 22265 40752 28187 40761
rect 22265 34848 22274 40752
rect 28178 34848 28187 40752
rect 22265 34839 28187 34848
rect 28294 40728 28341 40792
rect 28405 40728 28421 40792
rect 31493 40761 31597 41139
rect 34613 41108 34660 41172
rect 34724 41108 34740 41172
rect 34903 47052 40825 47061
rect 34903 41148 34912 47052
rect 40816 41148 40825 47052
rect 34903 41139 40825 41148
rect 40932 47028 40979 47092
rect 41043 47028 41059 47092
rect 44131 47061 44235 47250
rect 47251 47188 47355 47250
rect 47251 47172 47378 47188
rect 47251 47108 47298 47172
rect 47362 47108 47378 47172
rect 47251 47092 47378 47108
rect 40932 47012 41059 47028
rect 40932 46948 40979 47012
rect 41043 46948 41059 47012
rect 40932 46932 41059 46948
rect 40932 46868 40979 46932
rect 41043 46868 41059 46932
rect 40932 46852 41059 46868
rect 40932 46788 40979 46852
rect 41043 46788 41059 46852
rect 40932 46772 41059 46788
rect 40932 46708 40979 46772
rect 41043 46708 41059 46772
rect 40932 46692 41059 46708
rect 40932 46628 40979 46692
rect 41043 46628 41059 46692
rect 40932 46612 41059 46628
rect 40932 46548 40979 46612
rect 41043 46548 41059 46612
rect 40932 46532 41059 46548
rect 40932 46468 40979 46532
rect 41043 46468 41059 46532
rect 40932 46452 41059 46468
rect 40932 46388 40979 46452
rect 41043 46388 41059 46452
rect 40932 46372 41059 46388
rect 40932 46308 40979 46372
rect 41043 46308 41059 46372
rect 40932 46292 41059 46308
rect 40932 46228 40979 46292
rect 41043 46228 41059 46292
rect 40932 46212 41059 46228
rect 40932 46148 40979 46212
rect 41043 46148 41059 46212
rect 40932 46132 41059 46148
rect 40932 46068 40979 46132
rect 41043 46068 41059 46132
rect 40932 46052 41059 46068
rect 40932 45988 40979 46052
rect 41043 45988 41059 46052
rect 40932 45972 41059 45988
rect 40932 45908 40979 45972
rect 41043 45908 41059 45972
rect 40932 45892 41059 45908
rect 40932 45828 40979 45892
rect 41043 45828 41059 45892
rect 40932 45812 41059 45828
rect 40932 45748 40979 45812
rect 41043 45748 41059 45812
rect 40932 45732 41059 45748
rect 40932 45668 40979 45732
rect 41043 45668 41059 45732
rect 40932 45652 41059 45668
rect 40932 45588 40979 45652
rect 41043 45588 41059 45652
rect 40932 45572 41059 45588
rect 40932 45508 40979 45572
rect 41043 45508 41059 45572
rect 40932 45492 41059 45508
rect 40932 45428 40979 45492
rect 41043 45428 41059 45492
rect 40932 45412 41059 45428
rect 40932 45348 40979 45412
rect 41043 45348 41059 45412
rect 40932 45332 41059 45348
rect 40932 45268 40979 45332
rect 41043 45268 41059 45332
rect 40932 45252 41059 45268
rect 40932 45188 40979 45252
rect 41043 45188 41059 45252
rect 40932 45172 41059 45188
rect 40932 45108 40979 45172
rect 41043 45108 41059 45172
rect 40932 45092 41059 45108
rect 40932 45028 40979 45092
rect 41043 45028 41059 45092
rect 40932 45012 41059 45028
rect 40932 44948 40979 45012
rect 41043 44948 41059 45012
rect 40932 44932 41059 44948
rect 40932 44868 40979 44932
rect 41043 44868 41059 44932
rect 40932 44852 41059 44868
rect 40932 44788 40979 44852
rect 41043 44788 41059 44852
rect 40932 44772 41059 44788
rect 40932 44708 40979 44772
rect 41043 44708 41059 44772
rect 40932 44692 41059 44708
rect 40932 44628 40979 44692
rect 41043 44628 41059 44692
rect 40932 44612 41059 44628
rect 40932 44548 40979 44612
rect 41043 44548 41059 44612
rect 40932 44532 41059 44548
rect 40932 44468 40979 44532
rect 41043 44468 41059 44532
rect 40932 44452 41059 44468
rect 40932 44388 40979 44452
rect 41043 44388 41059 44452
rect 40932 44372 41059 44388
rect 40932 44308 40979 44372
rect 41043 44308 41059 44372
rect 40932 44292 41059 44308
rect 40932 44228 40979 44292
rect 41043 44228 41059 44292
rect 40932 44212 41059 44228
rect 40932 44148 40979 44212
rect 41043 44148 41059 44212
rect 40932 44132 41059 44148
rect 40932 44068 40979 44132
rect 41043 44068 41059 44132
rect 40932 44052 41059 44068
rect 40932 43988 40979 44052
rect 41043 43988 41059 44052
rect 40932 43972 41059 43988
rect 40932 43908 40979 43972
rect 41043 43908 41059 43972
rect 40932 43892 41059 43908
rect 40932 43828 40979 43892
rect 41043 43828 41059 43892
rect 40932 43812 41059 43828
rect 40932 43748 40979 43812
rect 41043 43748 41059 43812
rect 40932 43732 41059 43748
rect 40932 43668 40979 43732
rect 41043 43668 41059 43732
rect 40932 43652 41059 43668
rect 40932 43588 40979 43652
rect 41043 43588 41059 43652
rect 40932 43572 41059 43588
rect 40932 43508 40979 43572
rect 41043 43508 41059 43572
rect 40932 43492 41059 43508
rect 40932 43428 40979 43492
rect 41043 43428 41059 43492
rect 40932 43412 41059 43428
rect 40932 43348 40979 43412
rect 41043 43348 41059 43412
rect 40932 43332 41059 43348
rect 40932 43268 40979 43332
rect 41043 43268 41059 43332
rect 40932 43252 41059 43268
rect 40932 43188 40979 43252
rect 41043 43188 41059 43252
rect 40932 43172 41059 43188
rect 40932 43108 40979 43172
rect 41043 43108 41059 43172
rect 40932 43092 41059 43108
rect 40932 43028 40979 43092
rect 41043 43028 41059 43092
rect 40932 43012 41059 43028
rect 40932 42948 40979 43012
rect 41043 42948 41059 43012
rect 40932 42932 41059 42948
rect 40932 42868 40979 42932
rect 41043 42868 41059 42932
rect 40932 42852 41059 42868
rect 40932 42788 40979 42852
rect 41043 42788 41059 42852
rect 40932 42772 41059 42788
rect 40932 42708 40979 42772
rect 41043 42708 41059 42772
rect 40932 42692 41059 42708
rect 40932 42628 40979 42692
rect 41043 42628 41059 42692
rect 40932 42612 41059 42628
rect 40932 42548 40979 42612
rect 41043 42548 41059 42612
rect 40932 42532 41059 42548
rect 40932 42468 40979 42532
rect 41043 42468 41059 42532
rect 40932 42452 41059 42468
rect 40932 42388 40979 42452
rect 41043 42388 41059 42452
rect 40932 42372 41059 42388
rect 40932 42308 40979 42372
rect 41043 42308 41059 42372
rect 40932 42292 41059 42308
rect 40932 42228 40979 42292
rect 41043 42228 41059 42292
rect 40932 42212 41059 42228
rect 40932 42148 40979 42212
rect 41043 42148 41059 42212
rect 40932 42132 41059 42148
rect 40932 42068 40979 42132
rect 41043 42068 41059 42132
rect 40932 42052 41059 42068
rect 40932 41988 40979 42052
rect 41043 41988 41059 42052
rect 40932 41972 41059 41988
rect 40932 41908 40979 41972
rect 41043 41908 41059 41972
rect 40932 41892 41059 41908
rect 40932 41828 40979 41892
rect 41043 41828 41059 41892
rect 40932 41812 41059 41828
rect 40932 41748 40979 41812
rect 41043 41748 41059 41812
rect 40932 41732 41059 41748
rect 40932 41668 40979 41732
rect 41043 41668 41059 41732
rect 40932 41652 41059 41668
rect 40932 41588 40979 41652
rect 41043 41588 41059 41652
rect 40932 41572 41059 41588
rect 40932 41508 40979 41572
rect 41043 41508 41059 41572
rect 40932 41492 41059 41508
rect 40932 41428 40979 41492
rect 41043 41428 41059 41492
rect 40932 41412 41059 41428
rect 40932 41348 40979 41412
rect 41043 41348 41059 41412
rect 40932 41332 41059 41348
rect 40932 41268 40979 41332
rect 41043 41268 41059 41332
rect 40932 41252 41059 41268
rect 40932 41188 40979 41252
rect 41043 41188 41059 41252
rect 40932 41172 41059 41188
rect 34613 41092 34740 41108
rect 34613 41028 34660 41092
rect 34724 41028 34740 41092
rect 34613 41012 34740 41028
rect 34613 40888 34717 41012
rect 34613 40872 34740 40888
rect 34613 40808 34660 40872
rect 34724 40808 34740 40872
rect 34613 40792 34740 40808
rect 28294 40712 28421 40728
rect 28294 40648 28341 40712
rect 28405 40648 28421 40712
rect 28294 40632 28421 40648
rect 28294 40568 28341 40632
rect 28405 40568 28421 40632
rect 28294 40552 28421 40568
rect 28294 40488 28341 40552
rect 28405 40488 28421 40552
rect 28294 40472 28421 40488
rect 28294 40408 28341 40472
rect 28405 40408 28421 40472
rect 28294 40392 28421 40408
rect 28294 40328 28341 40392
rect 28405 40328 28421 40392
rect 28294 40312 28421 40328
rect 28294 40248 28341 40312
rect 28405 40248 28421 40312
rect 28294 40232 28421 40248
rect 28294 40168 28341 40232
rect 28405 40168 28421 40232
rect 28294 40152 28421 40168
rect 28294 40088 28341 40152
rect 28405 40088 28421 40152
rect 28294 40072 28421 40088
rect 28294 40008 28341 40072
rect 28405 40008 28421 40072
rect 28294 39992 28421 40008
rect 28294 39928 28341 39992
rect 28405 39928 28421 39992
rect 28294 39912 28421 39928
rect 28294 39848 28341 39912
rect 28405 39848 28421 39912
rect 28294 39832 28421 39848
rect 28294 39768 28341 39832
rect 28405 39768 28421 39832
rect 28294 39752 28421 39768
rect 28294 39688 28341 39752
rect 28405 39688 28421 39752
rect 28294 39672 28421 39688
rect 28294 39608 28341 39672
rect 28405 39608 28421 39672
rect 28294 39592 28421 39608
rect 28294 39528 28341 39592
rect 28405 39528 28421 39592
rect 28294 39512 28421 39528
rect 28294 39448 28341 39512
rect 28405 39448 28421 39512
rect 28294 39432 28421 39448
rect 28294 39368 28341 39432
rect 28405 39368 28421 39432
rect 28294 39352 28421 39368
rect 28294 39288 28341 39352
rect 28405 39288 28421 39352
rect 28294 39272 28421 39288
rect 28294 39208 28341 39272
rect 28405 39208 28421 39272
rect 28294 39192 28421 39208
rect 28294 39128 28341 39192
rect 28405 39128 28421 39192
rect 28294 39112 28421 39128
rect 28294 39048 28341 39112
rect 28405 39048 28421 39112
rect 28294 39032 28421 39048
rect 28294 38968 28341 39032
rect 28405 38968 28421 39032
rect 28294 38952 28421 38968
rect 28294 38888 28341 38952
rect 28405 38888 28421 38952
rect 28294 38872 28421 38888
rect 28294 38808 28341 38872
rect 28405 38808 28421 38872
rect 28294 38792 28421 38808
rect 28294 38728 28341 38792
rect 28405 38728 28421 38792
rect 28294 38712 28421 38728
rect 28294 38648 28341 38712
rect 28405 38648 28421 38712
rect 28294 38632 28421 38648
rect 28294 38568 28341 38632
rect 28405 38568 28421 38632
rect 28294 38552 28421 38568
rect 28294 38488 28341 38552
rect 28405 38488 28421 38552
rect 28294 38472 28421 38488
rect 28294 38408 28341 38472
rect 28405 38408 28421 38472
rect 28294 38392 28421 38408
rect 28294 38328 28341 38392
rect 28405 38328 28421 38392
rect 28294 38312 28421 38328
rect 28294 38248 28341 38312
rect 28405 38248 28421 38312
rect 28294 38232 28421 38248
rect 28294 38168 28341 38232
rect 28405 38168 28421 38232
rect 28294 38152 28421 38168
rect 28294 38088 28341 38152
rect 28405 38088 28421 38152
rect 28294 38072 28421 38088
rect 28294 38008 28341 38072
rect 28405 38008 28421 38072
rect 28294 37992 28421 38008
rect 28294 37928 28341 37992
rect 28405 37928 28421 37992
rect 28294 37912 28421 37928
rect 28294 37848 28341 37912
rect 28405 37848 28421 37912
rect 28294 37832 28421 37848
rect 28294 37768 28341 37832
rect 28405 37768 28421 37832
rect 28294 37752 28421 37768
rect 28294 37688 28341 37752
rect 28405 37688 28421 37752
rect 28294 37672 28421 37688
rect 28294 37608 28341 37672
rect 28405 37608 28421 37672
rect 28294 37592 28421 37608
rect 28294 37528 28341 37592
rect 28405 37528 28421 37592
rect 28294 37512 28421 37528
rect 28294 37448 28341 37512
rect 28405 37448 28421 37512
rect 28294 37432 28421 37448
rect 28294 37368 28341 37432
rect 28405 37368 28421 37432
rect 28294 37352 28421 37368
rect 28294 37288 28341 37352
rect 28405 37288 28421 37352
rect 28294 37272 28421 37288
rect 28294 37208 28341 37272
rect 28405 37208 28421 37272
rect 28294 37192 28421 37208
rect 28294 37128 28341 37192
rect 28405 37128 28421 37192
rect 28294 37112 28421 37128
rect 28294 37048 28341 37112
rect 28405 37048 28421 37112
rect 28294 37032 28421 37048
rect 28294 36968 28341 37032
rect 28405 36968 28421 37032
rect 28294 36952 28421 36968
rect 28294 36888 28341 36952
rect 28405 36888 28421 36952
rect 28294 36872 28421 36888
rect 28294 36808 28341 36872
rect 28405 36808 28421 36872
rect 28294 36792 28421 36808
rect 28294 36728 28341 36792
rect 28405 36728 28421 36792
rect 28294 36712 28421 36728
rect 28294 36648 28341 36712
rect 28405 36648 28421 36712
rect 28294 36632 28421 36648
rect 28294 36568 28341 36632
rect 28405 36568 28421 36632
rect 28294 36552 28421 36568
rect 28294 36488 28341 36552
rect 28405 36488 28421 36552
rect 28294 36472 28421 36488
rect 28294 36408 28341 36472
rect 28405 36408 28421 36472
rect 28294 36392 28421 36408
rect 28294 36328 28341 36392
rect 28405 36328 28421 36392
rect 28294 36312 28421 36328
rect 28294 36248 28341 36312
rect 28405 36248 28421 36312
rect 28294 36232 28421 36248
rect 28294 36168 28341 36232
rect 28405 36168 28421 36232
rect 28294 36152 28421 36168
rect 28294 36088 28341 36152
rect 28405 36088 28421 36152
rect 28294 36072 28421 36088
rect 28294 36008 28341 36072
rect 28405 36008 28421 36072
rect 28294 35992 28421 36008
rect 28294 35928 28341 35992
rect 28405 35928 28421 35992
rect 28294 35912 28421 35928
rect 28294 35848 28341 35912
rect 28405 35848 28421 35912
rect 28294 35832 28421 35848
rect 28294 35768 28341 35832
rect 28405 35768 28421 35832
rect 28294 35752 28421 35768
rect 28294 35688 28341 35752
rect 28405 35688 28421 35752
rect 28294 35672 28421 35688
rect 28294 35608 28341 35672
rect 28405 35608 28421 35672
rect 28294 35592 28421 35608
rect 28294 35528 28341 35592
rect 28405 35528 28421 35592
rect 28294 35512 28421 35528
rect 28294 35448 28341 35512
rect 28405 35448 28421 35512
rect 28294 35432 28421 35448
rect 28294 35368 28341 35432
rect 28405 35368 28421 35432
rect 28294 35352 28421 35368
rect 28294 35288 28341 35352
rect 28405 35288 28421 35352
rect 28294 35272 28421 35288
rect 28294 35208 28341 35272
rect 28405 35208 28421 35272
rect 28294 35192 28421 35208
rect 28294 35128 28341 35192
rect 28405 35128 28421 35192
rect 28294 35112 28421 35128
rect 28294 35048 28341 35112
rect 28405 35048 28421 35112
rect 28294 35032 28421 35048
rect 28294 34968 28341 35032
rect 28405 34968 28421 35032
rect 28294 34952 28421 34968
rect 28294 34888 28341 34952
rect 28405 34888 28421 34952
rect 28294 34872 28421 34888
rect 21975 34792 22102 34808
rect 21975 34728 22022 34792
rect 22086 34728 22102 34792
rect 21975 34712 22102 34728
rect 21975 34588 22079 34712
rect 21975 34572 22102 34588
rect 21975 34508 22022 34572
rect 22086 34508 22102 34572
rect 21975 34492 22102 34508
rect 15656 34412 15783 34428
rect 15656 34348 15703 34412
rect 15767 34348 15783 34412
rect 15656 34332 15783 34348
rect 15656 34268 15703 34332
rect 15767 34268 15783 34332
rect 15656 34252 15783 34268
rect 15656 34188 15703 34252
rect 15767 34188 15783 34252
rect 15656 34172 15783 34188
rect 15656 34108 15703 34172
rect 15767 34108 15783 34172
rect 15656 34092 15783 34108
rect 15656 34028 15703 34092
rect 15767 34028 15783 34092
rect 15656 34012 15783 34028
rect 15656 33948 15703 34012
rect 15767 33948 15783 34012
rect 15656 33932 15783 33948
rect 15656 33868 15703 33932
rect 15767 33868 15783 33932
rect 15656 33852 15783 33868
rect 15656 33788 15703 33852
rect 15767 33788 15783 33852
rect 15656 33772 15783 33788
rect 15656 33708 15703 33772
rect 15767 33708 15783 33772
rect 15656 33692 15783 33708
rect 15656 33628 15703 33692
rect 15767 33628 15783 33692
rect 15656 33612 15783 33628
rect 15656 33548 15703 33612
rect 15767 33548 15783 33612
rect 15656 33532 15783 33548
rect 15656 33468 15703 33532
rect 15767 33468 15783 33532
rect 15656 33452 15783 33468
rect 15656 33388 15703 33452
rect 15767 33388 15783 33452
rect 15656 33372 15783 33388
rect 15656 33308 15703 33372
rect 15767 33308 15783 33372
rect 15656 33292 15783 33308
rect 15656 33228 15703 33292
rect 15767 33228 15783 33292
rect 15656 33212 15783 33228
rect 15656 33148 15703 33212
rect 15767 33148 15783 33212
rect 15656 33132 15783 33148
rect 15656 33068 15703 33132
rect 15767 33068 15783 33132
rect 15656 33052 15783 33068
rect 15656 32988 15703 33052
rect 15767 32988 15783 33052
rect 15656 32972 15783 32988
rect 15656 32908 15703 32972
rect 15767 32908 15783 32972
rect 15656 32892 15783 32908
rect 15656 32828 15703 32892
rect 15767 32828 15783 32892
rect 15656 32812 15783 32828
rect 15656 32748 15703 32812
rect 15767 32748 15783 32812
rect 15656 32732 15783 32748
rect 15656 32668 15703 32732
rect 15767 32668 15783 32732
rect 15656 32652 15783 32668
rect 15656 32588 15703 32652
rect 15767 32588 15783 32652
rect 15656 32572 15783 32588
rect 15656 32508 15703 32572
rect 15767 32508 15783 32572
rect 15656 32492 15783 32508
rect 15656 32428 15703 32492
rect 15767 32428 15783 32492
rect 15656 32412 15783 32428
rect 15656 32348 15703 32412
rect 15767 32348 15783 32412
rect 15656 32332 15783 32348
rect 15656 32268 15703 32332
rect 15767 32268 15783 32332
rect 15656 32252 15783 32268
rect 15656 32188 15703 32252
rect 15767 32188 15783 32252
rect 15656 32172 15783 32188
rect 15656 32108 15703 32172
rect 15767 32108 15783 32172
rect 15656 32092 15783 32108
rect 15656 32028 15703 32092
rect 15767 32028 15783 32092
rect 15656 32012 15783 32028
rect 15656 31948 15703 32012
rect 15767 31948 15783 32012
rect 15656 31932 15783 31948
rect 15656 31868 15703 31932
rect 15767 31868 15783 31932
rect 15656 31852 15783 31868
rect 15656 31788 15703 31852
rect 15767 31788 15783 31852
rect 15656 31772 15783 31788
rect 15656 31708 15703 31772
rect 15767 31708 15783 31772
rect 15656 31692 15783 31708
rect 15656 31628 15703 31692
rect 15767 31628 15783 31692
rect 15656 31612 15783 31628
rect 15656 31548 15703 31612
rect 15767 31548 15783 31612
rect 15656 31532 15783 31548
rect 15656 31468 15703 31532
rect 15767 31468 15783 31532
rect 15656 31452 15783 31468
rect 15656 31388 15703 31452
rect 15767 31388 15783 31452
rect 15656 31372 15783 31388
rect 15656 31308 15703 31372
rect 15767 31308 15783 31372
rect 15656 31292 15783 31308
rect 15656 31228 15703 31292
rect 15767 31228 15783 31292
rect 15656 31212 15783 31228
rect 15656 31148 15703 31212
rect 15767 31148 15783 31212
rect 15656 31132 15783 31148
rect 15656 31068 15703 31132
rect 15767 31068 15783 31132
rect 15656 31052 15783 31068
rect 15656 30988 15703 31052
rect 15767 30988 15783 31052
rect 15656 30972 15783 30988
rect 15656 30908 15703 30972
rect 15767 30908 15783 30972
rect 15656 30892 15783 30908
rect 15656 30828 15703 30892
rect 15767 30828 15783 30892
rect 15656 30812 15783 30828
rect 15656 30748 15703 30812
rect 15767 30748 15783 30812
rect 15656 30732 15783 30748
rect 15656 30668 15703 30732
rect 15767 30668 15783 30732
rect 15656 30652 15783 30668
rect 15656 30588 15703 30652
rect 15767 30588 15783 30652
rect 15656 30572 15783 30588
rect 15656 30508 15703 30572
rect 15767 30508 15783 30572
rect 15656 30492 15783 30508
rect 15656 30428 15703 30492
rect 15767 30428 15783 30492
rect 15656 30412 15783 30428
rect 15656 30348 15703 30412
rect 15767 30348 15783 30412
rect 15656 30332 15783 30348
rect 15656 30268 15703 30332
rect 15767 30268 15783 30332
rect 15656 30252 15783 30268
rect 15656 30188 15703 30252
rect 15767 30188 15783 30252
rect 15656 30172 15783 30188
rect 15656 30108 15703 30172
rect 15767 30108 15783 30172
rect 15656 30092 15783 30108
rect 15656 30028 15703 30092
rect 15767 30028 15783 30092
rect 15656 30012 15783 30028
rect 15656 29948 15703 30012
rect 15767 29948 15783 30012
rect 15656 29932 15783 29948
rect 15656 29868 15703 29932
rect 15767 29868 15783 29932
rect 15656 29852 15783 29868
rect 15656 29788 15703 29852
rect 15767 29788 15783 29852
rect 15656 29772 15783 29788
rect 15656 29708 15703 29772
rect 15767 29708 15783 29772
rect 15656 29692 15783 29708
rect 15656 29628 15703 29692
rect 15767 29628 15783 29692
rect 15656 29612 15783 29628
rect 15656 29548 15703 29612
rect 15767 29548 15783 29612
rect 15656 29532 15783 29548
rect 15656 29468 15703 29532
rect 15767 29468 15783 29532
rect 15656 29452 15783 29468
rect 15656 29388 15703 29452
rect 15767 29388 15783 29452
rect 15656 29372 15783 29388
rect 15656 29308 15703 29372
rect 15767 29308 15783 29372
rect 15656 29292 15783 29308
rect 15656 29228 15703 29292
rect 15767 29228 15783 29292
rect 15656 29212 15783 29228
rect 15656 29148 15703 29212
rect 15767 29148 15783 29212
rect 15656 29132 15783 29148
rect 15656 29068 15703 29132
rect 15767 29068 15783 29132
rect 15656 29052 15783 29068
rect 15656 28988 15703 29052
rect 15767 28988 15783 29052
rect 15656 28972 15783 28988
rect 15656 28908 15703 28972
rect 15767 28908 15783 28972
rect 15656 28892 15783 28908
rect 15656 28828 15703 28892
rect 15767 28828 15783 28892
rect 15656 28812 15783 28828
rect 15656 28748 15703 28812
rect 15767 28748 15783 28812
rect 15656 28732 15783 28748
rect 15656 28668 15703 28732
rect 15767 28668 15783 28732
rect 15656 28652 15783 28668
rect 15656 28588 15703 28652
rect 15767 28588 15783 28652
rect 15656 28572 15783 28588
rect 9337 28492 9464 28508
rect 9337 28428 9384 28492
rect 9448 28428 9464 28492
rect 9337 28412 9464 28428
rect 9337 28288 9441 28412
rect 9337 28272 9464 28288
rect 9337 28208 9384 28272
rect 9448 28208 9464 28272
rect 9337 28192 9464 28208
rect 3018 28112 3145 28128
rect 3018 28048 3065 28112
rect 3129 28048 3145 28112
rect 3018 28032 3145 28048
rect 3018 27968 3065 28032
rect 3129 27968 3145 28032
rect 3018 27952 3145 27968
rect 3018 27888 3065 27952
rect 3129 27888 3145 27952
rect 3018 27872 3145 27888
rect 3018 27808 3065 27872
rect 3129 27808 3145 27872
rect 3018 27792 3145 27808
rect 3018 27728 3065 27792
rect 3129 27728 3145 27792
rect 3018 27712 3145 27728
rect 3018 27648 3065 27712
rect 3129 27648 3145 27712
rect 3018 27632 3145 27648
rect 3018 27568 3065 27632
rect 3129 27568 3145 27632
rect 3018 27552 3145 27568
rect 3018 27488 3065 27552
rect 3129 27488 3145 27552
rect 3018 27472 3145 27488
rect 3018 27408 3065 27472
rect 3129 27408 3145 27472
rect 3018 27392 3145 27408
rect 3018 27328 3065 27392
rect 3129 27328 3145 27392
rect 3018 27312 3145 27328
rect 3018 27248 3065 27312
rect 3129 27248 3145 27312
rect 3018 27232 3145 27248
rect 3018 27168 3065 27232
rect 3129 27168 3145 27232
rect 3018 27152 3145 27168
rect 3018 27088 3065 27152
rect 3129 27088 3145 27152
rect 3018 27072 3145 27088
rect 3018 27008 3065 27072
rect 3129 27008 3145 27072
rect 3018 26992 3145 27008
rect 3018 26928 3065 26992
rect 3129 26928 3145 26992
rect 3018 26912 3145 26928
rect 3018 26848 3065 26912
rect 3129 26848 3145 26912
rect 3018 26832 3145 26848
rect 3018 26768 3065 26832
rect 3129 26768 3145 26832
rect 3018 26752 3145 26768
rect 3018 26688 3065 26752
rect 3129 26688 3145 26752
rect 3018 26672 3145 26688
rect 3018 26608 3065 26672
rect 3129 26608 3145 26672
rect 3018 26592 3145 26608
rect 3018 26528 3065 26592
rect 3129 26528 3145 26592
rect 3018 26512 3145 26528
rect 3018 26448 3065 26512
rect 3129 26448 3145 26512
rect 3018 26432 3145 26448
rect 3018 26368 3065 26432
rect 3129 26368 3145 26432
rect 3018 26352 3145 26368
rect 3018 26288 3065 26352
rect 3129 26288 3145 26352
rect 3018 26272 3145 26288
rect 3018 26208 3065 26272
rect 3129 26208 3145 26272
rect 3018 26192 3145 26208
rect 3018 26128 3065 26192
rect 3129 26128 3145 26192
rect 3018 26112 3145 26128
rect 3018 26048 3065 26112
rect 3129 26048 3145 26112
rect 3018 26032 3145 26048
rect 3018 25968 3065 26032
rect 3129 25968 3145 26032
rect 3018 25952 3145 25968
rect 3018 25888 3065 25952
rect 3129 25888 3145 25952
rect 3018 25872 3145 25888
rect 3018 25808 3065 25872
rect 3129 25808 3145 25872
rect 3018 25792 3145 25808
rect 3018 25728 3065 25792
rect 3129 25728 3145 25792
rect 3018 25712 3145 25728
rect 3018 25648 3065 25712
rect 3129 25648 3145 25712
rect 3018 25632 3145 25648
rect 3018 25568 3065 25632
rect 3129 25568 3145 25632
rect 3018 25552 3145 25568
rect 3018 25488 3065 25552
rect 3129 25488 3145 25552
rect 3018 25472 3145 25488
rect 3018 25408 3065 25472
rect 3129 25408 3145 25472
rect 3018 25392 3145 25408
rect 3018 25328 3065 25392
rect 3129 25328 3145 25392
rect 3018 25312 3145 25328
rect 3018 25248 3065 25312
rect 3129 25248 3145 25312
rect 3018 25232 3145 25248
rect 3018 25168 3065 25232
rect 3129 25168 3145 25232
rect 3018 25152 3145 25168
rect 3018 25088 3065 25152
rect 3129 25088 3145 25152
rect 3018 25072 3145 25088
rect 3018 25008 3065 25072
rect 3129 25008 3145 25072
rect 3018 24992 3145 25008
rect 3018 24928 3065 24992
rect 3129 24928 3145 24992
rect 3018 24912 3145 24928
rect 3018 24848 3065 24912
rect 3129 24848 3145 24912
rect 3018 24832 3145 24848
rect 3018 24768 3065 24832
rect 3129 24768 3145 24832
rect 3018 24752 3145 24768
rect 3018 24688 3065 24752
rect 3129 24688 3145 24752
rect 3018 24672 3145 24688
rect 3018 24608 3065 24672
rect 3129 24608 3145 24672
rect 3018 24592 3145 24608
rect 3018 24528 3065 24592
rect 3129 24528 3145 24592
rect 3018 24512 3145 24528
rect 3018 24448 3065 24512
rect 3129 24448 3145 24512
rect 3018 24432 3145 24448
rect 3018 24368 3065 24432
rect 3129 24368 3145 24432
rect 3018 24352 3145 24368
rect 3018 24288 3065 24352
rect 3129 24288 3145 24352
rect 3018 24272 3145 24288
rect 3018 24208 3065 24272
rect 3129 24208 3145 24272
rect 3018 24192 3145 24208
rect 3018 24128 3065 24192
rect 3129 24128 3145 24192
rect 3018 24112 3145 24128
rect 3018 24048 3065 24112
rect 3129 24048 3145 24112
rect 3018 24032 3145 24048
rect 3018 23968 3065 24032
rect 3129 23968 3145 24032
rect 3018 23952 3145 23968
rect 3018 23888 3065 23952
rect 3129 23888 3145 23952
rect 3018 23872 3145 23888
rect 3018 23808 3065 23872
rect 3129 23808 3145 23872
rect 3018 23792 3145 23808
rect 3018 23728 3065 23792
rect 3129 23728 3145 23792
rect 3018 23712 3145 23728
rect 3018 23648 3065 23712
rect 3129 23648 3145 23712
rect 3018 23632 3145 23648
rect 3018 23568 3065 23632
rect 3129 23568 3145 23632
rect 3018 23552 3145 23568
rect 3018 23488 3065 23552
rect 3129 23488 3145 23552
rect 3018 23472 3145 23488
rect 3018 23408 3065 23472
rect 3129 23408 3145 23472
rect 3018 23392 3145 23408
rect 3018 23328 3065 23392
rect 3129 23328 3145 23392
rect 3018 23312 3145 23328
rect 3018 23248 3065 23312
rect 3129 23248 3145 23312
rect 3018 23232 3145 23248
rect 3018 23168 3065 23232
rect 3129 23168 3145 23232
rect 3018 23152 3145 23168
rect 3018 23088 3065 23152
rect 3129 23088 3145 23152
rect 3018 23072 3145 23088
rect 3018 23008 3065 23072
rect 3129 23008 3145 23072
rect 3018 22992 3145 23008
rect 3018 22928 3065 22992
rect 3129 22928 3145 22992
rect 3018 22912 3145 22928
rect 3018 22848 3065 22912
rect 3129 22848 3145 22912
rect 3018 22832 3145 22848
rect 3018 22768 3065 22832
rect 3129 22768 3145 22832
rect 3018 22752 3145 22768
rect 3018 22688 3065 22752
rect 3129 22688 3145 22752
rect 3018 22672 3145 22688
rect 3018 22608 3065 22672
rect 3129 22608 3145 22672
rect 3018 22592 3145 22608
rect 3018 22528 3065 22592
rect 3129 22528 3145 22592
rect 3018 22512 3145 22528
rect 3018 22448 3065 22512
rect 3129 22448 3145 22512
rect 3018 22432 3145 22448
rect 3018 22368 3065 22432
rect 3129 22368 3145 22432
rect 3018 22352 3145 22368
rect 3018 22288 3065 22352
rect 3129 22288 3145 22352
rect 3018 22272 3145 22288
rect -3301 22192 -3174 22208
rect -3301 22128 -3254 22192
rect -3190 22128 -3174 22192
rect -3301 22112 -3174 22128
rect -3301 21988 -3197 22112
rect -3301 21972 -3174 21988
rect -3301 21908 -3254 21972
rect -3190 21908 -3174 21972
rect -3301 21892 -3174 21908
rect -9620 21812 -9493 21828
rect -9620 21748 -9573 21812
rect -9509 21748 -9493 21812
rect -9620 21732 -9493 21748
rect -9620 21668 -9573 21732
rect -9509 21668 -9493 21732
rect -9620 21652 -9493 21668
rect -9620 21588 -9573 21652
rect -9509 21588 -9493 21652
rect -9620 21572 -9493 21588
rect -9620 21508 -9573 21572
rect -9509 21508 -9493 21572
rect -9620 21492 -9493 21508
rect -9620 21428 -9573 21492
rect -9509 21428 -9493 21492
rect -9620 21412 -9493 21428
rect -9620 21348 -9573 21412
rect -9509 21348 -9493 21412
rect -9620 21332 -9493 21348
rect -9620 21268 -9573 21332
rect -9509 21268 -9493 21332
rect -9620 21252 -9493 21268
rect -9620 21188 -9573 21252
rect -9509 21188 -9493 21252
rect -9620 21172 -9493 21188
rect -9620 21108 -9573 21172
rect -9509 21108 -9493 21172
rect -9620 21092 -9493 21108
rect -9620 21028 -9573 21092
rect -9509 21028 -9493 21092
rect -9620 21012 -9493 21028
rect -9620 20948 -9573 21012
rect -9509 20948 -9493 21012
rect -9620 20932 -9493 20948
rect -9620 20868 -9573 20932
rect -9509 20868 -9493 20932
rect -9620 20852 -9493 20868
rect -9620 20788 -9573 20852
rect -9509 20788 -9493 20852
rect -9620 20772 -9493 20788
rect -9620 20708 -9573 20772
rect -9509 20708 -9493 20772
rect -9620 20692 -9493 20708
rect -9620 20628 -9573 20692
rect -9509 20628 -9493 20692
rect -9620 20612 -9493 20628
rect -9620 20548 -9573 20612
rect -9509 20548 -9493 20612
rect -9620 20532 -9493 20548
rect -9620 20468 -9573 20532
rect -9509 20468 -9493 20532
rect -9620 20452 -9493 20468
rect -9620 20388 -9573 20452
rect -9509 20388 -9493 20452
rect -9620 20372 -9493 20388
rect -9620 20308 -9573 20372
rect -9509 20308 -9493 20372
rect -9620 20292 -9493 20308
rect -9620 20228 -9573 20292
rect -9509 20228 -9493 20292
rect -9620 20212 -9493 20228
rect -9620 20148 -9573 20212
rect -9509 20148 -9493 20212
rect -9620 20132 -9493 20148
rect -9620 20068 -9573 20132
rect -9509 20068 -9493 20132
rect -9620 20052 -9493 20068
rect -9620 19988 -9573 20052
rect -9509 19988 -9493 20052
rect -9620 19972 -9493 19988
rect -9620 19908 -9573 19972
rect -9509 19908 -9493 19972
rect -9620 19892 -9493 19908
rect -9620 19828 -9573 19892
rect -9509 19828 -9493 19892
rect -9620 19812 -9493 19828
rect -9620 19748 -9573 19812
rect -9509 19748 -9493 19812
rect -9620 19732 -9493 19748
rect -9620 19668 -9573 19732
rect -9509 19668 -9493 19732
rect -9620 19652 -9493 19668
rect -9620 19588 -9573 19652
rect -9509 19588 -9493 19652
rect -9620 19572 -9493 19588
rect -9620 19508 -9573 19572
rect -9509 19508 -9493 19572
rect -9620 19492 -9493 19508
rect -9620 19428 -9573 19492
rect -9509 19428 -9493 19492
rect -9620 19412 -9493 19428
rect -9620 19348 -9573 19412
rect -9509 19348 -9493 19412
rect -9620 19332 -9493 19348
rect -9620 19268 -9573 19332
rect -9509 19268 -9493 19332
rect -9620 19252 -9493 19268
rect -9620 19188 -9573 19252
rect -9509 19188 -9493 19252
rect -9620 19172 -9493 19188
rect -9620 19108 -9573 19172
rect -9509 19108 -9493 19172
rect -9620 19092 -9493 19108
rect -9620 19028 -9573 19092
rect -9509 19028 -9493 19092
rect -9620 19012 -9493 19028
rect -9620 18948 -9573 19012
rect -9509 18948 -9493 19012
rect -9620 18932 -9493 18948
rect -9620 18868 -9573 18932
rect -9509 18868 -9493 18932
rect -9620 18852 -9493 18868
rect -9620 18788 -9573 18852
rect -9509 18788 -9493 18852
rect -9620 18772 -9493 18788
rect -9620 18708 -9573 18772
rect -9509 18708 -9493 18772
rect -9620 18692 -9493 18708
rect -9620 18628 -9573 18692
rect -9509 18628 -9493 18692
rect -9620 18612 -9493 18628
rect -9620 18548 -9573 18612
rect -9509 18548 -9493 18612
rect -9620 18532 -9493 18548
rect -9620 18468 -9573 18532
rect -9509 18468 -9493 18532
rect -9620 18452 -9493 18468
rect -9620 18388 -9573 18452
rect -9509 18388 -9493 18452
rect -9620 18372 -9493 18388
rect -9620 18308 -9573 18372
rect -9509 18308 -9493 18372
rect -9620 18292 -9493 18308
rect -9620 18228 -9573 18292
rect -9509 18228 -9493 18292
rect -9620 18212 -9493 18228
rect -9620 18148 -9573 18212
rect -9509 18148 -9493 18212
rect -9620 18132 -9493 18148
rect -9620 18068 -9573 18132
rect -9509 18068 -9493 18132
rect -9620 18052 -9493 18068
rect -9620 17988 -9573 18052
rect -9509 17988 -9493 18052
rect -9620 17972 -9493 17988
rect -9620 17908 -9573 17972
rect -9509 17908 -9493 17972
rect -9620 17892 -9493 17908
rect -9620 17828 -9573 17892
rect -9509 17828 -9493 17892
rect -9620 17812 -9493 17828
rect -9620 17748 -9573 17812
rect -9509 17748 -9493 17812
rect -9620 17732 -9493 17748
rect -9620 17668 -9573 17732
rect -9509 17668 -9493 17732
rect -9620 17652 -9493 17668
rect -9620 17588 -9573 17652
rect -9509 17588 -9493 17652
rect -9620 17572 -9493 17588
rect -9620 17508 -9573 17572
rect -9509 17508 -9493 17572
rect -9620 17492 -9493 17508
rect -9620 17428 -9573 17492
rect -9509 17428 -9493 17492
rect -9620 17412 -9493 17428
rect -9620 17348 -9573 17412
rect -9509 17348 -9493 17412
rect -9620 17332 -9493 17348
rect -9620 17268 -9573 17332
rect -9509 17268 -9493 17332
rect -9620 17252 -9493 17268
rect -9620 17188 -9573 17252
rect -9509 17188 -9493 17252
rect -9620 17172 -9493 17188
rect -9620 17108 -9573 17172
rect -9509 17108 -9493 17172
rect -9620 17092 -9493 17108
rect -9620 17028 -9573 17092
rect -9509 17028 -9493 17092
rect -9620 17012 -9493 17028
rect -9620 16948 -9573 17012
rect -9509 16948 -9493 17012
rect -9620 16932 -9493 16948
rect -9620 16868 -9573 16932
rect -9509 16868 -9493 16932
rect -9620 16852 -9493 16868
rect -9620 16788 -9573 16852
rect -9509 16788 -9493 16852
rect -9620 16772 -9493 16788
rect -9620 16708 -9573 16772
rect -9509 16708 -9493 16772
rect -9620 16692 -9493 16708
rect -9620 16628 -9573 16692
rect -9509 16628 -9493 16692
rect -9620 16612 -9493 16628
rect -9620 16548 -9573 16612
rect -9509 16548 -9493 16612
rect -9620 16532 -9493 16548
rect -9620 16468 -9573 16532
rect -9509 16468 -9493 16532
rect -9620 16452 -9493 16468
rect -9620 16388 -9573 16452
rect -9509 16388 -9493 16452
rect -9620 16372 -9493 16388
rect -9620 16308 -9573 16372
rect -9509 16308 -9493 16372
rect -9620 16292 -9493 16308
rect -9620 16228 -9573 16292
rect -9509 16228 -9493 16292
rect -9620 16212 -9493 16228
rect -9620 16148 -9573 16212
rect -9509 16148 -9493 16212
rect -9620 16132 -9493 16148
rect -9620 16068 -9573 16132
rect -9509 16068 -9493 16132
rect -9620 16052 -9493 16068
rect -9620 15988 -9573 16052
rect -9509 15988 -9493 16052
rect -9620 15972 -9493 15988
rect -15939 15892 -15812 15908
rect -15939 15828 -15892 15892
rect -15828 15828 -15812 15892
rect -15939 15812 -15812 15828
rect -15939 15688 -15835 15812
rect -15939 15672 -15812 15688
rect -15939 15608 -15892 15672
rect -15828 15608 -15812 15672
rect -15939 15592 -15812 15608
rect -22258 15512 -22131 15528
rect -22258 15448 -22211 15512
rect -22147 15448 -22131 15512
rect -22258 15432 -22131 15448
rect -22258 15368 -22211 15432
rect -22147 15368 -22131 15432
rect -22258 15352 -22131 15368
rect -22258 15288 -22211 15352
rect -22147 15288 -22131 15352
rect -22258 15272 -22131 15288
rect -22258 15208 -22211 15272
rect -22147 15208 -22131 15272
rect -22258 15192 -22131 15208
rect -22258 15128 -22211 15192
rect -22147 15128 -22131 15192
rect -22258 15112 -22131 15128
rect -22258 15048 -22211 15112
rect -22147 15048 -22131 15112
rect -22258 15032 -22131 15048
rect -22258 14968 -22211 15032
rect -22147 14968 -22131 15032
rect -22258 14952 -22131 14968
rect -22258 14888 -22211 14952
rect -22147 14888 -22131 14952
rect -22258 14872 -22131 14888
rect -22258 14808 -22211 14872
rect -22147 14808 -22131 14872
rect -22258 14792 -22131 14808
rect -22258 14728 -22211 14792
rect -22147 14728 -22131 14792
rect -22258 14712 -22131 14728
rect -22258 14648 -22211 14712
rect -22147 14648 -22131 14712
rect -22258 14632 -22131 14648
rect -22258 14568 -22211 14632
rect -22147 14568 -22131 14632
rect -22258 14552 -22131 14568
rect -22258 14488 -22211 14552
rect -22147 14488 -22131 14552
rect -22258 14472 -22131 14488
rect -22258 14408 -22211 14472
rect -22147 14408 -22131 14472
rect -22258 14392 -22131 14408
rect -22258 14328 -22211 14392
rect -22147 14328 -22131 14392
rect -22258 14312 -22131 14328
rect -22258 14248 -22211 14312
rect -22147 14248 -22131 14312
rect -22258 14232 -22131 14248
rect -22258 14168 -22211 14232
rect -22147 14168 -22131 14232
rect -22258 14152 -22131 14168
rect -22258 14088 -22211 14152
rect -22147 14088 -22131 14152
rect -22258 14072 -22131 14088
rect -22258 14008 -22211 14072
rect -22147 14008 -22131 14072
rect -22258 13992 -22131 14008
rect -22258 13928 -22211 13992
rect -22147 13928 -22131 13992
rect -22258 13912 -22131 13928
rect -22258 13848 -22211 13912
rect -22147 13848 -22131 13912
rect -22258 13832 -22131 13848
rect -22258 13768 -22211 13832
rect -22147 13768 -22131 13832
rect -22258 13752 -22131 13768
rect -22258 13688 -22211 13752
rect -22147 13688 -22131 13752
rect -22258 13672 -22131 13688
rect -22258 13608 -22211 13672
rect -22147 13608 -22131 13672
rect -22258 13592 -22131 13608
rect -22258 13528 -22211 13592
rect -22147 13528 -22131 13592
rect -22258 13512 -22131 13528
rect -22258 13448 -22211 13512
rect -22147 13448 -22131 13512
rect -22258 13432 -22131 13448
rect -22258 13368 -22211 13432
rect -22147 13368 -22131 13432
rect -22258 13352 -22131 13368
rect -22258 13288 -22211 13352
rect -22147 13288 -22131 13352
rect -22258 13272 -22131 13288
rect -22258 13208 -22211 13272
rect -22147 13208 -22131 13272
rect -22258 13192 -22131 13208
rect -22258 13128 -22211 13192
rect -22147 13128 -22131 13192
rect -22258 13112 -22131 13128
rect -22258 13048 -22211 13112
rect -22147 13048 -22131 13112
rect -22258 13032 -22131 13048
rect -22258 12968 -22211 13032
rect -22147 12968 -22131 13032
rect -22258 12952 -22131 12968
rect -22258 12888 -22211 12952
rect -22147 12888 -22131 12952
rect -22258 12872 -22131 12888
rect -22258 12808 -22211 12872
rect -22147 12808 -22131 12872
rect -22258 12792 -22131 12808
rect -22258 12728 -22211 12792
rect -22147 12728 -22131 12792
rect -22258 12712 -22131 12728
rect -22258 12648 -22211 12712
rect -22147 12648 -22131 12712
rect -22258 12632 -22131 12648
rect -22258 12568 -22211 12632
rect -22147 12568 -22131 12632
rect -22258 12552 -22131 12568
rect -22258 12488 -22211 12552
rect -22147 12488 -22131 12552
rect -22258 12472 -22131 12488
rect -22258 12408 -22211 12472
rect -22147 12408 -22131 12472
rect -22258 12392 -22131 12408
rect -22258 12328 -22211 12392
rect -22147 12328 -22131 12392
rect -22258 12312 -22131 12328
rect -22258 12248 -22211 12312
rect -22147 12248 -22131 12312
rect -22258 12232 -22131 12248
rect -22258 12168 -22211 12232
rect -22147 12168 -22131 12232
rect -22258 12152 -22131 12168
rect -22258 12088 -22211 12152
rect -22147 12088 -22131 12152
rect -22258 12072 -22131 12088
rect -22258 12008 -22211 12072
rect -22147 12008 -22131 12072
rect -22258 11992 -22131 12008
rect -22258 11928 -22211 11992
rect -22147 11928 -22131 11992
rect -22258 11912 -22131 11928
rect -22258 11848 -22211 11912
rect -22147 11848 -22131 11912
rect -22258 11832 -22131 11848
rect -22258 11768 -22211 11832
rect -22147 11768 -22131 11832
rect -22258 11752 -22131 11768
rect -22258 11688 -22211 11752
rect -22147 11688 -22131 11752
rect -22258 11672 -22131 11688
rect -22258 11608 -22211 11672
rect -22147 11608 -22131 11672
rect -22258 11592 -22131 11608
rect -22258 11528 -22211 11592
rect -22147 11528 -22131 11592
rect -22258 11512 -22131 11528
rect -22258 11448 -22211 11512
rect -22147 11448 -22131 11512
rect -22258 11432 -22131 11448
rect -22258 11368 -22211 11432
rect -22147 11368 -22131 11432
rect -22258 11352 -22131 11368
rect -22258 11288 -22211 11352
rect -22147 11288 -22131 11352
rect -22258 11272 -22131 11288
rect -22258 11208 -22211 11272
rect -22147 11208 -22131 11272
rect -22258 11192 -22131 11208
rect -22258 11128 -22211 11192
rect -22147 11128 -22131 11192
rect -22258 11112 -22131 11128
rect -22258 11048 -22211 11112
rect -22147 11048 -22131 11112
rect -22258 11032 -22131 11048
rect -22258 10968 -22211 11032
rect -22147 10968 -22131 11032
rect -22258 10952 -22131 10968
rect -22258 10888 -22211 10952
rect -22147 10888 -22131 10952
rect -22258 10872 -22131 10888
rect -22258 10808 -22211 10872
rect -22147 10808 -22131 10872
rect -22258 10792 -22131 10808
rect -22258 10728 -22211 10792
rect -22147 10728 -22131 10792
rect -22258 10712 -22131 10728
rect -22258 10648 -22211 10712
rect -22147 10648 -22131 10712
rect -22258 10632 -22131 10648
rect -22258 10568 -22211 10632
rect -22147 10568 -22131 10632
rect -22258 10552 -22131 10568
rect -22258 10488 -22211 10552
rect -22147 10488 -22131 10552
rect -22258 10472 -22131 10488
rect -22258 10408 -22211 10472
rect -22147 10408 -22131 10472
rect -22258 10392 -22131 10408
rect -22258 10328 -22211 10392
rect -22147 10328 -22131 10392
rect -22258 10312 -22131 10328
rect -22258 10248 -22211 10312
rect -22147 10248 -22131 10312
rect -22258 10232 -22131 10248
rect -22258 10168 -22211 10232
rect -22147 10168 -22131 10232
rect -22258 10152 -22131 10168
rect -22258 10088 -22211 10152
rect -22147 10088 -22131 10152
rect -22258 10072 -22131 10088
rect -22258 10008 -22211 10072
rect -22147 10008 -22131 10072
rect -22258 9992 -22131 10008
rect -22258 9928 -22211 9992
rect -22147 9928 -22131 9992
rect -22258 9912 -22131 9928
rect -22258 9848 -22211 9912
rect -22147 9848 -22131 9912
rect -22258 9832 -22131 9848
rect -22258 9768 -22211 9832
rect -22147 9768 -22131 9832
rect -22258 9752 -22131 9768
rect -22258 9688 -22211 9752
rect -22147 9688 -22131 9752
rect -22258 9672 -22131 9688
rect -28577 9592 -28450 9608
rect -28577 9528 -28530 9592
rect -28466 9528 -28450 9592
rect -28577 9512 -28450 9528
rect -28577 9388 -28473 9512
rect -28577 9372 -28450 9388
rect -28577 9308 -28530 9372
rect -28466 9308 -28450 9372
rect -28577 9292 -28450 9308
rect -34896 9212 -34769 9228
rect -34896 9148 -34849 9212
rect -34785 9148 -34769 9212
rect -34896 9132 -34769 9148
rect -34896 9068 -34849 9132
rect -34785 9068 -34769 9132
rect -34896 9052 -34769 9068
rect -34896 8988 -34849 9052
rect -34785 8988 -34769 9052
rect -34896 8972 -34769 8988
rect -34896 8908 -34849 8972
rect -34785 8908 -34769 8972
rect -34896 8892 -34769 8908
rect -34896 8828 -34849 8892
rect -34785 8828 -34769 8892
rect -34896 8812 -34769 8828
rect -34896 8748 -34849 8812
rect -34785 8748 -34769 8812
rect -34896 8732 -34769 8748
rect -34896 8668 -34849 8732
rect -34785 8668 -34769 8732
rect -34896 8652 -34769 8668
rect -34896 8588 -34849 8652
rect -34785 8588 -34769 8652
rect -34896 8572 -34769 8588
rect -34896 8508 -34849 8572
rect -34785 8508 -34769 8572
rect -34896 8492 -34769 8508
rect -34896 8428 -34849 8492
rect -34785 8428 -34769 8492
rect -34896 8412 -34769 8428
rect -34896 8348 -34849 8412
rect -34785 8348 -34769 8412
rect -34896 8332 -34769 8348
rect -34896 8268 -34849 8332
rect -34785 8268 -34769 8332
rect -34896 8252 -34769 8268
rect -34896 8188 -34849 8252
rect -34785 8188 -34769 8252
rect -34896 8172 -34769 8188
rect -34896 8108 -34849 8172
rect -34785 8108 -34769 8172
rect -34896 8092 -34769 8108
rect -34896 8028 -34849 8092
rect -34785 8028 -34769 8092
rect -34896 8012 -34769 8028
rect -34896 7948 -34849 8012
rect -34785 7948 -34769 8012
rect -34896 7932 -34769 7948
rect -34896 7868 -34849 7932
rect -34785 7868 -34769 7932
rect -34896 7852 -34769 7868
rect -34896 7788 -34849 7852
rect -34785 7788 -34769 7852
rect -34896 7772 -34769 7788
rect -34896 7708 -34849 7772
rect -34785 7708 -34769 7772
rect -34896 7692 -34769 7708
rect -34896 7628 -34849 7692
rect -34785 7628 -34769 7692
rect -34896 7612 -34769 7628
rect -34896 7548 -34849 7612
rect -34785 7548 -34769 7612
rect -34896 7532 -34769 7548
rect -34896 7468 -34849 7532
rect -34785 7468 -34769 7532
rect -34896 7452 -34769 7468
rect -34896 7388 -34849 7452
rect -34785 7388 -34769 7452
rect -34896 7372 -34769 7388
rect -34896 7308 -34849 7372
rect -34785 7308 -34769 7372
rect -34896 7292 -34769 7308
rect -34896 7228 -34849 7292
rect -34785 7228 -34769 7292
rect -34896 7212 -34769 7228
rect -34896 7148 -34849 7212
rect -34785 7148 -34769 7212
rect -34896 7132 -34769 7148
rect -34896 7068 -34849 7132
rect -34785 7068 -34769 7132
rect -34896 7052 -34769 7068
rect -34896 6988 -34849 7052
rect -34785 6988 -34769 7052
rect -34896 6972 -34769 6988
rect -34896 6908 -34849 6972
rect -34785 6908 -34769 6972
rect -34896 6892 -34769 6908
rect -34896 6828 -34849 6892
rect -34785 6828 -34769 6892
rect -34896 6812 -34769 6828
rect -34896 6748 -34849 6812
rect -34785 6748 -34769 6812
rect -34896 6732 -34769 6748
rect -34896 6668 -34849 6732
rect -34785 6668 -34769 6732
rect -34896 6652 -34769 6668
rect -34896 6588 -34849 6652
rect -34785 6588 -34769 6652
rect -34896 6572 -34769 6588
rect -34896 6508 -34849 6572
rect -34785 6508 -34769 6572
rect -34896 6492 -34769 6508
rect -34896 6428 -34849 6492
rect -34785 6428 -34769 6492
rect -34896 6412 -34769 6428
rect -34896 6348 -34849 6412
rect -34785 6348 -34769 6412
rect -34896 6332 -34769 6348
rect -34896 6268 -34849 6332
rect -34785 6268 -34769 6332
rect -34896 6252 -34769 6268
rect -34896 6188 -34849 6252
rect -34785 6188 -34769 6252
rect -34896 6172 -34769 6188
rect -34896 6108 -34849 6172
rect -34785 6108 -34769 6172
rect -34896 6092 -34769 6108
rect -34896 6028 -34849 6092
rect -34785 6028 -34769 6092
rect -34896 6012 -34769 6028
rect -34896 5948 -34849 6012
rect -34785 5948 -34769 6012
rect -34896 5932 -34769 5948
rect -34896 5868 -34849 5932
rect -34785 5868 -34769 5932
rect -34896 5852 -34769 5868
rect -34896 5788 -34849 5852
rect -34785 5788 -34769 5852
rect -34896 5772 -34769 5788
rect -34896 5708 -34849 5772
rect -34785 5708 -34769 5772
rect -34896 5692 -34769 5708
rect -34896 5628 -34849 5692
rect -34785 5628 -34769 5692
rect -34896 5612 -34769 5628
rect -34896 5548 -34849 5612
rect -34785 5548 -34769 5612
rect -34896 5532 -34769 5548
rect -34896 5468 -34849 5532
rect -34785 5468 -34769 5532
rect -34896 5452 -34769 5468
rect -34896 5388 -34849 5452
rect -34785 5388 -34769 5452
rect -34896 5372 -34769 5388
rect -34896 5308 -34849 5372
rect -34785 5308 -34769 5372
rect -34896 5292 -34769 5308
rect -34896 5228 -34849 5292
rect -34785 5228 -34769 5292
rect -34896 5212 -34769 5228
rect -34896 5148 -34849 5212
rect -34785 5148 -34769 5212
rect -34896 5132 -34769 5148
rect -34896 5068 -34849 5132
rect -34785 5068 -34769 5132
rect -34896 5052 -34769 5068
rect -34896 4988 -34849 5052
rect -34785 4988 -34769 5052
rect -34896 4972 -34769 4988
rect -34896 4908 -34849 4972
rect -34785 4908 -34769 4972
rect -34896 4892 -34769 4908
rect -34896 4828 -34849 4892
rect -34785 4828 -34769 4892
rect -34896 4812 -34769 4828
rect -34896 4748 -34849 4812
rect -34785 4748 -34769 4812
rect -34896 4732 -34769 4748
rect -34896 4668 -34849 4732
rect -34785 4668 -34769 4732
rect -34896 4652 -34769 4668
rect -34896 4588 -34849 4652
rect -34785 4588 -34769 4652
rect -34896 4572 -34769 4588
rect -34896 4508 -34849 4572
rect -34785 4508 -34769 4572
rect -34896 4492 -34769 4508
rect -34896 4428 -34849 4492
rect -34785 4428 -34769 4492
rect -34896 4412 -34769 4428
rect -34896 4348 -34849 4412
rect -34785 4348 -34769 4412
rect -34896 4332 -34769 4348
rect -34896 4268 -34849 4332
rect -34785 4268 -34769 4332
rect -34896 4252 -34769 4268
rect -34896 4188 -34849 4252
rect -34785 4188 -34769 4252
rect -34896 4172 -34769 4188
rect -34896 4108 -34849 4172
rect -34785 4108 -34769 4172
rect -34896 4092 -34769 4108
rect -34896 4028 -34849 4092
rect -34785 4028 -34769 4092
rect -34896 4012 -34769 4028
rect -34896 3948 -34849 4012
rect -34785 3948 -34769 4012
rect -34896 3932 -34769 3948
rect -34896 3868 -34849 3932
rect -34785 3868 -34769 3932
rect -34896 3852 -34769 3868
rect -34896 3788 -34849 3852
rect -34785 3788 -34769 3852
rect -34896 3772 -34769 3788
rect -34896 3708 -34849 3772
rect -34785 3708 -34769 3772
rect -34896 3692 -34769 3708
rect -34896 3628 -34849 3692
rect -34785 3628 -34769 3692
rect -34896 3612 -34769 3628
rect -34896 3548 -34849 3612
rect -34785 3548 -34769 3612
rect -34896 3532 -34769 3548
rect -34896 3468 -34849 3532
rect -34785 3468 -34769 3532
rect -34896 3452 -34769 3468
rect -34896 3388 -34849 3452
rect -34785 3388 -34769 3452
rect -34896 3372 -34769 3388
rect -41215 3292 -41088 3308
rect -41215 3228 -41168 3292
rect -41104 3228 -41088 3292
rect -41215 3212 -41088 3228
rect -41215 3088 -41111 3212
rect -41215 3072 -41088 3088
rect -41215 3008 -41168 3072
rect -41104 3008 -41088 3072
rect -41215 2992 -41088 3008
rect -47244 2952 -41322 2961
rect -47244 -2952 -47235 2952
rect -41331 -2952 -41322 2952
rect -47244 -2961 -41322 -2952
rect -41215 2928 -41168 2992
rect -41104 2928 -41088 2992
rect -38016 2961 -37912 3339
rect -34896 3308 -34849 3372
rect -34785 3308 -34769 3372
rect -34606 9252 -28684 9261
rect -34606 3348 -34597 9252
rect -28693 3348 -28684 9252
rect -34606 3339 -28684 3348
rect -28577 9228 -28530 9292
rect -28466 9228 -28450 9292
rect -25378 9261 -25274 9639
rect -22258 9608 -22211 9672
rect -22147 9608 -22131 9672
rect -21968 15552 -16046 15561
rect -21968 9648 -21959 15552
rect -16055 9648 -16046 15552
rect -21968 9639 -16046 9648
rect -15939 15528 -15892 15592
rect -15828 15528 -15812 15592
rect -12740 15561 -12636 15939
rect -9620 15908 -9573 15972
rect -9509 15908 -9493 15972
rect -9330 21852 -3408 21861
rect -9330 15948 -9321 21852
rect -3417 15948 -3408 21852
rect -9330 15939 -3408 15948
rect -3301 21828 -3254 21892
rect -3190 21828 -3174 21892
rect -102 21861 2 22239
rect 3018 22208 3065 22272
rect 3129 22208 3145 22272
rect 3308 28152 9230 28161
rect 3308 22248 3317 28152
rect 9221 22248 9230 28152
rect 3308 22239 9230 22248
rect 9337 28128 9384 28192
rect 9448 28128 9464 28192
rect 12536 28161 12640 28539
rect 15656 28508 15703 28572
rect 15767 28508 15783 28572
rect 15946 34452 21868 34461
rect 15946 28548 15955 34452
rect 21859 28548 21868 34452
rect 15946 28539 21868 28548
rect 21975 34428 22022 34492
rect 22086 34428 22102 34492
rect 25174 34461 25278 34839
rect 28294 34808 28341 34872
rect 28405 34808 28421 34872
rect 28584 40752 34506 40761
rect 28584 34848 28593 40752
rect 34497 34848 34506 40752
rect 28584 34839 34506 34848
rect 34613 40728 34660 40792
rect 34724 40728 34740 40792
rect 37812 40761 37916 41139
rect 40932 41108 40979 41172
rect 41043 41108 41059 41172
rect 41222 47052 47144 47061
rect 41222 41148 41231 47052
rect 47135 41148 47144 47052
rect 41222 41139 47144 41148
rect 47251 47028 47298 47092
rect 47362 47028 47378 47092
rect 47251 47012 47378 47028
rect 47251 46948 47298 47012
rect 47362 46948 47378 47012
rect 47251 46932 47378 46948
rect 47251 46868 47298 46932
rect 47362 46868 47378 46932
rect 47251 46852 47378 46868
rect 47251 46788 47298 46852
rect 47362 46788 47378 46852
rect 47251 46772 47378 46788
rect 47251 46708 47298 46772
rect 47362 46708 47378 46772
rect 47251 46692 47378 46708
rect 47251 46628 47298 46692
rect 47362 46628 47378 46692
rect 47251 46612 47378 46628
rect 47251 46548 47298 46612
rect 47362 46548 47378 46612
rect 47251 46532 47378 46548
rect 47251 46468 47298 46532
rect 47362 46468 47378 46532
rect 47251 46452 47378 46468
rect 47251 46388 47298 46452
rect 47362 46388 47378 46452
rect 47251 46372 47378 46388
rect 47251 46308 47298 46372
rect 47362 46308 47378 46372
rect 47251 46292 47378 46308
rect 47251 46228 47298 46292
rect 47362 46228 47378 46292
rect 47251 46212 47378 46228
rect 47251 46148 47298 46212
rect 47362 46148 47378 46212
rect 47251 46132 47378 46148
rect 47251 46068 47298 46132
rect 47362 46068 47378 46132
rect 47251 46052 47378 46068
rect 47251 45988 47298 46052
rect 47362 45988 47378 46052
rect 47251 45972 47378 45988
rect 47251 45908 47298 45972
rect 47362 45908 47378 45972
rect 47251 45892 47378 45908
rect 47251 45828 47298 45892
rect 47362 45828 47378 45892
rect 47251 45812 47378 45828
rect 47251 45748 47298 45812
rect 47362 45748 47378 45812
rect 47251 45732 47378 45748
rect 47251 45668 47298 45732
rect 47362 45668 47378 45732
rect 47251 45652 47378 45668
rect 47251 45588 47298 45652
rect 47362 45588 47378 45652
rect 47251 45572 47378 45588
rect 47251 45508 47298 45572
rect 47362 45508 47378 45572
rect 47251 45492 47378 45508
rect 47251 45428 47298 45492
rect 47362 45428 47378 45492
rect 47251 45412 47378 45428
rect 47251 45348 47298 45412
rect 47362 45348 47378 45412
rect 47251 45332 47378 45348
rect 47251 45268 47298 45332
rect 47362 45268 47378 45332
rect 47251 45252 47378 45268
rect 47251 45188 47298 45252
rect 47362 45188 47378 45252
rect 47251 45172 47378 45188
rect 47251 45108 47298 45172
rect 47362 45108 47378 45172
rect 47251 45092 47378 45108
rect 47251 45028 47298 45092
rect 47362 45028 47378 45092
rect 47251 45012 47378 45028
rect 47251 44948 47298 45012
rect 47362 44948 47378 45012
rect 47251 44932 47378 44948
rect 47251 44868 47298 44932
rect 47362 44868 47378 44932
rect 47251 44852 47378 44868
rect 47251 44788 47298 44852
rect 47362 44788 47378 44852
rect 47251 44772 47378 44788
rect 47251 44708 47298 44772
rect 47362 44708 47378 44772
rect 47251 44692 47378 44708
rect 47251 44628 47298 44692
rect 47362 44628 47378 44692
rect 47251 44612 47378 44628
rect 47251 44548 47298 44612
rect 47362 44548 47378 44612
rect 47251 44532 47378 44548
rect 47251 44468 47298 44532
rect 47362 44468 47378 44532
rect 47251 44452 47378 44468
rect 47251 44388 47298 44452
rect 47362 44388 47378 44452
rect 47251 44372 47378 44388
rect 47251 44308 47298 44372
rect 47362 44308 47378 44372
rect 47251 44292 47378 44308
rect 47251 44228 47298 44292
rect 47362 44228 47378 44292
rect 47251 44212 47378 44228
rect 47251 44148 47298 44212
rect 47362 44148 47378 44212
rect 47251 44132 47378 44148
rect 47251 44068 47298 44132
rect 47362 44068 47378 44132
rect 47251 44052 47378 44068
rect 47251 43988 47298 44052
rect 47362 43988 47378 44052
rect 47251 43972 47378 43988
rect 47251 43908 47298 43972
rect 47362 43908 47378 43972
rect 47251 43892 47378 43908
rect 47251 43828 47298 43892
rect 47362 43828 47378 43892
rect 47251 43812 47378 43828
rect 47251 43748 47298 43812
rect 47362 43748 47378 43812
rect 47251 43732 47378 43748
rect 47251 43668 47298 43732
rect 47362 43668 47378 43732
rect 47251 43652 47378 43668
rect 47251 43588 47298 43652
rect 47362 43588 47378 43652
rect 47251 43572 47378 43588
rect 47251 43508 47298 43572
rect 47362 43508 47378 43572
rect 47251 43492 47378 43508
rect 47251 43428 47298 43492
rect 47362 43428 47378 43492
rect 47251 43412 47378 43428
rect 47251 43348 47298 43412
rect 47362 43348 47378 43412
rect 47251 43332 47378 43348
rect 47251 43268 47298 43332
rect 47362 43268 47378 43332
rect 47251 43252 47378 43268
rect 47251 43188 47298 43252
rect 47362 43188 47378 43252
rect 47251 43172 47378 43188
rect 47251 43108 47298 43172
rect 47362 43108 47378 43172
rect 47251 43092 47378 43108
rect 47251 43028 47298 43092
rect 47362 43028 47378 43092
rect 47251 43012 47378 43028
rect 47251 42948 47298 43012
rect 47362 42948 47378 43012
rect 47251 42932 47378 42948
rect 47251 42868 47298 42932
rect 47362 42868 47378 42932
rect 47251 42852 47378 42868
rect 47251 42788 47298 42852
rect 47362 42788 47378 42852
rect 47251 42772 47378 42788
rect 47251 42708 47298 42772
rect 47362 42708 47378 42772
rect 47251 42692 47378 42708
rect 47251 42628 47298 42692
rect 47362 42628 47378 42692
rect 47251 42612 47378 42628
rect 47251 42548 47298 42612
rect 47362 42548 47378 42612
rect 47251 42532 47378 42548
rect 47251 42468 47298 42532
rect 47362 42468 47378 42532
rect 47251 42452 47378 42468
rect 47251 42388 47298 42452
rect 47362 42388 47378 42452
rect 47251 42372 47378 42388
rect 47251 42308 47298 42372
rect 47362 42308 47378 42372
rect 47251 42292 47378 42308
rect 47251 42228 47298 42292
rect 47362 42228 47378 42292
rect 47251 42212 47378 42228
rect 47251 42148 47298 42212
rect 47362 42148 47378 42212
rect 47251 42132 47378 42148
rect 47251 42068 47298 42132
rect 47362 42068 47378 42132
rect 47251 42052 47378 42068
rect 47251 41988 47298 42052
rect 47362 41988 47378 42052
rect 47251 41972 47378 41988
rect 47251 41908 47298 41972
rect 47362 41908 47378 41972
rect 47251 41892 47378 41908
rect 47251 41828 47298 41892
rect 47362 41828 47378 41892
rect 47251 41812 47378 41828
rect 47251 41748 47298 41812
rect 47362 41748 47378 41812
rect 47251 41732 47378 41748
rect 47251 41668 47298 41732
rect 47362 41668 47378 41732
rect 47251 41652 47378 41668
rect 47251 41588 47298 41652
rect 47362 41588 47378 41652
rect 47251 41572 47378 41588
rect 47251 41508 47298 41572
rect 47362 41508 47378 41572
rect 47251 41492 47378 41508
rect 47251 41428 47298 41492
rect 47362 41428 47378 41492
rect 47251 41412 47378 41428
rect 47251 41348 47298 41412
rect 47362 41348 47378 41412
rect 47251 41332 47378 41348
rect 47251 41268 47298 41332
rect 47362 41268 47378 41332
rect 47251 41252 47378 41268
rect 47251 41188 47298 41252
rect 47362 41188 47378 41252
rect 47251 41172 47378 41188
rect 40932 41092 41059 41108
rect 40932 41028 40979 41092
rect 41043 41028 41059 41092
rect 40932 41012 41059 41028
rect 40932 40888 41036 41012
rect 40932 40872 41059 40888
rect 40932 40808 40979 40872
rect 41043 40808 41059 40872
rect 40932 40792 41059 40808
rect 34613 40712 34740 40728
rect 34613 40648 34660 40712
rect 34724 40648 34740 40712
rect 34613 40632 34740 40648
rect 34613 40568 34660 40632
rect 34724 40568 34740 40632
rect 34613 40552 34740 40568
rect 34613 40488 34660 40552
rect 34724 40488 34740 40552
rect 34613 40472 34740 40488
rect 34613 40408 34660 40472
rect 34724 40408 34740 40472
rect 34613 40392 34740 40408
rect 34613 40328 34660 40392
rect 34724 40328 34740 40392
rect 34613 40312 34740 40328
rect 34613 40248 34660 40312
rect 34724 40248 34740 40312
rect 34613 40232 34740 40248
rect 34613 40168 34660 40232
rect 34724 40168 34740 40232
rect 34613 40152 34740 40168
rect 34613 40088 34660 40152
rect 34724 40088 34740 40152
rect 34613 40072 34740 40088
rect 34613 40008 34660 40072
rect 34724 40008 34740 40072
rect 34613 39992 34740 40008
rect 34613 39928 34660 39992
rect 34724 39928 34740 39992
rect 34613 39912 34740 39928
rect 34613 39848 34660 39912
rect 34724 39848 34740 39912
rect 34613 39832 34740 39848
rect 34613 39768 34660 39832
rect 34724 39768 34740 39832
rect 34613 39752 34740 39768
rect 34613 39688 34660 39752
rect 34724 39688 34740 39752
rect 34613 39672 34740 39688
rect 34613 39608 34660 39672
rect 34724 39608 34740 39672
rect 34613 39592 34740 39608
rect 34613 39528 34660 39592
rect 34724 39528 34740 39592
rect 34613 39512 34740 39528
rect 34613 39448 34660 39512
rect 34724 39448 34740 39512
rect 34613 39432 34740 39448
rect 34613 39368 34660 39432
rect 34724 39368 34740 39432
rect 34613 39352 34740 39368
rect 34613 39288 34660 39352
rect 34724 39288 34740 39352
rect 34613 39272 34740 39288
rect 34613 39208 34660 39272
rect 34724 39208 34740 39272
rect 34613 39192 34740 39208
rect 34613 39128 34660 39192
rect 34724 39128 34740 39192
rect 34613 39112 34740 39128
rect 34613 39048 34660 39112
rect 34724 39048 34740 39112
rect 34613 39032 34740 39048
rect 34613 38968 34660 39032
rect 34724 38968 34740 39032
rect 34613 38952 34740 38968
rect 34613 38888 34660 38952
rect 34724 38888 34740 38952
rect 34613 38872 34740 38888
rect 34613 38808 34660 38872
rect 34724 38808 34740 38872
rect 34613 38792 34740 38808
rect 34613 38728 34660 38792
rect 34724 38728 34740 38792
rect 34613 38712 34740 38728
rect 34613 38648 34660 38712
rect 34724 38648 34740 38712
rect 34613 38632 34740 38648
rect 34613 38568 34660 38632
rect 34724 38568 34740 38632
rect 34613 38552 34740 38568
rect 34613 38488 34660 38552
rect 34724 38488 34740 38552
rect 34613 38472 34740 38488
rect 34613 38408 34660 38472
rect 34724 38408 34740 38472
rect 34613 38392 34740 38408
rect 34613 38328 34660 38392
rect 34724 38328 34740 38392
rect 34613 38312 34740 38328
rect 34613 38248 34660 38312
rect 34724 38248 34740 38312
rect 34613 38232 34740 38248
rect 34613 38168 34660 38232
rect 34724 38168 34740 38232
rect 34613 38152 34740 38168
rect 34613 38088 34660 38152
rect 34724 38088 34740 38152
rect 34613 38072 34740 38088
rect 34613 38008 34660 38072
rect 34724 38008 34740 38072
rect 34613 37992 34740 38008
rect 34613 37928 34660 37992
rect 34724 37928 34740 37992
rect 34613 37912 34740 37928
rect 34613 37848 34660 37912
rect 34724 37848 34740 37912
rect 34613 37832 34740 37848
rect 34613 37768 34660 37832
rect 34724 37768 34740 37832
rect 34613 37752 34740 37768
rect 34613 37688 34660 37752
rect 34724 37688 34740 37752
rect 34613 37672 34740 37688
rect 34613 37608 34660 37672
rect 34724 37608 34740 37672
rect 34613 37592 34740 37608
rect 34613 37528 34660 37592
rect 34724 37528 34740 37592
rect 34613 37512 34740 37528
rect 34613 37448 34660 37512
rect 34724 37448 34740 37512
rect 34613 37432 34740 37448
rect 34613 37368 34660 37432
rect 34724 37368 34740 37432
rect 34613 37352 34740 37368
rect 34613 37288 34660 37352
rect 34724 37288 34740 37352
rect 34613 37272 34740 37288
rect 34613 37208 34660 37272
rect 34724 37208 34740 37272
rect 34613 37192 34740 37208
rect 34613 37128 34660 37192
rect 34724 37128 34740 37192
rect 34613 37112 34740 37128
rect 34613 37048 34660 37112
rect 34724 37048 34740 37112
rect 34613 37032 34740 37048
rect 34613 36968 34660 37032
rect 34724 36968 34740 37032
rect 34613 36952 34740 36968
rect 34613 36888 34660 36952
rect 34724 36888 34740 36952
rect 34613 36872 34740 36888
rect 34613 36808 34660 36872
rect 34724 36808 34740 36872
rect 34613 36792 34740 36808
rect 34613 36728 34660 36792
rect 34724 36728 34740 36792
rect 34613 36712 34740 36728
rect 34613 36648 34660 36712
rect 34724 36648 34740 36712
rect 34613 36632 34740 36648
rect 34613 36568 34660 36632
rect 34724 36568 34740 36632
rect 34613 36552 34740 36568
rect 34613 36488 34660 36552
rect 34724 36488 34740 36552
rect 34613 36472 34740 36488
rect 34613 36408 34660 36472
rect 34724 36408 34740 36472
rect 34613 36392 34740 36408
rect 34613 36328 34660 36392
rect 34724 36328 34740 36392
rect 34613 36312 34740 36328
rect 34613 36248 34660 36312
rect 34724 36248 34740 36312
rect 34613 36232 34740 36248
rect 34613 36168 34660 36232
rect 34724 36168 34740 36232
rect 34613 36152 34740 36168
rect 34613 36088 34660 36152
rect 34724 36088 34740 36152
rect 34613 36072 34740 36088
rect 34613 36008 34660 36072
rect 34724 36008 34740 36072
rect 34613 35992 34740 36008
rect 34613 35928 34660 35992
rect 34724 35928 34740 35992
rect 34613 35912 34740 35928
rect 34613 35848 34660 35912
rect 34724 35848 34740 35912
rect 34613 35832 34740 35848
rect 34613 35768 34660 35832
rect 34724 35768 34740 35832
rect 34613 35752 34740 35768
rect 34613 35688 34660 35752
rect 34724 35688 34740 35752
rect 34613 35672 34740 35688
rect 34613 35608 34660 35672
rect 34724 35608 34740 35672
rect 34613 35592 34740 35608
rect 34613 35528 34660 35592
rect 34724 35528 34740 35592
rect 34613 35512 34740 35528
rect 34613 35448 34660 35512
rect 34724 35448 34740 35512
rect 34613 35432 34740 35448
rect 34613 35368 34660 35432
rect 34724 35368 34740 35432
rect 34613 35352 34740 35368
rect 34613 35288 34660 35352
rect 34724 35288 34740 35352
rect 34613 35272 34740 35288
rect 34613 35208 34660 35272
rect 34724 35208 34740 35272
rect 34613 35192 34740 35208
rect 34613 35128 34660 35192
rect 34724 35128 34740 35192
rect 34613 35112 34740 35128
rect 34613 35048 34660 35112
rect 34724 35048 34740 35112
rect 34613 35032 34740 35048
rect 34613 34968 34660 35032
rect 34724 34968 34740 35032
rect 34613 34952 34740 34968
rect 34613 34888 34660 34952
rect 34724 34888 34740 34952
rect 34613 34872 34740 34888
rect 28294 34792 28421 34808
rect 28294 34728 28341 34792
rect 28405 34728 28421 34792
rect 28294 34712 28421 34728
rect 28294 34588 28398 34712
rect 28294 34572 28421 34588
rect 28294 34508 28341 34572
rect 28405 34508 28421 34572
rect 28294 34492 28421 34508
rect 21975 34412 22102 34428
rect 21975 34348 22022 34412
rect 22086 34348 22102 34412
rect 21975 34332 22102 34348
rect 21975 34268 22022 34332
rect 22086 34268 22102 34332
rect 21975 34252 22102 34268
rect 21975 34188 22022 34252
rect 22086 34188 22102 34252
rect 21975 34172 22102 34188
rect 21975 34108 22022 34172
rect 22086 34108 22102 34172
rect 21975 34092 22102 34108
rect 21975 34028 22022 34092
rect 22086 34028 22102 34092
rect 21975 34012 22102 34028
rect 21975 33948 22022 34012
rect 22086 33948 22102 34012
rect 21975 33932 22102 33948
rect 21975 33868 22022 33932
rect 22086 33868 22102 33932
rect 21975 33852 22102 33868
rect 21975 33788 22022 33852
rect 22086 33788 22102 33852
rect 21975 33772 22102 33788
rect 21975 33708 22022 33772
rect 22086 33708 22102 33772
rect 21975 33692 22102 33708
rect 21975 33628 22022 33692
rect 22086 33628 22102 33692
rect 21975 33612 22102 33628
rect 21975 33548 22022 33612
rect 22086 33548 22102 33612
rect 21975 33532 22102 33548
rect 21975 33468 22022 33532
rect 22086 33468 22102 33532
rect 21975 33452 22102 33468
rect 21975 33388 22022 33452
rect 22086 33388 22102 33452
rect 21975 33372 22102 33388
rect 21975 33308 22022 33372
rect 22086 33308 22102 33372
rect 21975 33292 22102 33308
rect 21975 33228 22022 33292
rect 22086 33228 22102 33292
rect 21975 33212 22102 33228
rect 21975 33148 22022 33212
rect 22086 33148 22102 33212
rect 21975 33132 22102 33148
rect 21975 33068 22022 33132
rect 22086 33068 22102 33132
rect 21975 33052 22102 33068
rect 21975 32988 22022 33052
rect 22086 32988 22102 33052
rect 21975 32972 22102 32988
rect 21975 32908 22022 32972
rect 22086 32908 22102 32972
rect 21975 32892 22102 32908
rect 21975 32828 22022 32892
rect 22086 32828 22102 32892
rect 21975 32812 22102 32828
rect 21975 32748 22022 32812
rect 22086 32748 22102 32812
rect 21975 32732 22102 32748
rect 21975 32668 22022 32732
rect 22086 32668 22102 32732
rect 21975 32652 22102 32668
rect 21975 32588 22022 32652
rect 22086 32588 22102 32652
rect 21975 32572 22102 32588
rect 21975 32508 22022 32572
rect 22086 32508 22102 32572
rect 21975 32492 22102 32508
rect 21975 32428 22022 32492
rect 22086 32428 22102 32492
rect 21975 32412 22102 32428
rect 21975 32348 22022 32412
rect 22086 32348 22102 32412
rect 21975 32332 22102 32348
rect 21975 32268 22022 32332
rect 22086 32268 22102 32332
rect 21975 32252 22102 32268
rect 21975 32188 22022 32252
rect 22086 32188 22102 32252
rect 21975 32172 22102 32188
rect 21975 32108 22022 32172
rect 22086 32108 22102 32172
rect 21975 32092 22102 32108
rect 21975 32028 22022 32092
rect 22086 32028 22102 32092
rect 21975 32012 22102 32028
rect 21975 31948 22022 32012
rect 22086 31948 22102 32012
rect 21975 31932 22102 31948
rect 21975 31868 22022 31932
rect 22086 31868 22102 31932
rect 21975 31852 22102 31868
rect 21975 31788 22022 31852
rect 22086 31788 22102 31852
rect 21975 31772 22102 31788
rect 21975 31708 22022 31772
rect 22086 31708 22102 31772
rect 21975 31692 22102 31708
rect 21975 31628 22022 31692
rect 22086 31628 22102 31692
rect 21975 31612 22102 31628
rect 21975 31548 22022 31612
rect 22086 31548 22102 31612
rect 21975 31532 22102 31548
rect 21975 31468 22022 31532
rect 22086 31468 22102 31532
rect 21975 31452 22102 31468
rect 21975 31388 22022 31452
rect 22086 31388 22102 31452
rect 21975 31372 22102 31388
rect 21975 31308 22022 31372
rect 22086 31308 22102 31372
rect 21975 31292 22102 31308
rect 21975 31228 22022 31292
rect 22086 31228 22102 31292
rect 21975 31212 22102 31228
rect 21975 31148 22022 31212
rect 22086 31148 22102 31212
rect 21975 31132 22102 31148
rect 21975 31068 22022 31132
rect 22086 31068 22102 31132
rect 21975 31052 22102 31068
rect 21975 30988 22022 31052
rect 22086 30988 22102 31052
rect 21975 30972 22102 30988
rect 21975 30908 22022 30972
rect 22086 30908 22102 30972
rect 21975 30892 22102 30908
rect 21975 30828 22022 30892
rect 22086 30828 22102 30892
rect 21975 30812 22102 30828
rect 21975 30748 22022 30812
rect 22086 30748 22102 30812
rect 21975 30732 22102 30748
rect 21975 30668 22022 30732
rect 22086 30668 22102 30732
rect 21975 30652 22102 30668
rect 21975 30588 22022 30652
rect 22086 30588 22102 30652
rect 21975 30572 22102 30588
rect 21975 30508 22022 30572
rect 22086 30508 22102 30572
rect 21975 30492 22102 30508
rect 21975 30428 22022 30492
rect 22086 30428 22102 30492
rect 21975 30412 22102 30428
rect 21975 30348 22022 30412
rect 22086 30348 22102 30412
rect 21975 30332 22102 30348
rect 21975 30268 22022 30332
rect 22086 30268 22102 30332
rect 21975 30252 22102 30268
rect 21975 30188 22022 30252
rect 22086 30188 22102 30252
rect 21975 30172 22102 30188
rect 21975 30108 22022 30172
rect 22086 30108 22102 30172
rect 21975 30092 22102 30108
rect 21975 30028 22022 30092
rect 22086 30028 22102 30092
rect 21975 30012 22102 30028
rect 21975 29948 22022 30012
rect 22086 29948 22102 30012
rect 21975 29932 22102 29948
rect 21975 29868 22022 29932
rect 22086 29868 22102 29932
rect 21975 29852 22102 29868
rect 21975 29788 22022 29852
rect 22086 29788 22102 29852
rect 21975 29772 22102 29788
rect 21975 29708 22022 29772
rect 22086 29708 22102 29772
rect 21975 29692 22102 29708
rect 21975 29628 22022 29692
rect 22086 29628 22102 29692
rect 21975 29612 22102 29628
rect 21975 29548 22022 29612
rect 22086 29548 22102 29612
rect 21975 29532 22102 29548
rect 21975 29468 22022 29532
rect 22086 29468 22102 29532
rect 21975 29452 22102 29468
rect 21975 29388 22022 29452
rect 22086 29388 22102 29452
rect 21975 29372 22102 29388
rect 21975 29308 22022 29372
rect 22086 29308 22102 29372
rect 21975 29292 22102 29308
rect 21975 29228 22022 29292
rect 22086 29228 22102 29292
rect 21975 29212 22102 29228
rect 21975 29148 22022 29212
rect 22086 29148 22102 29212
rect 21975 29132 22102 29148
rect 21975 29068 22022 29132
rect 22086 29068 22102 29132
rect 21975 29052 22102 29068
rect 21975 28988 22022 29052
rect 22086 28988 22102 29052
rect 21975 28972 22102 28988
rect 21975 28908 22022 28972
rect 22086 28908 22102 28972
rect 21975 28892 22102 28908
rect 21975 28828 22022 28892
rect 22086 28828 22102 28892
rect 21975 28812 22102 28828
rect 21975 28748 22022 28812
rect 22086 28748 22102 28812
rect 21975 28732 22102 28748
rect 21975 28668 22022 28732
rect 22086 28668 22102 28732
rect 21975 28652 22102 28668
rect 21975 28588 22022 28652
rect 22086 28588 22102 28652
rect 21975 28572 22102 28588
rect 15656 28492 15783 28508
rect 15656 28428 15703 28492
rect 15767 28428 15783 28492
rect 15656 28412 15783 28428
rect 15656 28288 15760 28412
rect 15656 28272 15783 28288
rect 15656 28208 15703 28272
rect 15767 28208 15783 28272
rect 15656 28192 15783 28208
rect 9337 28112 9464 28128
rect 9337 28048 9384 28112
rect 9448 28048 9464 28112
rect 9337 28032 9464 28048
rect 9337 27968 9384 28032
rect 9448 27968 9464 28032
rect 9337 27952 9464 27968
rect 9337 27888 9384 27952
rect 9448 27888 9464 27952
rect 9337 27872 9464 27888
rect 9337 27808 9384 27872
rect 9448 27808 9464 27872
rect 9337 27792 9464 27808
rect 9337 27728 9384 27792
rect 9448 27728 9464 27792
rect 9337 27712 9464 27728
rect 9337 27648 9384 27712
rect 9448 27648 9464 27712
rect 9337 27632 9464 27648
rect 9337 27568 9384 27632
rect 9448 27568 9464 27632
rect 9337 27552 9464 27568
rect 9337 27488 9384 27552
rect 9448 27488 9464 27552
rect 9337 27472 9464 27488
rect 9337 27408 9384 27472
rect 9448 27408 9464 27472
rect 9337 27392 9464 27408
rect 9337 27328 9384 27392
rect 9448 27328 9464 27392
rect 9337 27312 9464 27328
rect 9337 27248 9384 27312
rect 9448 27248 9464 27312
rect 9337 27232 9464 27248
rect 9337 27168 9384 27232
rect 9448 27168 9464 27232
rect 9337 27152 9464 27168
rect 9337 27088 9384 27152
rect 9448 27088 9464 27152
rect 9337 27072 9464 27088
rect 9337 27008 9384 27072
rect 9448 27008 9464 27072
rect 9337 26992 9464 27008
rect 9337 26928 9384 26992
rect 9448 26928 9464 26992
rect 9337 26912 9464 26928
rect 9337 26848 9384 26912
rect 9448 26848 9464 26912
rect 9337 26832 9464 26848
rect 9337 26768 9384 26832
rect 9448 26768 9464 26832
rect 9337 26752 9464 26768
rect 9337 26688 9384 26752
rect 9448 26688 9464 26752
rect 9337 26672 9464 26688
rect 9337 26608 9384 26672
rect 9448 26608 9464 26672
rect 9337 26592 9464 26608
rect 9337 26528 9384 26592
rect 9448 26528 9464 26592
rect 9337 26512 9464 26528
rect 9337 26448 9384 26512
rect 9448 26448 9464 26512
rect 9337 26432 9464 26448
rect 9337 26368 9384 26432
rect 9448 26368 9464 26432
rect 9337 26352 9464 26368
rect 9337 26288 9384 26352
rect 9448 26288 9464 26352
rect 9337 26272 9464 26288
rect 9337 26208 9384 26272
rect 9448 26208 9464 26272
rect 9337 26192 9464 26208
rect 9337 26128 9384 26192
rect 9448 26128 9464 26192
rect 9337 26112 9464 26128
rect 9337 26048 9384 26112
rect 9448 26048 9464 26112
rect 9337 26032 9464 26048
rect 9337 25968 9384 26032
rect 9448 25968 9464 26032
rect 9337 25952 9464 25968
rect 9337 25888 9384 25952
rect 9448 25888 9464 25952
rect 9337 25872 9464 25888
rect 9337 25808 9384 25872
rect 9448 25808 9464 25872
rect 9337 25792 9464 25808
rect 9337 25728 9384 25792
rect 9448 25728 9464 25792
rect 9337 25712 9464 25728
rect 9337 25648 9384 25712
rect 9448 25648 9464 25712
rect 9337 25632 9464 25648
rect 9337 25568 9384 25632
rect 9448 25568 9464 25632
rect 9337 25552 9464 25568
rect 9337 25488 9384 25552
rect 9448 25488 9464 25552
rect 9337 25472 9464 25488
rect 9337 25408 9384 25472
rect 9448 25408 9464 25472
rect 9337 25392 9464 25408
rect 9337 25328 9384 25392
rect 9448 25328 9464 25392
rect 9337 25312 9464 25328
rect 9337 25248 9384 25312
rect 9448 25248 9464 25312
rect 9337 25232 9464 25248
rect 9337 25168 9384 25232
rect 9448 25168 9464 25232
rect 9337 25152 9464 25168
rect 9337 25088 9384 25152
rect 9448 25088 9464 25152
rect 9337 25072 9464 25088
rect 9337 25008 9384 25072
rect 9448 25008 9464 25072
rect 9337 24992 9464 25008
rect 9337 24928 9384 24992
rect 9448 24928 9464 24992
rect 9337 24912 9464 24928
rect 9337 24848 9384 24912
rect 9448 24848 9464 24912
rect 9337 24832 9464 24848
rect 9337 24768 9384 24832
rect 9448 24768 9464 24832
rect 9337 24752 9464 24768
rect 9337 24688 9384 24752
rect 9448 24688 9464 24752
rect 9337 24672 9464 24688
rect 9337 24608 9384 24672
rect 9448 24608 9464 24672
rect 9337 24592 9464 24608
rect 9337 24528 9384 24592
rect 9448 24528 9464 24592
rect 9337 24512 9464 24528
rect 9337 24448 9384 24512
rect 9448 24448 9464 24512
rect 9337 24432 9464 24448
rect 9337 24368 9384 24432
rect 9448 24368 9464 24432
rect 9337 24352 9464 24368
rect 9337 24288 9384 24352
rect 9448 24288 9464 24352
rect 9337 24272 9464 24288
rect 9337 24208 9384 24272
rect 9448 24208 9464 24272
rect 9337 24192 9464 24208
rect 9337 24128 9384 24192
rect 9448 24128 9464 24192
rect 9337 24112 9464 24128
rect 9337 24048 9384 24112
rect 9448 24048 9464 24112
rect 9337 24032 9464 24048
rect 9337 23968 9384 24032
rect 9448 23968 9464 24032
rect 9337 23952 9464 23968
rect 9337 23888 9384 23952
rect 9448 23888 9464 23952
rect 9337 23872 9464 23888
rect 9337 23808 9384 23872
rect 9448 23808 9464 23872
rect 9337 23792 9464 23808
rect 9337 23728 9384 23792
rect 9448 23728 9464 23792
rect 9337 23712 9464 23728
rect 9337 23648 9384 23712
rect 9448 23648 9464 23712
rect 9337 23632 9464 23648
rect 9337 23568 9384 23632
rect 9448 23568 9464 23632
rect 9337 23552 9464 23568
rect 9337 23488 9384 23552
rect 9448 23488 9464 23552
rect 9337 23472 9464 23488
rect 9337 23408 9384 23472
rect 9448 23408 9464 23472
rect 9337 23392 9464 23408
rect 9337 23328 9384 23392
rect 9448 23328 9464 23392
rect 9337 23312 9464 23328
rect 9337 23248 9384 23312
rect 9448 23248 9464 23312
rect 9337 23232 9464 23248
rect 9337 23168 9384 23232
rect 9448 23168 9464 23232
rect 9337 23152 9464 23168
rect 9337 23088 9384 23152
rect 9448 23088 9464 23152
rect 9337 23072 9464 23088
rect 9337 23008 9384 23072
rect 9448 23008 9464 23072
rect 9337 22992 9464 23008
rect 9337 22928 9384 22992
rect 9448 22928 9464 22992
rect 9337 22912 9464 22928
rect 9337 22848 9384 22912
rect 9448 22848 9464 22912
rect 9337 22832 9464 22848
rect 9337 22768 9384 22832
rect 9448 22768 9464 22832
rect 9337 22752 9464 22768
rect 9337 22688 9384 22752
rect 9448 22688 9464 22752
rect 9337 22672 9464 22688
rect 9337 22608 9384 22672
rect 9448 22608 9464 22672
rect 9337 22592 9464 22608
rect 9337 22528 9384 22592
rect 9448 22528 9464 22592
rect 9337 22512 9464 22528
rect 9337 22448 9384 22512
rect 9448 22448 9464 22512
rect 9337 22432 9464 22448
rect 9337 22368 9384 22432
rect 9448 22368 9464 22432
rect 9337 22352 9464 22368
rect 9337 22288 9384 22352
rect 9448 22288 9464 22352
rect 9337 22272 9464 22288
rect 3018 22192 3145 22208
rect 3018 22128 3065 22192
rect 3129 22128 3145 22192
rect 3018 22112 3145 22128
rect 3018 21988 3122 22112
rect 3018 21972 3145 21988
rect 3018 21908 3065 21972
rect 3129 21908 3145 21972
rect 3018 21892 3145 21908
rect -3301 21812 -3174 21828
rect -3301 21748 -3254 21812
rect -3190 21748 -3174 21812
rect -3301 21732 -3174 21748
rect -3301 21668 -3254 21732
rect -3190 21668 -3174 21732
rect -3301 21652 -3174 21668
rect -3301 21588 -3254 21652
rect -3190 21588 -3174 21652
rect -3301 21572 -3174 21588
rect -3301 21508 -3254 21572
rect -3190 21508 -3174 21572
rect -3301 21492 -3174 21508
rect -3301 21428 -3254 21492
rect -3190 21428 -3174 21492
rect -3301 21412 -3174 21428
rect -3301 21348 -3254 21412
rect -3190 21348 -3174 21412
rect -3301 21332 -3174 21348
rect -3301 21268 -3254 21332
rect -3190 21268 -3174 21332
rect -3301 21252 -3174 21268
rect -3301 21188 -3254 21252
rect -3190 21188 -3174 21252
rect -3301 21172 -3174 21188
rect -3301 21108 -3254 21172
rect -3190 21108 -3174 21172
rect -3301 21092 -3174 21108
rect -3301 21028 -3254 21092
rect -3190 21028 -3174 21092
rect -3301 21012 -3174 21028
rect -3301 20948 -3254 21012
rect -3190 20948 -3174 21012
rect -3301 20932 -3174 20948
rect -3301 20868 -3254 20932
rect -3190 20868 -3174 20932
rect -3301 20852 -3174 20868
rect -3301 20788 -3254 20852
rect -3190 20788 -3174 20852
rect -3301 20772 -3174 20788
rect -3301 20708 -3254 20772
rect -3190 20708 -3174 20772
rect -3301 20692 -3174 20708
rect -3301 20628 -3254 20692
rect -3190 20628 -3174 20692
rect -3301 20612 -3174 20628
rect -3301 20548 -3254 20612
rect -3190 20548 -3174 20612
rect -3301 20532 -3174 20548
rect -3301 20468 -3254 20532
rect -3190 20468 -3174 20532
rect -3301 20452 -3174 20468
rect -3301 20388 -3254 20452
rect -3190 20388 -3174 20452
rect -3301 20372 -3174 20388
rect -3301 20308 -3254 20372
rect -3190 20308 -3174 20372
rect -3301 20292 -3174 20308
rect -3301 20228 -3254 20292
rect -3190 20228 -3174 20292
rect -3301 20212 -3174 20228
rect -3301 20148 -3254 20212
rect -3190 20148 -3174 20212
rect -3301 20132 -3174 20148
rect -3301 20068 -3254 20132
rect -3190 20068 -3174 20132
rect -3301 20052 -3174 20068
rect -3301 19988 -3254 20052
rect -3190 19988 -3174 20052
rect -3301 19972 -3174 19988
rect -3301 19908 -3254 19972
rect -3190 19908 -3174 19972
rect -3301 19892 -3174 19908
rect -3301 19828 -3254 19892
rect -3190 19828 -3174 19892
rect -3301 19812 -3174 19828
rect -3301 19748 -3254 19812
rect -3190 19748 -3174 19812
rect -3301 19732 -3174 19748
rect -3301 19668 -3254 19732
rect -3190 19668 -3174 19732
rect -3301 19652 -3174 19668
rect -3301 19588 -3254 19652
rect -3190 19588 -3174 19652
rect -3301 19572 -3174 19588
rect -3301 19508 -3254 19572
rect -3190 19508 -3174 19572
rect -3301 19492 -3174 19508
rect -3301 19428 -3254 19492
rect -3190 19428 -3174 19492
rect -3301 19412 -3174 19428
rect -3301 19348 -3254 19412
rect -3190 19348 -3174 19412
rect -3301 19332 -3174 19348
rect -3301 19268 -3254 19332
rect -3190 19268 -3174 19332
rect -3301 19252 -3174 19268
rect -3301 19188 -3254 19252
rect -3190 19188 -3174 19252
rect -3301 19172 -3174 19188
rect -3301 19108 -3254 19172
rect -3190 19108 -3174 19172
rect -3301 19092 -3174 19108
rect -3301 19028 -3254 19092
rect -3190 19028 -3174 19092
rect -3301 19012 -3174 19028
rect -3301 18948 -3254 19012
rect -3190 18948 -3174 19012
rect -3301 18932 -3174 18948
rect -3301 18868 -3254 18932
rect -3190 18868 -3174 18932
rect -3301 18852 -3174 18868
rect -3301 18788 -3254 18852
rect -3190 18788 -3174 18852
rect -3301 18772 -3174 18788
rect -3301 18708 -3254 18772
rect -3190 18708 -3174 18772
rect -3301 18692 -3174 18708
rect -3301 18628 -3254 18692
rect -3190 18628 -3174 18692
rect -3301 18612 -3174 18628
rect -3301 18548 -3254 18612
rect -3190 18548 -3174 18612
rect -3301 18532 -3174 18548
rect -3301 18468 -3254 18532
rect -3190 18468 -3174 18532
rect -3301 18452 -3174 18468
rect -3301 18388 -3254 18452
rect -3190 18388 -3174 18452
rect -3301 18372 -3174 18388
rect -3301 18308 -3254 18372
rect -3190 18308 -3174 18372
rect -3301 18292 -3174 18308
rect -3301 18228 -3254 18292
rect -3190 18228 -3174 18292
rect -3301 18212 -3174 18228
rect -3301 18148 -3254 18212
rect -3190 18148 -3174 18212
rect -3301 18132 -3174 18148
rect -3301 18068 -3254 18132
rect -3190 18068 -3174 18132
rect -3301 18052 -3174 18068
rect -3301 17988 -3254 18052
rect -3190 17988 -3174 18052
rect -3301 17972 -3174 17988
rect -3301 17908 -3254 17972
rect -3190 17908 -3174 17972
rect -3301 17892 -3174 17908
rect -3301 17828 -3254 17892
rect -3190 17828 -3174 17892
rect -3301 17812 -3174 17828
rect -3301 17748 -3254 17812
rect -3190 17748 -3174 17812
rect -3301 17732 -3174 17748
rect -3301 17668 -3254 17732
rect -3190 17668 -3174 17732
rect -3301 17652 -3174 17668
rect -3301 17588 -3254 17652
rect -3190 17588 -3174 17652
rect -3301 17572 -3174 17588
rect -3301 17508 -3254 17572
rect -3190 17508 -3174 17572
rect -3301 17492 -3174 17508
rect -3301 17428 -3254 17492
rect -3190 17428 -3174 17492
rect -3301 17412 -3174 17428
rect -3301 17348 -3254 17412
rect -3190 17348 -3174 17412
rect -3301 17332 -3174 17348
rect -3301 17268 -3254 17332
rect -3190 17268 -3174 17332
rect -3301 17252 -3174 17268
rect -3301 17188 -3254 17252
rect -3190 17188 -3174 17252
rect -3301 17172 -3174 17188
rect -3301 17108 -3254 17172
rect -3190 17108 -3174 17172
rect -3301 17092 -3174 17108
rect -3301 17028 -3254 17092
rect -3190 17028 -3174 17092
rect -3301 17012 -3174 17028
rect -3301 16948 -3254 17012
rect -3190 16948 -3174 17012
rect -3301 16932 -3174 16948
rect -3301 16868 -3254 16932
rect -3190 16868 -3174 16932
rect -3301 16852 -3174 16868
rect -3301 16788 -3254 16852
rect -3190 16788 -3174 16852
rect -3301 16772 -3174 16788
rect -3301 16708 -3254 16772
rect -3190 16708 -3174 16772
rect -3301 16692 -3174 16708
rect -3301 16628 -3254 16692
rect -3190 16628 -3174 16692
rect -3301 16612 -3174 16628
rect -3301 16548 -3254 16612
rect -3190 16548 -3174 16612
rect -3301 16532 -3174 16548
rect -3301 16468 -3254 16532
rect -3190 16468 -3174 16532
rect -3301 16452 -3174 16468
rect -3301 16388 -3254 16452
rect -3190 16388 -3174 16452
rect -3301 16372 -3174 16388
rect -3301 16308 -3254 16372
rect -3190 16308 -3174 16372
rect -3301 16292 -3174 16308
rect -3301 16228 -3254 16292
rect -3190 16228 -3174 16292
rect -3301 16212 -3174 16228
rect -3301 16148 -3254 16212
rect -3190 16148 -3174 16212
rect -3301 16132 -3174 16148
rect -3301 16068 -3254 16132
rect -3190 16068 -3174 16132
rect -3301 16052 -3174 16068
rect -3301 15988 -3254 16052
rect -3190 15988 -3174 16052
rect -3301 15972 -3174 15988
rect -9620 15892 -9493 15908
rect -9620 15828 -9573 15892
rect -9509 15828 -9493 15892
rect -9620 15812 -9493 15828
rect -9620 15688 -9516 15812
rect -9620 15672 -9493 15688
rect -9620 15608 -9573 15672
rect -9509 15608 -9493 15672
rect -9620 15592 -9493 15608
rect -15939 15512 -15812 15528
rect -15939 15448 -15892 15512
rect -15828 15448 -15812 15512
rect -15939 15432 -15812 15448
rect -15939 15368 -15892 15432
rect -15828 15368 -15812 15432
rect -15939 15352 -15812 15368
rect -15939 15288 -15892 15352
rect -15828 15288 -15812 15352
rect -15939 15272 -15812 15288
rect -15939 15208 -15892 15272
rect -15828 15208 -15812 15272
rect -15939 15192 -15812 15208
rect -15939 15128 -15892 15192
rect -15828 15128 -15812 15192
rect -15939 15112 -15812 15128
rect -15939 15048 -15892 15112
rect -15828 15048 -15812 15112
rect -15939 15032 -15812 15048
rect -15939 14968 -15892 15032
rect -15828 14968 -15812 15032
rect -15939 14952 -15812 14968
rect -15939 14888 -15892 14952
rect -15828 14888 -15812 14952
rect -15939 14872 -15812 14888
rect -15939 14808 -15892 14872
rect -15828 14808 -15812 14872
rect -15939 14792 -15812 14808
rect -15939 14728 -15892 14792
rect -15828 14728 -15812 14792
rect -15939 14712 -15812 14728
rect -15939 14648 -15892 14712
rect -15828 14648 -15812 14712
rect -15939 14632 -15812 14648
rect -15939 14568 -15892 14632
rect -15828 14568 -15812 14632
rect -15939 14552 -15812 14568
rect -15939 14488 -15892 14552
rect -15828 14488 -15812 14552
rect -15939 14472 -15812 14488
rect -15939 14408 -15892 14472
rect -15828 14408 -15812 14472
rect -15939 14392 -15812 14408
rect -15939 14328 -15892 14392
rect -15828 14328 -15812 14392
rect -15939 14312 -15812 14328
rect -15939 14248 -15892 14312
rect -15828 14248 -15812 14312
rect -15939 14232 -15812 14248
rect -15939 14168 -15892 14232
rect -15828 14168 -15812 14232
rect -15939 14152 -15812 14168
rect -15939 14088 -15892 14152
rect -15828 14088 -15812 14152
rect -15939 14072 -15812 14088
rect -15939 14008 -15892 14072
rect -15828 14008 -15812 14072
rect -15939 13992 -15812 14008
rect -15939 13928 -15892 13992
rect -15828 13928 -15812 13992
rect -15939 13912 -15812 13928
rect -15939 13848 -15892 13912
rect -15828 13848 -15812 13912
rect -15939 13832 -15812 13848
rect -15939 13768 -15892 13832
rect -15828 13768 -15812 13832
rect -15939 13752 -15812 13768
rect -15939 13688 -15892 13752
rect -15828 13688 -15812 13752
rect -15939 13672 -15812 13688
rect -15939 13608 -15892 13672
rect -15828 13608 -15812 13672
rect -15939 13592 -15812 13608
rect -15939 13528 -15892 13592
rect -15828 13528 -15812 13592
rect -15939 13512 -15812 13528
rect -15939 13448 -15892 13512
rect -15828 13448 -15812 13512
rect -15939 13432 -15812 13448
rect -15939 13368 -15892 13432
rect -15828 13368 -15812 13432
rect -15939 13352 -15812 13368
rect -15939 13288 -15892 13352
rect -15828 13288 -15812 13352
rect -15939 13272 -15812 13288
rect -15939 13208 -15892 13272
rect -15828 13208 -15812 13272
rect -15939 13192 -15812 13208
rect -15939 13128 -15892 13192
rect -15828 13128 -15812 13192
rect -15939 13112 -15812 13128
rect -15939 13048 -15892 13112
rect -15828 13048 -15812 13112
rect -15939 13032 -15812 13048
rect -15939 12968 -15892 13032
rect -15828 12968 -15812 13032
rect -15939 12952 -15812 12968
rect -15939 12888 -15892 12952
rect -15828 12888 -15812 12952
rect -15939 12872 -15812 12888
rect -15939 12808 -15892 12872
rect -15828 12808 -15812 12872
rect -15939 12792 -15812 12808
rect -15939 12728 -15892 12792
rect -15828 12728 -15812 12792
rect -15939 12712 -15812 12728
rect -15939 12648 -15892 12712
rect -15828 12648 -15812 12712
rect -15939 12632 -15812 12648
rect -15939 12568 -15892 12632
rect -15828 12568 -15812 12632
rect -15939 12552 -15812 12568
rect -15939 12488 -15892 12552
rect -15828 12488 -15812 12552
rect -15939 12472 -15812 12488
rect -15939 12408 -15892 12472
rect -15828 12408 -15812 12472
rect -15939 12392 -15812 12408
rect -15939 12328 -15892 12392
rect -15828 12328 -15812 12392
rect -15939 12312 -15812 12328
rect -15939 12248 -15892 12312
rect -15828 12248 -15812 12312
rect -15939 12232 -15812 12248
rect -15939 12168 -15892 12232
rect -15828 12168 -15812 12232
rect -15939 12152 -15812 12168
rect -15939 12088 -15892 12152
rect -15828 12088 -15812 12152
rect -15939 12072 -15812 12088
rect -15939 12008 -15892 12072
rect -15828 12008 -15812 12072
rect -15939 11992 -15812 12008
rect -15939 11928 -15892 11992
rect -15828 11928 -15812 11992
rect -15939 11912 -15812 11928
rect -15939 11848 -15892 11912
rect -15828 11848 -15812 11912
rect -15939 11832 -15812 11848
rect -15939 11768 -15892 11832
rect -15828 11768 -15812 11832
rect -15939 11752 -15812 11768
rect -15939 11688 -15892 11752
rect -15828 11688 -15812 11752
rect -15939 11672 -15812 11688
rect -15939 11608 -15892 11672
rect -15828 11608 -15812 11672
rect -15939 11592 -15812 11608
rect -15939 11528 -15892 11592
rect -15828 11528 -15812 11592
rect -15939 11512 -15812 11528
rect -15939 11448 -15892 11512
rect -15828 11448 -15812 11512
rect -15939 11432 -15812 11448
rect -15939 11368 -15892 11432
rect -15828 11368 -15812 11432
rect -15939 11352 -15812 11368
rect -15939 11288 -15892 11352
rect -15828 11288 -15812 11352
rect -15939 11272 -15812 11288
rect -15939 11208 -15892 11272
rect -15828 11208 -15812 11272
rect -15939 11192 -15812 11208
rect -15939 11128 -15892 11192
rect -15828 11128 -15812 11192
rect -15939 11112 -15812 11128
rect -15939 11048 -15892 11112
rect -15828 11048 -15812 11112
rect -15939 11032 -15812 11048
rect -15939 10968 -15892 11032
rect -15828 10968 -15812 11032
rect -15939 10952 -15812 10968
rect -15939 10888 -15892 10952
rect -15828 10888 -15812 10952
rect -15939 10872 -15812 10888
rect -15939 10808 -15892 10872
rect -15828 10808 -15812 10872
rect -15939 10792 -15812 10808
rect -15939 10728 -15892 10792
rect -15828 10728 -15812 10792
rect -15939 10712 -15812 10728
rect -15939 10648 -15892 10712
rect -15828 10648 -15812 10712
rect -15939 10632 -15812 10648
rect -15939 10568 -15892 10632
rect -15828 10568 -15812 10632
rect -15939 10552 -15812 10568
rect -15939 10488 -15892 10552
rect -15828 10488 -15812 10552
rect -15939 10472 -15812 10488
rect -15939 10408 -15892 10472
rect -15828 10408 -15812 10472
rect -15939 10392 -15812 10408
rect -15939 10328 -15892 10392
rect -15828 10328 -15812 10392
rect -15939 10312 -15812 10328
rect -15939 10248 -15892 10312
rect -15828 10248 -15812 10312
rect -15939 10232 -15812 10248
rect -15939 10168 -15892 10232
rect -15828 10168 -15812 10232
rect -15939 10152 -15812 10168
rect -15939 10088 -15892 10152
rect -15828 10088 -15812 10152
rect -15939 10072 -15812 10088
rect -15939 10008 -15892 10072
rect -15828 10008 -15812 10072
rect -15939 9992 -15812 10008
rect -15939 9928 -15892 9992
rect -15828 9928 -15812 9992
rect -15939 9912 -15812 9928
rect -15939 9848 -15892 9912
rect -15828 9848 -15812 9912
rect -15939 9832 -15812 9848
rect -15939 9768 -15892 9832
rect -15828 9768 -15812 9832
rect -15939 9752 -15812 9768
rect -15939 9688 -15892 9752
rect -15828 9688 -15812 9752
rect -15939 9672 -15812 9688
rect -22258 9592 -22131 9608
rect -22258 9528 -22211 9592
rect -22147 9528 -22131 9592
rect -22258 9512 -22131 9528
rect -22258 9388 -22154 9512
rect -22258 9372 -22131 9388
rect -22258 9308 -22211 9372
rect -22147 9308 -22131 9372
rect -22258 9292 -22131 9308
rect -28577 9212 -28450 9228
rect -28577 9148 -28530 9212
rect -28466 9148 -28450 9212
rect -28577 9132 -28450 9148
rect -28577 9068 -28530 9132
rect -28466 9068 -28450 9132
rect -28577 9052 -28450 9068
rect -28577 8988 -28530 9052
rect -28466 8988 -28450 9052
rect -28577 8972 -28450 8988
rect -28577 8908 -28530 8972
rect -28466 8908 -28450 8972
rect -28577 8892 -28450 8908
rect -28577 8828 -28530 8892
rect -28466 8828 -28450 8892
rect -28577 8812 -28450 8828
rect -28577 8748 -28530 8812
rect -28466 8748 -28450 8812
rect -28577 8732 -28450 8748
rect -28577 8668 -28530 8732
rect -28466 8668 -28450 8732
rect -28577 8652 -28450 8668
rect -28577 8588 -28530 8652
rect -28466 8588 -28450 8652
rect -28577 8572 -28450 8588
rect -28577 8508 -28530 8572
rect -28466 8508 -28450 8572
rect -28577 8492 -28450 8508
rect -28577 8428 -28530 8492
rect -28466 8428 -28450 8492
rect -28577 8412 -28450 8428
rect -28577 8348 -28530 8412
rect -28466 8348 -28450 8412
rect -28577 8332 -28450 8348
rect -28577 8268 -28530 8332
rect -28466 8268 -28450 8332
rect -28577 8252 -28450 8268
rect -28577 8188 -28530 8252
rect -28466 8188 -28450 8252
rect -28577 8172 -28450 8188
rect -28577 8108 -28530 8172
rect -28466 8108 -28450 8172
rect -28577 8092 -28450 8108
rect -28577 8028 -28530 8092
rect -28466 8028 -28450 8092
rect -28577 8012 -28450 8028
rect -28577 7948 -28530 8012
rect -28466 7948 -28450 8012
rect -28577 7932 -28450 7948
rect -28577 7868 -28530 7932
rect -28466 7868 -28450 7932
rect -28577 7852 -28450 7868
rect -28577 7788 -28530 7852
rect -28466 7788 -28450 7852
rect -28577 7772 -28450 7788
rect -28577 7708 -28530 7772
rect -28466 7708 -28450 7772
rect -28577 7692 -28450 7708
rect -28577 7628 -28530 7692
rect -28466 7628 -28450 7692
rect -28577 7612 -28450 7628
rect -28577 7548 -28530 7612
rect -28466 7548 -28450 7612
rect -28577 7532 -28450 7548
rect -28577 7468 -28530 7532
rect -28466 7468 -28450 7532
rect -28577 7452 -28450 7468
rect -28577 7388 -28530 7452
rect -28466 7388 -28450 7452
rect -28577 7372 -28450 7388
rect -28577 7308 -28530 7372
rect -28466 7308 -28450 7372
rect -28577 7292 -28450 7308
rect -28577 7228 -28530 7292
rect -28466 7228 -28450 7292
rect -28577 7212 -28450 7228
rect -28577 7148 -28530 7212
rect -28466 7148 -28450 7212
rect -28577 7132 -28450 7148
rect -28577 7068 -28530 7132
rect -28466 7068 -28450 7132
rect -28577 7052 -28450 7068
rect -28577 6988 -28530 7052
rect -28466 6988 -28450 7052
rect -28577 6972 -28450 6988
rect -28577 6908 -28530 6972
rect -28466 6908 -28450 6972
rect -28577 6892 -28450 6908
rect -28577 6828 -28530 6892
rect -28466 6828 -28450 6892
rect -28577 6812 -28450 6828
rect -28577 6748 -28530 6812
rect -28466 6748 -28450 6812
rect -28577 6732 -28450 6748
rect -28577 6668 -28530 6732
rect -28466 6668 -28450 6732
rect -28577 6652 -28450 6668
rect -28577 6588 -28530 6652
rect -28466 6588 -28450 6652
rect -28577 6572 -28450 6588
rect -28577 6508 -28530 6572
rect -28466 6508 -28450 6572
rect -28577 6492 -28450 6508
rect -28577 6428 -28530 6492
rect -28466 6428 -28450 6492
rect -28577 6412 -28450 6428
rect -28577 6348 -28530 6412
rect -28466 6348 -28450 6412
rect -28577 6332 -28450 6348
rect -28577 6268 -28530 6332
rect -28466 6268 -28450 6332
rect -28577 6252 -28450 6268
rect -28577 6188 -28530 6252
rect -28466 6188 -28450 6252
rect -28577 6172 -28450 6188
rect -28577 6108 -28530 6172
rect -28466 6108 -28450 6172
rect -28577 6092 -28450 6108
rect -28577 6028 -28530 6092
rect -28466 6028 -28450 6092
rect -28577 6012 -28450 6028
rect -28577 5948 -28530 6012
rect -28466 5948 -28450 6012
rect -28577 5932 -28450 5948
rect -28577 5868 -28530 5932
rect -28466 5868 -28450 5932
rect -28577 5852 -28450 5868
rect -28577 5788 -28530 5852
rect -28466 5788 -28450 5852
rect -28577 5772 -28450 5788
rect -28577 5708 -28530 5772
rect -28466 5708 -28450 5772
rect -28577 5692 -28450 5708
rect -28577 5628 -28530 5692
rect -28466 5628 -28450 5692
rect -28577 5612 -28450 5628
rect -28577 5548 -28530 5612
rect -28466 5548 -28450 5612
rect -28577 5532 -28450 5548
rect -28577 5468 -28530 5532
rect -28466 5468 -28450 5532
rect -28577 5452 -28450 5468
rect -28577 5388 -28530 5452
rect -28466 5388 -28450 5452
rect -28577 5372 -28450 5388
rect -28577 5308 -28530 5372
rect -28466 5308 -28450 5372
rect -28577 5292 -28450 5308
rect -28577 5228 -28530 5292
rect -28466 5228 -28450 5292
rect -28577 5212 -28450 5228
rect -28577 5148 -28530 5212
rect -28466 5148 -28450 5212
rect -28577 5132 -28450 5148
rect -28577 5068 -28530 5132
rect -28466 5068 -28450 5132
rect -28577 5052 -28450 5068
rect -28577 4988 -28530 5052
rect -28466 4988 -28450 5052
rect -28577 4972 -28450 4988
rect -28577 4908 -28530 4972
rect -28466 4908 -28450 4972
rect -28577 4892 -28450 4908
rect -28577 4828 -28530 4892
rect -28466 4828 -28450 4892
rect -28577 4812 -28450 4828
rect -28577 4748 -28530 4812
rect -28466 4748 -28450 4812
rect -28577 4732 -28450 4748
rect -28577 4668 -28530 4732
rect -28466 4668 -28450 4732
rect -28577 4652 -28450 4668
rect -28577 4588 -28530 4652
rect -28466 4588 -28450 4652
rect -28577 4572 -28450 4588
rect -28577 4508 -28530 4572
rect -28466 4508 -28450 4572
rect -28577 4492 -28450 4508
rect -28577 4428 -28530 4492
rect -28466 4428 -28450 4492
rect -28577 4412 -28450 4428
rect -28577 4348 -28530 4412
rect -28466 4348 -28450 4412
rect -28577 4332 -28450 4348
rect -28577 4268 -28530 4332
rect -28466 4268 -28450 4332
rect -28577 4252 -28450 4268
rect -28577 4188 -28530 4252
rect -28466 4188 -28450 4252
rect -28577 4172 -28450 4188
rect -28577 4108 -28530 4172
rect -28466 4108 -28450 4172
rect -28577 4092 -28450 4108
rect -28577 4028 -28530 4092
rect -28466 4028 -28450 4092
rect -28577 4012 -28450 4028
rect -28577 3948 -28530 4012
rect -28466 3948 -28450 4012
rect -28577 3932 -28450 3948
rect -28577 3868 -28530 3932
rect -28466 3868 -28450 3932
rect -28577 3852 -28450 3868
rect -28577 3788 -28530 3852
rect -28466 3788 -28450 3852
rect -28577 3772 -28450 3788
rect -28577 3708 -28530 3772
rect -28466 3708 -28450 3772
rect -28577 3692 -28450 3708
rect -28577 3628 -28530 3692
rect -28466 3628 -28450 3692
rect -28577 3612 -28450 3628
rect -28577 3548 -28530 3612
rect -28466 3548 -28450 3612
rect -28577 3532 -28450 3548
rect -28577 3468 -28530 3532
rect -28466 3468 -28450 3532
rect -28577 3452 -28450 3468
rect -28577 3388 -28530 3452
rect -28466 3388 -28450 3452
rect -28577 3372 -28450 3388
rect -34896 3292 -34769 3308
rect -34896 3228 -34849 3292
rect -34785 3228 -34769 3292
rect -34896 3212 -34769 3228
rect -34896 3088 -34792 3212
rect -34896 3072 -34769 3088
rect -34896 3008 -34849 3072
rect -34785 3008 -34769 3072
rect -34896 2992 -34769 3008
rect -41215 2912 -41088 2928
rect -41215 2848 -41168 2912
rect -41104 2848 -41088 2912
rect -41215 2832 -41088 2848
rect -41215 2768 -41168 2832
rect -41104 2768 -41088 2832
rect -41215 2752 -41088 2768
rect -41215 2688 -41168 2752
rect -41104 2688 -41088 2752
rect -41215 2672 -41088 2688
rect -41215 2608 -41168 2672
rect -41104 2608 -41088 2672
rect -41215 2592 -41088 2608
rect -41215 2528 -41168 2592
rect -41104 2528 -41088 2592
rect -41215 2512 -41088 2528
rect -41215 2448 -41168 2512
rect -41104 2448 -41088 2512
rect -41215 2432 -41088 2448
rect -41215 2368 -41168 2432
rect -41104 2368 -41088 2432
rect -41215 2352 -41088 2368
rect -41215 2288 -41168 2352
rect -41104 2288 -41088 2352
rect -41215 2272 -41088 2288
rect -41215 2208 -41168 2272
rect -41104 2208 -41088 2272
rect -41215 2192 -41088 2208
rect -41215 2128 -41168 2192
rect -41104 2128 -41088 2192
rect -41215 2112 -41088 2128
rect -41215 2048 -41168 2112
rect -41104 2048 -41088 2112
rect -41215 2032 -41088 2048
rect -41215 1968 -41168 2032
rect -41104 1968 -41088 2032
rect -41215 1952 -41088 1968
rect -41215 1888 -41168 1952
rect -41104 1888 -41088 1952
rect -41215 1872 -41088 1888
rect -41215 1808 -41168 1872
rect -41104 1808 -41088 1872
rect -41215 1792 -41088 1808
rect -41215 1728 -41168 1792
rect -41104 1728 -41088 1792
rect -41215 1712 -41088 1728
rect -41215 1648 -41168 1712
rect -41104 1648 -41088 1712
rect -41215 1632 -41088 1648
rect -41215 1568 -41168 1632
rect -41104 1568 -41088 1632
rect -41215 1552 -41088 1568
rect -41215 1488 -41168 1552
rect -41104 1488 -41088 1552
rect -41215 1472 -41088 1488
rect -41215 1408 -41168 1472
rect -41104 1408 -41088 1472
rect -41215 1392 -41088 1408
rect -41215 1328 -41168 1392
rect -41104 1328 -41088 1392
rect -41215 1312 -41088 1328
rect -41215 1248 -41168 1312
rect -41104 1248 -41088 1312
rect -41215 1232 -41088 1248
rect -41215 1168 -41168 1232
rect -41104 1168 -41088 1232
rect -41215 1152 -41088 1168
rect -41215 1088 -41168 1152
rect -41104 1088 -41088 1152
rect -41215 1072 -41088 1088
rect -41215 1008 -41168 1072
rect -41104 1008 -41088 1072
rect -41215 992 -41088 1008
rect -41215 928 -41168 992
rect -41104 928 -41088 992
rect -41215 912 -41088 928
rect -41215 848 -41168 912
rect -41104 848 -41088 912
rect -41215 832 -41088 848
rect -41215 768 -41168 832
rect -41104 768 -41088 832
rect -41215 752 -41088 768
rect -41215 688 -41168 752
rect -41104 688 -41088 752
rect -41215 672 -41088 688
rect -41215 608 -41168 672
rect -41104 608 -41088 672
rect -41215 592 -41088 608
rect -41215 528 -41168 592
rect -41104 528 -41088 592
rect -41215 512 -41088 528
rect -41215 448 -41168 512
rect -41104 448 -41088 512
rect -41215 432 -41088 448
rect -41215 368 -41168 432
rect -41104 368 -41088 432
rect -41215 352 -41088 368
rect -41215 288 -41168 352
rect -41104 288 -41088 352
rect -41215 272 -41088 288
rect -41215 208 -41168 272
rect -41104 208 -41088 272
rect -41215 192 -41088 208
rect -41215 128 -41168 192
rect -41104 128 -41088 192
rect -41215 112 -41088 128
rect -41215 48 -41168 112
rect -41104 48 -41088 112
rect -41215 32 -41088 48
rect -41215 -32 -41168 32
rect -41104 -32 -41088 32
rect -41215 -48 -41088 -32
rect -41215 -112 -41168 -48
rect -41104 -112 -41088 -48
rect -41215 -128 -41088 -112
rect -41215 -192 -41168 -128
rect -41104 -192 -41088 -128
rect -41215 -208 -41088 -192
rect -41215 -272 -41168 -208
rect -41104 -272 -41088 -208
rect -41215 -288 -41088 -272
rect -41215 -352 -41168 -288
rect -41104 -352 -41088 -288
rect -41215 -368 -41088 -352
rect -41215 -432 -41168 -368
rect -41104 -432 -41088 -368
rect -41215 -448 -41088 -432
rect -41215 -512 -41168 -448
rect -41104 -512 -41088 -448
rect -41215 -528 -41088 -512
rect -41215 -592 -41168 -528
rect -41104 -592 -41088 -528
rect -41215 -608 -41088 -592
rect -41215 -672 -41168 -608
rect -41104 -672 -41088 -608
rect -41215 -688 -41088 -672
rect -41215 -752 -41168 -688
rect -41104 -752 -41088 -688
rect -41215 -768 -41088 -752
rect -41215 -832 -41168 -768
rect -41104 -832 -41088 -768
rect -41215 -848 -41088 -832
rect -41215 -912 -41168 -848
rect -41104 -912 -41088 -848
rect -41215 -928 -41088 -912
rect -41215 -992 -41168 -928
rect -41104 -992 -41088 -928
rect -41215 -1008 -41088 -992
rect -41215 -1072 -41168 -1008
rect -41104 -1072 -41088 -1008
rect -41215 -1088 -41088 -1072
rect -41215 -1152 -41168 -1088
rect -41104 -1152 -41088 -1088
rect -41215 -1168 -41088 -1152
rect -41215 -1232 -41168 -1168
rect -41104 -1232 -41088 -1168
rect -41215 -1248 -41088 -1232
rect -41215 -1312 -41168 -1248
rect -41104 -1312 -41088 -1248
rect -41215 -1328 -41088 -1312
rect -41215 -1392 -41168 -1328
rect -41104 -1392 -41088 -1328
rect -41215 -1408 -41088 -1392
rect -41215 -1472 -41168 -1408
rect -41104 -1472 -41088 -1408
rect -41215 -1488 -41088 -1472
rect -41215 -1552 -41168 -1488
rect -41104 -1552 -41088 -1488
rect -41215 -1568 -41088 -1552
rect -41215 -1632 -41168 -1568
rect -41104 -1632 -41088 -1568
rect -41215 -1648 -41088 -1632
rect -41215 -1712 -41168 -1648
rect -41104 -1712 -41088 -1648
rect -41215 -1728 -41088 -1712
rect -41215 -1792 -41168 -1728
rect -41104 -1792 -41088 -1728
rect -41215 -1808 -41088 -1792
rect -41215 -1872 -41168 -1808
rect -41104 -1872 -41088 -1808
rect -41215 -1888 -41088 -1872
rect -41215 -1952 -41168 -1888
rect -41104 -1952 -41088 -1888
rect -41215 -1968 -41088 -1952
rect -41215 -2032 -41168 -1968
rect -41104 -2032 -41088 -1968
rect -41215 -2048 -41088 -2032
rect -41215 -2112 -41168 -2048
rect -41104 -2112 -41088 -2048
rect -41215 -2128 -41088 -2112
rect -41215 -2192 -41168 -2128
rect -41104 -2192 -41088 -2128
rect -41215 -2208 -41088 -2192
rect -41215 -2272 -41168 -2208
rect -41104 -2272 -41088 -2208
rect -41215 -2288 -41088 -2272
rect -41215 -2352 -41168 -2288
rect -41104 -2352 -41088 -2288
rect -41215 -2368 -41088 -2352
rect -41215 -2432 -41168 -2368
rect -41104 -2432 -41088 -2368
rect -41215 -2448 -41088 -2432
rect -41215 -2512 -41168 -2448
rect -41104 -2512 -41088 -2448
rect -41215 -2528 -41088 -2512
rect -41215 -2592 -41168 -2528
rect -41104 -2592 -41088 -2528
rect -41215 -2608 -41088 -2592
rect -41215 -2672 -41168 -2608
rect -41104 -2672 -41088 -2608
rect -41215 -2688 -41088 -2672
rect -41215 -2752 -41168 -2688
rect -41104 -2752 -41088 -2688
rect -41215 -2768 -41088 -2752
rect -41215 -2832 -41168 -2768
rect -41104 -2832 -41088 -2768
rect -41215 -2848 -41088 -2832
rect -41215 -2912 -41168 -2848
rect -41104 -2912 -41088 -2848
rect -41215 -2928 -41088 -2912
rect -44335 -3339 -44231 -2961
rect -41215 -2992 -41168 -2928
rect -41104 -2992 -41088 -2928
rect -40925 2952 -35003 2961
rect -40925 -2952 -40916 2952
rect -35012 -2952 -35003 2952
rect -40925 -2961 -35003 -2952
rect -34896 2928 -34849 2992
rect -34785 2928 -34769 2992
rect -31697 2961 -31593 3339
rect -28577 3308 -28530 3372
rect -28466 3308 -28450 3372
rect -28287 9252 -22365 9261
rect -28287 3348 -28278 9252
rect -22374 3348 -22365 9252
rect -28287 3339 -22365 3348
rect -22258 9228 -22211 9292
rect -22147 9228 -22131 9292
rect -19059 9261 -18955 9639
rect -15939 9608 -15892 9672
rect -15828 9608 -15812 9672
rect -15649 15552 -9727 15561
rect -15649 9648 -15640 15552
rect -9736 9648 -9727 15552
rect -15649 9639 -9727 9648
rect -9620 15528 -9573 15592
rect -9509 15528 -9493 15592
rect -6421 15561 -6317 15939
rect -3301 15908 -3254 15972
rect -3190 15908 -3174 15972
rect -3011 21852 2911 21861
rect -3011 15948 -3002 21852
rect 2902 15948 2911 21852
rect -3011 15939 2911 15948
rect 3018 21828 3065 21892
rect 3129 21828 3145 21892
rect 6217 21861 6321 22239
rect 9337 22208 9384 22272
rect 9448 22208 9464 22272
rect 9627 28152 15549 28161
rect 9627 22248 9636 28152
rect 15540 22248 15549 28152
rect 9627 22239 15549 22248
rect 15656 28128 15703 28192
rect 15767 28128 15783 28192
rect 18855 28161 18959 28539
rect 21975 28508 22022 28572
rect 22086 28508 22102 28572
rect 22265 34452 28187 34461
rect 22265 28548 22274 34452
rect 28178 28548 28187 34452
rect 22265 28539 28187 28548
rect 28294 34428 28341 34492
rect 28405 34428 28421 34492
rect 31493 34461 31597 34839
rect 34613 34808 34660 34872
rect 34724 34808 34740 34872
rect 34903 40752 40825 40761
rect 34903 34848 34912 40752
rect 40816 34848 40825 40752
rect 34903 34839 40825 34848
rect 40932 40728 40979 40792
rect 41043 40728 41059 40792
rect 44131 40761 44235 41139
rect 47251 41108 47298 41172
rect 47362 41108 47378 41172
rect 47251 41092 47378 41108
rect 47251 41028 47298 41092
rect 47362 41028 47378 41092
rect 47251 41012 47378 41028
rect 47251 40888 47355 41012
rect 47251 40872 47378 40888
rect 47251 40808 47298 40872
rect 47362 40808 47378 40872
rect 47251 40792 47378 40808
rect 40932 40712 41059 40728
rect 40932 40648 40979 40712
rect 41043 40648 41059 40712
rect 40932 40632 41059 40648
rect 40932 40568 40979 40632
rect 41043 40568 41059 40632
rect 40932 40552 41059 40568
rect 40932 40488 40979 40552
rect 41043 40488 41059 40552
rect 40932 40472 41059 40488
rect 40932 40408 40979 40472
rect 41043 40408 41059 40472
rect 40932 40392 41059 40408
rect 40932 40328 40979 40392
rect 41043 40328 41059 40392
rect 40932 40312 41059 40328
rect 40932 40248 40979 40312
rect 41043 40248 41059 40312
rect 40932 40232 41059 40248
rect 40932 40168 40979 40232
rect 41043 40168 41059 40232
rect 40932 40152 41059 40168
rect 40932 40088 40979 40152
rect 41043 40088 41059 40152
rect 40932 40072 41059 40088
rect 40932 40008 40979 40072
rect 41043 40008 41059 40072
rect 40932 39992 41059 40008
rect 40932 39928 40979 39992
rect 41043 39928 41059 39992
rect 40932 39912 41059 39928
rect 40932 39848 40979 39912
rect 41043 39848 41059 39912
rect 40932 39832 41059 39848
rect 40932 39768 40979 39832
rect 41043 39768 41059 39832
rect 40932 39752 41059 39768
rect 40932 39688 40979 39752
rect 41043 39688 41059 39752
rect 40932 39672 41059 39688
rect 40932 39608 40979 39672
rect 41043 39608 41059 39672
rect 40932 39592 41059 39608
rect 40932 39528 40979 39592
rect 41043 39528 41059 39592
rect 40932 39512 41059 39528
rect 40932 39448 40979 39512
rect 41043 39448 41059 39512
rect 40932 39432 41059 39448
rect 40932 39368 40979 39432
rect 41043 39368 41059 39432
rect 40932 39352 41059 39368
rect 40932 39288 40979 39352
rect 41043 39288 41059 39352
rect 40932 39272 41059 39288
rect 40932 39208 40979 39272
rect 41043 39208 41059 39272
rect 40932 39192 41059 39208
rect 40932 39128 40979 39192
rect 41043 39128 41059 39192
rect 40932 39112 41059 39128
rect 40932 39048 40979 39112
rect 41043 39048 41059 39112
rect 40932 39032 41059 39048
rect 40932 38968 40979 39032
rect 41043 38968 41059 39032
rect 40932 38952 41059 38968
rect 40932 38888 40979 38952
rect 41043 38888 41059 38952
rect 40932 38872 41059 38888
rect 40932 38808 40979 38872
rect 41043 38808 41059 38872
rect 40932 38792 41059 38808
rect 40932 38728 40979 38792
rect 41043 38728 41059 38792
rect 40932 38712 41059 38728
rect 40932 38648 40979 38712
rect 41043 38648 41059 38712
rect 40932 38632 41059 38648
rect 40932 38568 40979 38632
rect 41043 38568 41059 38632
rect 40932 38552 41059 38568
rect 40932 38488 40979 38552
rect 41043 38488 41059 38552
rect 40932 38472 41059 38488
rect 40932 38408 40979 38472
rect 41043 38408 41059 38472
rect 40932 38392 41059 38408
rect 40932 38328 40979 38392
rect 41043 38328 41059 38392
rect 40932 38312 41059 38328
rect 40932 38248 40979 38312
rect 41043 38248 41059 38312
rect 40932 38232 41059 38248
rect 40932 38168 40979 38232
rect 41043 38168 41059 38232
rect 40932 38152 41059 38168
rect 40932 38088 40979 38152
rect 41043 38088 41059 38152
rect 40932 38072 41059 38088
rect 40932 38008 40979 38072
rect 41043 38008 41059 38072
rect 40932 37992 41059 38008
rect 40932 37928 40979 37992
rect 41043 37928 41059 37992
rect 40932 37912 41059 37928
rect 40932 37848 40979 37912
rect 41043 37848 41059 37912
rect 40932 37832 41059 37848
rect 40932 37768 40979 37832
rect 41043 37768 41059 37832
rect 40932 37752 41059 37768
rect 40932 37688 40979 37752
rect 41043 37688 41059 37752
rect 40932 37672 41059 37688
rect 40932 37608 40979 37672
rect 41043 37608 41059 37672
rect 40932 37592 41059 37608
rect 40932 37528 40979 37592
rect 41043 37528 41059 37592
rect 40932 37512 41059 37528
rect 40932 37448 40979 37512
rect 41043 37448 41059 37512
rect 40932 37432 41059 37448
rect 40932 37368 40979 37432
rect 41043 37368 41059 37432
rect 40932 37352 41059 37368
rect 40932 37288 40979 37352
rect 41043 37288 41059 37352
rect 40932 37272 41059 37288
rect 40932 37208 40979 37272
rect 41043 37208 41059 37272
rect 40932 37192 41059 37208
rect 40932 37128 40979 37192
rect 41043 37128 41059 37192
rect 40932 37112 41059 37128
rect 40932 37048 40979 37112
rect 41043 37048 41059 37112
rect 40932 37032 41059 37048
rect 40932 36968 40979 37032
rect 41043 36968 41059 37032
rect 40932 36952 41059 36968
rect 40932 36888 40979 36952
rect 41043 36888 41059 36952
rect 40932 36872 41059 36888
rect 40932 36808 40979 36872
rect 41043 36808 41059 36872
rect 40932 36792 41059 36808
rect 40932 36728 40979 36792
rect 41043 36728 41059 36792
rect 40932 36712 41059 36728
rect 40932 36648 40979 36712
rect 41043 36648 41059 36712
rect 40932 36632 41059 36648
rect 40932 36568 40979 36632
rect 41043 36568 41059 36632
rect 40932 36552 41059 36568
rect 40932 36488 40979 36552
rect 41043 36488 41059 36552
rect 40932 36472 41059 36488
rect 40932 36408 40979 36472
rect 41043 36408 41059 36472
rect 40932 36392 41059 36408
rect 40932 36328 40979 36392
rect 41043 36328 41059 36392
rect 40932 36312 41059 36328
rect 40932 36248 40979 36312
rect 41043 36248 41059 36312
rect 40932 36232 41059 36248
rect 40932 36168 40979 36232
rect 41043 36168 41059 36232
rect 40932 36152 41059 36168
rect 40932 36088 40979 36152
rect 41043 36088 41059 36152
rect 40932 36072 41059 36088
rect 40932 36008 40979 36072
rect 41043 36008 41059 36072
rect 40932 35992 41059 36008
rect 40932 35928 40979 35992
rect 41043 35928 41059 35992
rect 40932 35912 41059 35928
rect 40932 35848 40979 35912
rect 41043 35848 41059 35912
rect 40932 35832 41059 35848
rect 40932 35768 40979 35832
rect 41043 35768 41059 35832
rect 40932 35752 41059 35768
rect 40932 35688 40979 35752
rect 41043 35688 41059 35752
rect 40932 35672 41059 35688
rect 40932 35608 40979 35672
rect 41043 35608 41059 35672
rect 40932 35592 41059 35608
rect 40932 35528 40979 35592
rect 41043 35528 41059 35592
rect 40932 35512 41059 35528
rect 40932 35448 40979 35512
rect 41043 35448 41059 35512
rect 40932 35432 41059 35448
rect 40932 35368 40979 35432
rect 41043 35368 41059 35432
rect 40932 35352 41059 35368
rect 40932 35288 40979 35352
rect 41043 35288 41059 35352
rect 40932 35272 41059 35288
rect 40932 35208 40979 35272
rect 41043 35208 41059 35272
rect 40932 35192 41059 35208
rect 40932 35128 40979 35192
rect 41043 35128 41059 35192
rect 40932 35112 41059 35128
rect 40932 35048 40979 35112
rect 41043 35048 41059 35112
rect 40932 35032 41059 35048
rect 40932 34968 40979 35032
rect 41043 34968 41059 35032
rect 40932 34952 41059 34968
rect 40932 34888 40979 34952
rect 41043 34888 41059 34952
rect 40932 34872 41059 34888
rect 34613 34792 34740 34808
rect 34613 34728 34660 34792
rect 34724 34728 34740 34792
rect 34613 34712 34740 34728
rect 34613 34588 34717 34712
rect 34613 34572 34740 34588
rect 34613 34508 34660 34572
rect 34724 34508 34740 34572
rect 34613 34492 34740 34508
rect 28294 34412 28421 34428
rect 28294 34348 28341 34412
rect 28405 34348 28421 34412
rect 28294 34332 28421 34348
rect 28294 34268 28341 34332
rect 28405 34268 28421 34332
rect 28294 34252 28421 34268
rect 28294 34188 28341 34252
rect 28405 34188 28421 34252
rect 28294 34172 28421 34188
rect 28294 34108 28341 34172
rect 28405 34108 28421 34172
rect 28294 34092 28421 34108
rect 28294 34028 28341 34092
rect 28405 34028 28421 34092
rect 28294 34012 28421 34028
rect 28294 33948 28341 34012
rect 28405 33948 28421 34012
rect 28294 33932 28421 33948
rect 28294 33868 28341 33932
rect 28405 33868 28421 33932
rect 28294 33852 28421 33868
rect 28294 33788 28341 33852
rect 28405 33788 28421 33852
rect 28294 33772 28421 33788
rect 28294 33708 28341 33772
rect 28405 33708 28421 33772
rect 28294 33692 28421 33708
rect 28294 33628 28341 33692
rect 28405 33628 28421 33692
rect 28294 33612 28421 33628
rect 28294 33548 28341 33612
rect 28405 33548 28421 33612
rect 28294 33532 28421 33548
rect 28294 33468 28341 33532
rect 28405 33468 28421 33532
rect 28294 33452 28421 33468
rect 28294 33388 28341 33452
rect 28405 33388 28421 33452
rect 28294 33372 28421 33388
rect 28294 33308 28341 33372
rect 28405 33308 28421 33372
rect 28294 33292 28421 33308
rect 28294 33228 28341 33292
rect 28405 33228 28421 33292
rect 28294 33212 28421 33228
rect 28294 33148 28341 33212
rect 28405 33148 28421 33212
rect 28294 33132 28421 33148
rect 28294 33068 28341 33132
rect 28405 33068 28421 33132
rect 28294 33052 28421 33068
rect 28294 32988 28341 33052
rect 28405 32988 28421 33052
rect 28294 32972 28421 32988
rect 28294 32908 28341 32972
rect 28405 32908 28421 32972
rect 28294 32892 28421 32908
rect 28294 32828 28341 32892
rect 28405 32828 28421 32892
rect 28294 32812 28421 32828
rect 28294 32748 28341 32812
rect 28405 32748 28421 32812
rect 28294 32732 28421 32748
rect 28294 32668 28341 32732
rect 28405 32668 28421 32732
rect 28294 32652 28421 32668
rect 28294 32588 28341 32652
rect 28405 32588 28421 32652
rect 28294 32572 28421 32588
rect 28294 32508 28341 32572
rect 28405 32508 28421 32572
rect 28294 32492 28421 32508
rect 28294 32428 28341 32492
rect 28405 32428 28421 32492
rect 28294 32412 28421 32428
rect 28294 32348 28341 32412
rect 28405 32348 28421 32412
rect 28294 32332 28421 32348
rect 28294 32268 28341 32332
rect 28405 32268 28421 32332
rect 28294 32252 28421 32268
rect 28294 32188 28341 32252
rect 28405 32188 28421 32252
rect 28294 32172 28421 32188
rect 28294 32108 28341 32172
rect 28405 32108 28421 32172
rect 28294 32092 28421 32108
rect 28294 32028 28341 32092
rect 28405 32028 28421 32092
rect 28294 32012 28421 32028
rect 28294 31948 28341 32012
rect 28405 31948 28421 32012
rect 28294 31932 28421 31948
rect 28294 31868 28341 31932
rect 28405 31868 28421 31932
rect 28294 31852 28421 31868
rect 28294 31788 28341 31852
rect 28405 31788 28421 31852
rect 28294 31772 28421 31788
rect 28294 31708 28341 31772
rect 28405 31708 28421 31772
rect 28294 31692 28421 31708
rect 28294 31628 28341 31692
rect 28405 31628 28421 31692
rect 28294 31612 28421 31628
rect 28294 31548 28341 31612
rect 28405 31548 28421 31612
rect 28294 31532 28421 31548
rect 28294 31468 28341 31532
rect 28405 31468 28421 31532
rect 28294 31452 28421 31468
rect 28294 31388 28341 31452
rect 28405 31388 28421 31452
rect 28294 31372 28421 31388
rect 28294 31308 28341 31372
rect 28405 31308 28421 31372
rect 28294 31292 28421 31308
rect 28294 31228 28341 31292
rect 28405 31228 28421 31292
rect 28294 31212 28421 31228
rect 28294 31148 28341 31212
rect 28405 31148 28421 31212
rect 28294 31132 28421 31148
rect 28294 31068 28341 31132
rect 28405 31068 28421 31132
rect 28294 31052 28421 31068
rect 28294 30988 28341 31052
rect 28405 30988 28421 31052
rect 28294 30972 28421 30988
rect 28294 30908 28341 30972
rect 28405 30908 28421 30972
rect 28294 30892 28421 30908
rect 28294 30828 28341 30892
rect 28405 30828 28421 30892
rect 28294 30812 28421 30828
rect 28294 30748 28341 30812
rect 28405 30748 28421 30812
rect 28294 30732 28421 30748
rect 28294 30668 28341 30732
rect 28405 30668 28421 30732
rect 28294 30652 28421 30668
rect 28294 30588 28341 30652
rect 28405 30588 28421 30652
rect 28294 30572 28421 30588
rect 28294 30508 28341 30572
rect 28405 30508 28421 30572
rect 28294 30492 28421 30508
rect 28294 30428 28341 30492
rect 28405 30428 28421 30492
rect 28294 30412 28421 30428
rect 28294 30348 28341 30412
rect 28405 30348 28421 30412
rect 28294 30332 28421 30348
rect 28294 30268 28341 30332
rect 28405 30268 28421 30332
rect 28294 30252 28421 30268
rect 28294 30188 28341 30252
rect 28405 30188 28421 30252
rect 28294 30172 28421 30188
rect 28294 30108 28341 30172
rect 28405 30108 28421 30172
rect 28294 30092 28421 30108
rect 28294 30028 28341 30092
rect 28405 30028 28421 30092
rect 28294 30012 28421 30028
rect 28294 29948 28341 30012
rect 28405 29948 28421 30012
rect 28294 29932 28421 29948
rect 28294 29868 28341 29932
rect 28405 29868 28421 29932
rect 28294 29852 28421 29868
rect 28294 29788 28341 29852
rect 28405 29788 28421 29852
rect 28294 29772 28421 29788
rect 28294 29708 28341 29772
rect 28405 29708 28421 29772
rect 28294 29692 28421 29708
rect 28294 29628 28341 29692
rect 28405 29628 28421 29692
rect 28294 29612 28421 29628
rect 28294 29548 28341 29612
rect 28405 29548 28421 29612
rect 28294 29532 28421 29548
rect 28294 29468 28341 29532
rect 28405 29468 28421 29532
rect 28294 29452 28421 29468
rect 28294 29388 28341 29452
rect 28405 29388 28421 29452
rect 28294 29372 28421 29388
rect 28294 29308 28341 29372
rect 28405 29308 28421 29372
rect 28294 29292 28421 29308
rect 28294 29228 28341 29292
rect 28405 29228 28421 29292
rect 28294 29212 28421 29228
rect 28294 29148 28341 29212
rect 28405 29148 28421 29212
rect 28294 29132 28421 29148
rect 28294 29068 28341 29132
rect 28405 29068 28421 29132
rect 28294 29052 28421 29068
rect 28294 28988 28341 29052
rect 28405 28988 28421 29052
rect 28294 28972 28421 28988
rect 28294 28908 28341 28972
rect 28405 28908 28421 28972
rect 28294 28892 28421 28908
rect 28294 28828 28341 28892
rect 28405 28828 28421 28892
rect 28294 28812 28421 28828
rect 28294 28748 28341 28812
rect 28405 28748 28421 28812
rect 28294 28732 28421 28748
rect 28294 28668 28341 28732
rect 28405 28668 28421 28732
rect 28294 28652 28421 28668
rect 28294 28588 28341 28652
rect 28405 28588 28421 28652
rect 28294 28572 28421 28588
rect 21975 28492 22102 28508
rect 21975 28428 22022 28492
rect 22086 28428 22102 28492
rect 21975 28412 22102 28428
rect 21975 28288 22079 28412
rect 21975 28272 22102 28288
rect 21975 28208 22022 28272
rect 22086 28208 22102 28272
rect 21975 28192 22102 28208
rect 15656 28112 15783 28128
rect 15656 28048 15703 28112
rect 15767 28048 15783 28112
rect 15656 28032 15783 28048
rect 15656 27968 15703 28032
rect 15767 27968 15783 28032
rect 15656 27952 15783 27968
rect 15656 27888 15703 27952
rect 15767 27888 15783 27952
rect 15656 27872 15783 27888
rect 15656 27808 15703 27872
rect 15767 27808 15783 27872
rect 15656 27792 15783 27808
rect 15656 27728 15703 27792
rect 15767 27728 15783 27792
rect 15656 27712 15783 27728
rect 15656 27648 15703 27712
rect 15767 27648 15783 27712
rect 15656 27632 15783 27648
rect 15656 27568 15703 27632
rect 15767 27568 15783 27632
rect 15656 27552 15783 27568
rect 15656 27488 15703 27552
rect 15767 27488 15783 27552
rect 15656 27472 15783 27488
rect 15656 27408 15703 27472
rect 15767 27408 15783 27472
rect 15656 27392 15783 27408
rect 15656 27328 15703 27392
rect 15767 27328 15783 27392
rect 15656 27312 15783 27328
rect 15656 27248 15703 27312
rect 15767 27248 15783 27312
rect 15656 27232 15783 27248
rect 15656 27168 15703 27232
rect 15767 27168 15783 27232
rect 15656 27152 15783 27168
rect 15656 27088 15703 27152
rect 15767 27088 15783 27152
rect 15656 27072 15783 27088
rect 15656 27008 15703 27072
rect 15767 27008 15783 27072
rect 15656 26992 15783 27008
rect 15656 26928 15703 26992
rect 15767 26928 15783 26992
rect 15656 26912 15783 26928
rect 15656 26848 15703 26912
rect 15767 26848 15783 26912
rect 15656 26832 15783 26848
rect 15656 26768 15703 26832
rect 15767 26768 15783 26832
rect 15656 26752 15783 26768
rect 15656 26688 15703 26752
rect 15767 26688 15783 26752
rect 15656 26672 15783 26688
rect 15656 26608 15703 26672
rect 15767 26608 15783 26672
rect 15656 26592 15783 26608
rect 15656 26528 15703 26592
rect 15767 26528 15783 26592
rect 15656 26512 15783 26528
rect 15656 26448 15703 26512
rect 15767 26448 15783 26512
rect 15656 26432 15783 26448
rect 15656 26368 15703 26432
rect 15767 26368 15783 26432
rect 15656 26352 15783 26368
rect 15656 26288 15703 26352
rect 15767 26288 15783 26352
rect 15656 26272 15783 26288
rect 15656 26208 15703 26272
rect 15767 26208 15783 26272
rect 15656 26192 15783 26208
rect 15656 26128 15703 26192
rect 15767 26128 15783 26192
rect 15656 26112 15783 26128
rect 15656 26048 15703 26112
rect 15767 26048 15783 26112
rect 15656 26032 15783 26048
rect 15656 25968 15703 26032
rect 15767 25968 15783 26032
rect 15656 25952 15783 25968
rect 15656 25888 15703 25952
rect 15767 25888 15783 25952
rect 15656 25872 15783 25888
rect 15656 25808 15703 25872
rect 15767 25808 15783 25872
rect 15656 25792 15783 25808
rect 15656 25728 15703 25792
rect 15767 25728 15783 25792
rect 15656 25712 15783 25728
rect 15656 25648 15703 25712
rect 15767 25648 15783 25712
rect 15656 25632 15783 25648
rect 15656 25568 15703 25632
rect 15767 25568 15783 25632
rect 15656 25552 15783 25568
rect 15656 25488 15703 25552
rect 15767 25488 15783 25552
rect 15656 25472 15783 25488
rect 15656 25408 15703 25472
rect 15767 25408 15783 25472
rect 15656 25392 15783 25408
rect 15656 25328 15703 25392
rect 15767 25328 15783 25392
rect 15656 25312 15783 25328
rect 15656 25248 15703 25312
rect 15767 25248 15783 25312
rect 15656 25232 15783 25248
rect 15656 25168 15703 25232
rect 15767 25168 15783 25232
rect 15656 25152 15783 25168
rect 15656 25088 15703 25152
rect 15767 25088 15783 25152
rect 15656 25072 15783 25088
rect 15656 25008 15703 25072
rect 15767 25008 15783 25072
rect 15656 24992 15783 25008
rect 15656 24928 15703 24992
rect 15767 24928 15783 24992
rect 15656 24912 15783 24928
rect 15656 24848 15703 24912
rect 15767 24848 15783 24912
rect 15656 24832 15783 24848
rect 15656 24768 15703 24832
rect 15767 24768 15783 24832
rect 15656 24752 15783 24768
rect 15656 24688 15703 24752
rect 15767 24688 15783 24752
rect 15656 24672 15783 24688
rect 15656 24608 15703 24672
rect 15767 24608 15783 24672
rect 15656 24592 15783 24608
rect 15656 24528 15703 24592
rect 15767 24528 15783 24592
rect 15656 24512 15783 24528
rect 15656 24448 15703 24512
rect 15767 24448 15783 24512
rect 15656 24432 15783 24448
rect 15656 24368 15703 24432
rect 15767 24368 15783 24432
rect 15656 24352 15783 24368
rect 15656 24288 15703 24352
rect 15767 24288 15783 24352
rect 15656 24272 15783 24288
rect 15656 24208 15703 24272
rect 15767 24208 15783 24272
rect 15656 24192 15783 24208
rect 15656 24128 15703 24192
rect 15767 24128 15783 24192
rect 15656 24112 15783 24128
rect 15656 24048 15703 24112
rect 15767 24048 15783 24112
rect 15656 24032 15783 24048
rect 15656 23968 15703 24032
rect 15767 23968 15783 24032
rect 15656 23952 15783 23968
rect 15656 23888 15703 23952
rect 15767 23888 15783 23952
rect 15656 23872 15783 23888
rect 15656 23808 15703 23872
rect 15767 23808 15783 23872
rect 15656 23792 15783 23808
rect 15656 23728 15703 23792
rect 15767 23728 15783 23792
rect 15656 23712 15783 23728
rect 15656 23648 15703 23712
rect 15767 23648 15783 23712
rect 15656 23632 15783 23648
rect 15656 23568 15703 23632
rect 15767 23568 15783 23632
rect 15656 23552 15783 23568
rect 15656 23488 15703 23552
rect 15767 23488 15783 23552
rect 15656 23472 15783 23488
rect 15656 23408 15703 23472
rect 15767 23408 15783 23472
rect 15656 23392 15783 23408
rect 15656 23328 15703 23392
rect 15767 23328 15783 23392
rect 15656 23312 15783 23328
rect 15656 23248 15703 23312
rect 15767 23248 15783 23312
rect 15656 23232 15783 23248
rect 15656 23168 15703 23232
rect 15767 23168 15783 23232
rect 15656 23152 15783 23168
rect 15656 23088 15703 23152
rect 15767 23088 15783 23152
rect 15656 23072 15783 23088
rect 15656 23008 15703 23072
rect 15767 23008 15783 23072
rect 15656 22992 15783 23008
rect 15656 22928 15703 22992
rect 15767 22928 15783 22992
rect 15656 22912 15783 22928
rect 15656 22848 15703 22912
rect 15767 22848 15783 22912
rect 15656 22832 15783 22848
rect 15656 22768 15703 22832
rect 15767 22768 15783 22832
rect 15656 22752 15783 22768
rect 15656 22688 15703 22752
rect 15767 22688 15783 22752
rect 15656 22672 15783 22688
rect 15656 22608 15703 22672
rect 15767 22608 15783 22672
rect 15656 22592 15783 22608
rect 15656 22528 15703 22592
rect 15767 22528 15783 22592
rect 15656 22512 15783 22528
rect 15656 22448 15703 22512
rect 15767 22448 15783 22512
rect 15656 22432 15783 22448
rect 15656 22368 15703 22432
rect 15767 22368 15783 22432
rect 15656 22352 15783 22368
rect 15656 22288 15703 22352
rect 15767 22288 15783 22352
rect 15656 22272 15783 22288
rect 9337 22192 9464 22208
rect 9337 22128 9384 22192
rect 9448 22128 9464 22192
rect 9337 22112 9464 22128
rect 9337 21988 9441 22112
rect 9337 21972 9464 21988
rect 9337 21908 9384 21972
rect 9448 21908 9464 21972
rect 9337 21892 9464 21908
rect 3018 21812 3145 21828
rect 3018 21748 3065 21812
rect 3129 21748 3145 21812
rect 3018 21732 3145 21748
rect 3018 21668 3065 21732
rect 3129 21668 3145 21732
rect 3018 21652 3145 21668
rect 3018 21588 3065 21652
rect 3129 21588 3145 21652
rect 3018 21572 3145 21588
rect 3018 21508 3065 21572
rect 3129 21508 3145 21572
rect 3018 21492 3145 21508
rect 3018 21428 3065 21492
rect 3129 21428 3145 21492
rect 3018 21412 3145 21428
rect 3018 21348 3065 21412
rect 3129 21348 3145 21412
rect 3018 21332 3145 21348
rect 3018 21268 3065 21332
rect 3129 21268 3145 21332
rect 3018 21252 3145 21268
rect 3018 21188 3065 21252
rect 3129 21188 3145 21252
rect 3018 21172 3145 21188
rect 3018 21108 3065 21172
rect 3129 21108 3145 21172
rect 3018 21092 3145 21108
rect 3018 21028 3065 21092
rect 3129 21028 3145 21092
rect 3018 21012 3145 21028
rect 3018 20948 3065 21012
rect 3129 20948 3145 21012
rect 3018 20932 3145 20948
rect 3018 20868 3065 20932
rect 3129 20868 3145 20932
rect 3018 20852 3145 20868
rect 3018 20788 3065 20852
rect 3129 20788 3145 20852
rect 3018 20772 3145 20788
rect 3018 20708 3065 20772
rect 3129 20708 3145 20772
rect 3018 20692 3145 20708
rect 3018 20628 3065 20692
rect 3129 20628 3145 20692
rect 3018 20612 3145 20628
rect 3018 20548 3065 20612
rect 3129 20548 3145 20612
rect 3018 20532 3145 20548
rect 3018 20468 3065 20532
rect 3129 20468 3145 20532
rect 3018 20452 3145 20468
rect 3018 20388 3065 20452
rect 3129 20388 3145 20452
rect 3018 20372 3145 20388
rect 3018 20308 3065 20372
rect 3129 20308 3145 20372
rect 3018 20292 3145 20308
rect 3018 20228 3065 20292
rect 3129 20228 3145 20292
rect 3018 20212 3145 20228
rect 3018 20148 3065 20212
rect 3129 20148 3145 20212
rect 3018 20132 3145 20148
rect 3018 20068 3065 20132
rect 3129 20068 3145 20132
rect 3018 20052 3145 20068
rect 3018 19988 3065 20052
rect 3129 19988 3145 20052
rect 3018 19972 3145 19988
rect 3018 19908 3065 19972
rect 3129 19908 3145 19972
rect 3018 19892 3145 19908
rect 3018 19828 3065 19892
rect 3129 19828 3145 19892
rect 3018 19812 3145 19828
rect 3018 19748 3065 19812
rect 3129 19748 3145 19812
rect 3018 19732 3145 19748
rect 3018 19668 3065 19732
rect 3129 19668 3145 19732
rect 3018 19652 3145 19668
rect 3018 19588 3065 19652
rect 3129 19588 3145 19652
rect 3018 19572 3145 19588
rect 3018 19508 3065 19572
rect 3129 19508 3145 19572
rect 3018 19492 3145 19508
rect 3018 19428 3065 19492
rect 3129 19428 3145 19492
rect 3018 19412 3145 19428
rect 3018 19348 3065 19412
rect 3129 19348 3145 19412
rect 3018 19332 3145 19348
rect 3018 19268 3065 19332
rect 3129 19268 3145 19332
rect 3018 19252 3145 19268
rect 3018 19188 3065 19252
rect 3129 19188 3145 19252
rect 3018 19172 3145 19188
rect 3018 19108 3065 19172
rect 3129 19108 3145 19172
rect 3018 19092 3145 19108
rect 3018 19028 3065 19092
rect 3129 19028 3145 19092
rect 3018 19012 3145 19028
rect 3018 18948 3065 19012
rect 3129 18948 3145 19012
rect 3018 18932 3145 18948
rect 3018 18868 3065 18932
rect 3129 18868 3145 18932
rect 3018 18852 3145 18868
rect 3018 18788 3065 18852
rect 3129 18788 3145 18852
rect 3018 18772 3145 18788
rect 3018 18708 3065 18772
rect 3129 18708 3145 18772
rect 3018 18692 3145 18708
rect 3018 18628 3065 18692
rect 3129 18628 3145 18692
rect 3018 18612 3145 18628
rect 3018 18548 3065 18612
rect 3129 18548 3145 18612
rect 3018 18532 3145 18548
rect 3018 18468 3065 18532
rect 3129 18468 3145 18532
rect 3018 18452 3145 18468
rect 3018 18388 3065 18452
rect 3129 18388 3145 18452
rect 3018 18372 3145 18388
rect 3018 18308 3065 18372
rect 3129 18308 3145 18372
rect 3018 18292 3145 18308
rect 3018 18228 3065 18292
rect 3129 18228 3145 18292
rect 3018 18212 3145 18228
rect 3018 18148 3065 18212
rect 3129 18148 3145 18212
rect 3018 18132 3145 18148
rect 3018 18068 3065 18132
rect 3129 18068 3145 18132
rect 3018 18052 3145 18068
rect 3018 17988 3065 18052
rect 3129 17988 3145 18052
rect 3018 17972 3145 17988
rect 3018 17908 3065 17972
rect 3129 17908 3145 17972
rect 3018 17892 3145 17908
rect 3018 17828 3065 17892
rect 3129 17828 3145 17892
rect 3018 17812 3145 17828
rect 3018 17748 3065 17812
rect 3129 17748 3145 17812
rect 3018 17732 3145 17748
rect 3018 17668 3065 17732
rect 3129 17668 3145 17732
rect 3018 17652 3145 17668
rect 3018 17588 3065 17652
rect 3129 17588 3145 17652
rect 3018 17572 3145 17588
rect 3018 17508 3065 17572
rect 3129 17508 3145 17572
rect 3018 17492 3145 17508
rect 3018 17428 3065 17492
rect 3129 17428 3145 17492
rect 3018 17412 3145 17428
rect 3018 17348 3065 17412
rect 3129 17348 3145 17412
rect 3018 17332 3145 17348
rect 3018 17268 3065 17332
rect 3129 17268 3145 17332
rect 3018 17252 3145 17268
rect 3018 17188 3065 17252
rect 3129 17188 3145 17252
rect 3018 17172 3145 17188
rect 3018 17108 3065 17172
rect 3129 17108 3145 17172
rect 3018 17092 3145 17108
rect 3018 17028 3065 17092
rect 3129 17028 3145 17092
rect 3018 17012 3145 17028
rect 3018 16948 3065 17012
rect 3129 16948 3145 17012
rect 3018 16932 3145 16948
rect 3018 16868 3065 16932
rect 3129 16868 3145 16932
rect 3018 16852 3145 16868
rect 3018 16788 3065 16852
rect 3129 16788 3145 16852
rect 3018 16772 3145 16788
rect 3018 16708 3065 16772
rect 3129 16708 3145 16772
rect 3018 16692 3145 16708
rect 3018 16628 3065 16692
rect 3129 16628 3145 16692
rect 3018 16612 3145 16628
rect 3018 16548 3065 16612
rect 3129 16548 3145 16612
rect 3018 16532 3145 16548
rect 3018 16468 3065 16532
rect 3129 16468 3145 16532
rect 3018 16452 3145 16468
rect 3018 16388 3065 16452
rect 3129 16388 3145 16452
rect 3018 16372 3145 16388
rect 3018 16308 3065 16372
rect 3129 16308 3145 16372
rect 3018 16292 3145 16308
rect 3018 16228 3065 16292
rect 3129 16228 3145 16292
rect 3018 16212 3145 16228
rect 3018 16148 3065 16212
rect 3129 16148 3145 16212
rect 3018 16132 3145 16148
rect 3018 16068 3065 16132
rect 3129 16068 3145 16132
rect 3018 16052 3145 16068
rect 3018 15988 3065 16052
rect 3129 15988 3145 16052
rect 3018 15972 3145 15988
rect -3301 15892 -3174 15908
rect -3301 15828 -3254 15892
rect -3190 15828 -3174 15892
rect -3301 15812 -3174 15828
rect -3301 15688 -3197 15812
rect -3301 15672 -3174 15688
rect -3301 15608 -3254 15672
rect -3190 15608 -3174 15672
rect -3301 15592 -3174 15608
rect -9620 15512 -9493 15528
rect -9620 15448 -9573 15512
rect -9509 15448 -9493 15512
rect -9620 15432 -9493 15448
rect -9620 15368 -9573 15432
rect -9509 15368 -9493 15432
rect -9620 15352 -9493 15368
rect -9620 15288 -9573 15352
rect -9509 15288 -9493 15352
rect -9620 15272 -9493 15288
rect -9620 15208 -9573 15272
rect -9509 15208 -9493 15272
rect -9620 15192 -9493 15208
rect -9620 15128 -9573 15192
rect -9509 15128 -9493 15192
rect -9620 15112 -9493 15128
rect -9620 15048 -9573 15112
rect -9509 15048 -9493 15112
rect -9620 15032 -9493 15048
rect -9620 14968 -9573 15032
rect -9509 14968 -9493 15032
rect -9620 14952 -9493 14968
rect -9620 14888 -9573 14952
rect -9509 14888 -9493 14952
rect -9620 14872 -9493 14888
rect -9620 14808 -9573 14872
rect -9509 14808 -9493 14872
rect -9620 14792 -9493 14808
rect -9620 14728 -9573 14792
rect -9509 14728 -9493 14792
rect -9620 14712 -9493 14728
rect -9620 14648 -9573 14712
rect -9509 14648 -9493 14712
rect -9620 14632 -9493 14648
rect -9620 14568 -9573 14632
rect -9509 14568 -9493 14632
rect -9620 14552 -9493 14568
rect -9620 14488 -9573 14552
rect -9509 14488 -9493 14552
rect -9620 14472 -9493 14488
rect -9620 14408 -9573 14472
rect -9509 14408 -9493 14472
rect -9620 14392 -9493 14408
rect -9620 14328 -9573 14392
rect -9509 14328 -9493 14392
rect -9620 14312 -9493 14328
rect -9620 14248 -9573 14312
rect -9509 14248 -9493 14312
rect -9620 14232 -9493 14248
rect -9620 14168 -9573 14232
rect -9509 14168 -9493 14232
rect -9620 14152 -9493 14168
rect -9620 14088 -9573 14152
rect -9509 14088 -9493 14152
rect -9620 14072 -9493 14088
rect -9620 14008 -9573 14072
rect -9509 14008 -9493 14072
rect -9620 13992 -9493 14008
rect -9620 13928 -9573 13992
rect -9509 13928 -9493 13992
rect -9620 13912 -9493 13928
rect -9620 13848 -9573 13912
rect -9509 13848 -9493 13912
rect -9620 13832 -9493 13848
rect -9620 13768 -9573 13832
rect -9509 13768 -9493 13832
rect -9620 13752 -9493 13768
rect -9620 13688 -9573 13752
rect -9509 13688 -9493 13752
rect -9620 13672 -9493 13688
rect -9620 13608 -9573 13672
rect -9509 13608 -9493 13672
rect -9620 13592 -9493 13608
rect -9620 13528 -9573 13592
rect -9509 13528 -9493 13592
rect -9620 13512 -9493 13528
rect -9620 13448 -9573 13512
rect -9509 13448 -9493 13512
rect -9620 13432 -9493 13448
rect -9620 13368 -9573 13432
rect -9509 13368 -9493 13432
rect -9620 13352 -9493 13368
rect -9620 13288 -9573 13352
rect -9509 13288 -9493 13352
rect -9620 13272 -9493 13288
rect -9620 13208 -9573 13272
rect -9509 13208 -9493 13272
rect -9620 13192 -9493 13208
rect -9620 13128 -9573 13192
rect -9509 13128 -9493 13192
rect -9620 13112 -9493 13128
rect -9620 13048 -9573 13112
rect -9509 13048 -9493 13112
rect -9620 13032 -9493 13048
rect -9620 12968 -9573 13032
rect -9509 12968 -9493 13032
rect -9620 12952 -9493 12968
rect -9620 12888 -9573 12952
rect -9509 12888 -9493 12952
rect -9620 12872 -9493 12888
rect -9620 12808 -9573 12872
rect -9509 12808 -9493 12872
rect -9620 12792 -9493 12808
rect -9620 12728 -9573 12792
rect -9509 12728 -9493 12792
rect -9620 12712 -9493 12728
rect -9620 12648 -9573 12712
rect -9509 12648 -9493 12712
rect -9620 12632 -9493 12648
rect -9620 12568 -9573 12632
rect -9509 12568 -9493 12632
rect -9620 12552 -9493 12568
rect -9620 12488 -9573 12552
rect -9509 12488 -9493 12552
rect -9620 12472 -9493 12488
rect -9620 12408 -9573 12472
rect -9509 12408 -9493 12472
rect -9620 12392 -9493 12408
rect -9620 12328 -9573 12392
rect -9509 12328 -9493 12392
rect -9620 12312 -9493 12328
rect -9620 12248 -9573 12312
rect -9509 12248 -9493 12312
rect -9620 12232 -9493 12248
rect -9620 12168 -9573 12232
rect -9509 12168 -9493 12232
rect -9620 12152 -9493 12168
rect -9620 12088 -9573 12152
rect -9509 12088 -9493 12152
rect -9620 12072 -9493 12088
rect -9620 12008 -9573 12072
rect -9509 12008 -9493 12072
rect -9620 11992 -9493 12008
rect -9620 11928 -9573 11992
rect -9509 11928 -9493 11992
rect -9620 11912 -9493 11928
rect -9620 11848 -9573 11912
rect -9509 11848 -9493 11912
rect -9620 11832 -9493 11848
rect -9620 11768 -9573 11832
rect -9509 11768 -9493 11832
rect -9620 11752 -9493 11768
rect -9620 11688 -9573 11752
rect -9509 11688 -9493 11752
rect -9620 11672 -9493 11688
rect -9620 11608 -9573 11672
rect -9509 11608 -9493 11672
rect -9620 11592 -9493 11608
rect -9620 11528 -9573 11592
rect -9509 11528 -9493 11592
rect -9620 11512 -9493 11528
rect -9620 11448 -9573 11512
rect -9509 11448 -9493 11512
rect -9620 11432 -9493 11448
rect -9620 11368 -9573 11432
rect -9509 11368 -9493 11432
rect -9620 11352 -9493 11368
rect -9620 11288 -9573 11352
rect -9509 11288 -9493 11352
rect -9620 11272 -9493 11288
rect -9620 11208 -9573 11272
rect -9509 11208 -9493 11272
rect -9620 11192 -9493 11208
rect -9620 11128 -9573 11192
rect -9509 11128 -9493 11192
rect -9620 11112 -9493 11128
rect -9620 11048 -9573 11112
rect -9509 11048 -9493 11112
rect -9620 11032 -9493 11048
rect -9620 10968 -9573 11032
rect -9509 10968 -9493 11032
rect -9620 10952 -9493 10968
rect -9620 10888 -9573 10952
rect -9509 10888 -9493 10952
rect -9620 10872 -9493 10888
rect -9620 10808 -9573 10872
rect -9509 10808 -9493 10872
rect -9620 10792 -9493 10808
rect -9620 10728 -9573 10792
rect -9509 10728 -9493 10792
rect -9620 10712 -9493 10728
rect -9620 10648 -9573 10712
rect -9509 10648 -9493 10712
rect -9620 10632 -9493 10648
rect -9620 10568 -9573 10632
rect -9509 10568 -9493 10632
rect -9620 10552 -9493 10568
rect -9620 10488 -9573 10552
rect -9509 10488 -9493 10552
rect -9620 10472 -9493 10488
rect -9620 10408 -9573 10472
rect -9509 10408 -9493 10472
rect -9620 10392 -9493 10408
rect -9620 10328 -9573 10392
rect -9509 10328 -9493 10392
rect -9620 10312 -9493 10328
rect -9620 10248 -9573 10312
rect -9509 10248 -9493 10312
rect -9620 10232 -9493 10248
rect -9620 10168 -9573 10232
rect -9509 10168 -9493 10232
rect -9620 10152 -9493 10168
rect -9620 10088 -9573 10152
rect -9509 10088 -9493 10152
rect -9620 10072 -9493 10088
rect -9620 10008 -9573 10072
rect -9509 10008 -9493 10072
rect -9620 9992 -9493 10008
rect -9620 9928 -9573 9992
rect -9509 9928 -9493 9992
rect -9620 9912 -9493 9928
rect -9620 9848 -9573 9912
rect -9509 9848 -9493 9912
rect -9620 9832 -9493 9848
rect -9620 9768 -9573 9832
rect -9509 9768 -9493 9832
rect -9620 9752 -9493 9768
rect -9620 9688 -9573 9752
rect -9509 9688 -9493 9752
rect -9620 9672 -9493 9688
rect -15939 9592 -15812 9608
rect -15939 9528 -15892 9592
rect -15828 9528 -15812 9592
rect -15939 9512 -15812 9528
rect -15939 9388 -15835 9512
rect -15939 9372 -15812 9388
rect -15939 9308 -15892 9372
rect -15828 9308 -15812 9372
rect -15939 9292 -15812 9308
rect -22258 9212 -22131 9228
rect -22258 9148 -22211 9212
rect -22147 9148 -22131 9212
rect -22258 9132 -22131 9148
rect -22258 9068 -22211 9132
rect -22147 9068 -22131 9132
rect -22258 9052 -22131 9068
rect -22258 8988 -22211 9052
rect -22147 8988 -22131 9052
rect -22258 8972 -22131 8988
rect -22258 8908 -22211 8972
rect -22147 8908 -22131 8972
rect -22258 8892 -22131 8908
rect -22258 8828 -22211 8892
rect -22147 8828 -22131 8892
rect -22258 8812 -22131 8828
rect -22258 8748 -22211 8812
rect -22147 8748 -22131 8812
rect -22258 8732 -22131 8748
rect -22258 8668 -22211 8732
rect -22147 8668 -22131 8732
rect -22258 8652 -22131 8668
rect -22258 8588 -22211 8652
rect -22147 8588 -22131 8652
rect -22258 8572 -22131 8588
rect -22258 8508 -22211 8572
rect -22147 8508 -22131 8572
rect -22258 8492 -22131 8508
rect -22258 8428 -22211 8492
rect -22147 8428 -22131 8492
rect -22258 8412 -22131 8428
rect -22258 8348 -22211 8412
rect -22147 8348 -22131 8412
rect -22258 8332 -22131 8348
rect -22258 8268 -22211 8332
rect -22147 8268 -22131 8332
rect -22258 8252 -22131 8268
rect -22258 8188 -22211 8252
rect -22147 8188 -22131 8252
rect -22258 8172 -22131 8188
rect -22258 8108 -22211 8172
rect -22147 8108 -22131 8172
rect -22258 8092 -22131 8108
rect -22258 8028 -22211 8092
rect -22147 8028 -22131 8092
rect -22258 8012 -22131 8028
rect -22258 7948 -22211 8012
rect -22147 7948 -22131 8012
rect -22258 7932 -22131 7948
rect -22258 7868 -22211 7932
rect -22147 7868 -22131 7932
rect -22258 7852 -22131 7868
rect -22258 7788 -22211 7852
rect -22147 7788 -22131 7852
rect -22258 7772 -22131 7788
rect -22258 7708 -22211 7772
rect -22147 7708 -22131 7772
rect -22258 7692 -22131 7708
rect -22258 7628 -22211 7692
rect -22147 7628 -22131 7692
rect -22258 7612 -22131 7628
rect -22258 7548 -22211 7612
rect -22147 7548 -22131 7612
rect -22258 7532 -22131 7548
rect -22258 7468 -22211 7532
rect -22147 7468 -22131 7532
rect -22258 7452 -22131 7468
rect -22258 7388 -22211 7452
rect -22147 7388 -22131 7452
rect -22258 7372 -22131 7388
rect -22258 7308 -22211 7372
rect -22147 7308 -22131 7372
rect -22258 7292 -22131 7308
rect -22258 7228 -22211 7292
rect -22147 7228 -22131 7292
rect -22258 7212 -22131 7228
rect -22258 7148 -22211 7212
rect -22147 7148 -22131 7212
rect -22258 7132 -22131 7148
rect -22258 7068 -22211 7132
rect -22147 7068 -22131 7132
rect -22258 7052 -22131 7068
rect -22258 6988 -22211 7052
rect -22147 6988 -22131 7052
rect -22258 6972 -22131 6988
rect -22258 6908 -22211 6972
rect -22147 6908 -22131 6972
rect -22258 6892 -22131 6908
rect -22258 6828 -22211 6892
rect -22147 6828 -22131 6892
rect -22258 6812 -22131 6828
rect -22258 6748 -22211 6812
rect -22147 6748 -22131 6812
rect -22258 6732 -22131 6748
rect -22258 6668 -22211 6732
rect -22147 6668 -22131 6732
rect -22258 6652 -22131 6668
rect -22258 6588 -22211 6652
rect -22147 6588 -22131 6652
rect -22258 6572 -22131 6588
rect -22258 6508 -22211 6572
rect -22147 6508 -22131 6572
rect -22258 6492 -22131 6508
rect -22258 6428 -22211 6492
rect -22147 6428 -22131 6492
rect -22258 6412 -22131 6428
rect -22258 6348 -22211 6412
rect -22147 6348 -22131 6412
rect -22258 6332 -22131 6348
rect -22258 6268 -22211 6332
rect -22147 6268 -22131 6332
rect -22258 6252 -22131 6268
rect -22258 6188 -22211 6252
rect -22147 6188 -22131 6252
rect -22258 6172 -22131 6188
rect -22258 6108 -22211 6172
rect -22147 6108 -22131 6172
rect -22258 6092 -22131 6108
rect -22258 6028 -22211 6092
rect -22147 6028 -22131 6092
rect -22258 6012 -22131 6028
rect -22258 5948 -22211 6012
rect -22147 5948 -22131 6012
rect -22258 5932 -22131 5948
rect -22258 5868 -22211 5932
rect -22147 5868 -22131 5932
rect -22258 5852 -22131 5868
rect -22258 5788 -22211 5852
rect -22147 5788 -22131 5852
rect -22258 5772 -22131 5788
rect -22258 5708 -22211 5772
rect -22147 5708 -22131 5772
rect -22258 5692 -22131 5708
rect -22258 5628 -22211 5692
rect -22147 5628 -22131 5692
rect -22258 5612 -22131 5628
rect -22258 5548 -22211 5612
rect -22147 5548 -22131 5612
rect -22258 5532 -22131 5548
rect -22258 5468 -22211 5532
rect -22147 5468 -22131 5532
rect -22258 5452 -22131 5468
rect -22258 5388 -22211 5452
rect -22147 5388 -22131 5452
rect -22258 5372 -22131 5388
rect -22258 5308 -22211 5372
rect -22147 5308 -22131 5372
rect -22258 5292 -22131 5308
rect -22258 5228 -22211 5292
rect -22147 5228 -22131 5292
rect -22258 5212 -22131 5228
rect -22258 5148 -22211 5212
rect -22147 5148 -22131 5212
rect -22258 5132 -22131 5148
rect -22258 5068 -22211 5132
rect -22147 5068 -22131 5132
rect -22258 5052 -22131 5068
rect -22258 4988 -22211 5052
rect -22147 4988 -22131 5052
rect -22258 4972 -22131 4988
rect -22258 4908 -22211 4972
rect -22147 4908 -22131 4972
rect -22258 4892 -22131 4908
rect -22258 4828 -22211 4892
rect -22147 4828 -22131 4892
rect -22258 4812 -22131 4828
rect -22258 4748 -22211 4812
rect -22147 4748 -22131 4812
rect -22258 4732 -22131 4748
rect -22258 4668 -22211 4732
rect -22147 4668 -22131 4732
rect -22258 4652 -22131 4668
rect -22258 4588 -22211 4652
rect -22147 4588 -22131 4652
rect -22258 4572 -22131 4588
rect -22258 4508 -22211 4572
rect -22147 4508 -22131 4572
rect -22258 4492 -22131 4508
rect -22258 4428 -22211 4492
rect -22147 4428 -22131 4492
rect -22258 4412 -22131 4428
rect -22258 4348 -22211 4412
rect -22147 4348 -22131 4412
rect -22258 4332 -22131 4348
rect -22258 4268 -22211 4332
rect -22147 4268 -22131 4332
rect -22258 4252 -22131 4268
rect -22258 4188 -22211 4252
rect -22147 4188 -22131 4252
rect -22258 4172 -22131 4188
rect -22258 4108 -22211 4172
rect -22147 4108 -22131 4172
rect -22258 4092 -22131 4108
rect -22258 4028 -22211 4092
rect -22147 4028 -22131 4092
rect -22258 4012 -22131 4028
rect -22258 3948 -22211 4012
rect -22147 3948 -22131 4012
rect -22258 3932 -22131 3948
rect -22258 3868 -22211 3932
rect -22147 3868 -22131 3932
rect -22258 3852 -22131 3868
rect -22258 3788 -22211 3852
rect -22147 3788 -22131 3852
rect -22258 3772 -22131 3788
rect -22258 3708 -22211 3772
rect -22147 3708 -22131 3772
rect -22258 3692 -22131 3708
rect -22258 3628 -22211 3692
rect -22147 3628 -22131 3692
rect -22258 3612 -22131 3628
rect -22258 3548 -22211 3612
rect -22147 3548 -22131 3612
rect -22258 3532 -22131 3548
rect -22258 3468 -22211 3532
rect -22147 3468 -22131 3532
rect -22258 3452 -22131 3468
rect -22258 3388 -22211 3452
rect -22147 3388 -22131 3452
rect -22258 3372 -22131 3388
rect -28577 3292 -28450 3308
rect -28577 3228 -28530 3292
rect -28466 3228 -28450 3292
rect -28577 3212 -28450 3228
rect -28577 3088 -28473 3212
rect -28577 3072 -28450 3088
rect -28577 3008 -28530 3072
rect -28466 3008 -28450 3072
rect -28577 2992 -28450 3008
rect -34896 2912 -34769 2928
rect -34896 2848 -34849 2912
rect -34785 2848 -34769 2912
rect -34896 2832 -34769 2848
rect -34896 2768 -34849 2832
rect -34785 2768 -34769 2832
rect -34896 2752 -34769 2768
rect -34896 2688 -34849 2752
rect -34785 2688 -34769 2752
rect -34896 2672 -34769 2688
rect -34896 2608 -34849 2672
rect -34785 2608 -34769 2672
rect -34896 2592 -34769 2608
rect -34896 2528 -34849 2592
rect -34785 2528 -34769 2592
rect -34896 2512 -34769 2528
rect -34896 2448 -34849 2512
rect -34785 2448 -34769 2512
rect -34896 2432 -34769 2448
rect -34896 2368 -34849 2432
rect -34785 2368 -34769 2432
rect -34896 2352 -34769 2368
rect -34896 2288 -34849 2352
rect -34785 2288 -34769 2352
rect -34896 2272 -34769 2288
rect -34896 2208 -34849 2272
rect -34785 2208 -34769 2272
rect -34896 2192 -34769 2208
rect -34896 2128 -34849 2192
rect -34785 2128 -34769 2192
rect -34896 2112 -34769 2128
rect -34896 2048 -34849 2112
rect -34785 2048 -34769 2112
rect -34896 2032 -34769 2048
rect -34896 1968 -34849 2032
rect -34785 1968 -34769 2032
rect -34896 1952 -34769 1968
rect -34896 1888 -34849 1952
rect -34785 1888 -34769 1952
rect -34896 1872 -34769 1888
rect -34896 1808 -34849 1872
rect -34785 1808 -34769 1872
rect -34896 1792 -34769 1808
rect -34896 1728 -34849 1792
rect -34785 1728 -34769 1792
rect -34896 1712 -34769 1728
rect -34896 1648 -34849 1712
rect -34785 1648 -34769 1712
rect -34896 1632 -34769 1648
rect -34896 1568 -34849 1632
rect -34785 1568 -34769 1632
rect -34896 1552 -34769 1568
rect -34896 1488 -34849 1552
rect -34785 1488 -34769 1552
rect -34896 1472 -34769 1488
rect -34896 1408 -34849 1472
rect -34785 1408 -34769 1472
rect -34896 1392 -34769 1408
rect -34896 1328 -34849 1392
rect -34785 1328 -34769 1392
rect -34896 1312 -34769 1328
rect -34896 1248 -34849 1312
rect -34785 1248 -34769 1312
rect -34896 1232 -34769 1248
rect -34896 1168 -34849 1232
rect -34785 1168 -34769 1232
rect -34896 1152 -34769 1168
rect -34896 1088 -34849 1152
rect -34785 1088 -34769 1152
rect -34896 1072 -34769 1088
rect -34896 1008 -34849 1072
rect -34785 1008 -34769 1072
rect -34896 992 -34769 1008
rect -34896 928 -34849 992
rect -34785 928 -34769 992
rect -34896 912 -34769 928
rect -34896 848 -34849 912
rect -34785 848 -34769 912
rect -34896 832 -34769 848
rect -34896 768 -34849 832
rect -34785 768 -34769 832
rect -34896 752 -34769 768
rect -34896 688 -34849 752
rect -34785 688 -34769 752
rect -34896 672 -34769 688
rect -34896 608 -34849 672
rect -34785 608 -34769 672
rect -34896 592 -34769 608
rect -34896 528 -34849 592
rect -34785 528 -34769 592
rect -34896 512 -34769 528
rect -34896 448 -34849 512
rect -34785 448 -34769 512
rect -34896 432 -34769 448
rect -34896 368 -34849 432
rect -34785 368 -34769 432
rect -34896 352 -34769 368
rect -34896 288 -34849 352
rect -34785 288 -34769 352
rect -34896 272 -34769 288
rect -34896 208 -34849 272
rect -34785 208 -34769 272
rect -34896 192 -34769 208
rect -34896 128 -34849 192
rect -34785 128 -34769 192
rect -34896 112 -34769 128
rect -34896 48 -34849 112
rect -34785 48 -34769 112
rect -34896 32 -34769 48
rect -34896 -32 -34849 32
rect -34785 -32 -34769 32
rect -34896 -48 -34769 -32
rect -34896 -112 -34849 -48
rect -34785 -112 -34769 -48
rect -34896 -128 -34769 -112
rect -34896 -192 -34849 -128
rect -34785 -192 -34769 -128
rect -34896 -208 -34769 -192
rect -34896 -272 -34849 -208
rect -34785 -272 -34769 -208
rect -34896 -288 -34769 -272
rect -34896 -352 -34849 -288
rect -34785 -352 -34769 -288
rect -34896 -368 -34769 -352
rect -34896 -432 -34849 -368
rect -34785 -432 -34769 -368
rect -34896 -448 -34769 -432
rect -34896 -512 -34849 -448
rect -34785 -512 -34769 -448
rect -34896 -528 -34769 -512
rect -34896 -592 -34849 -528
rect -34785 -592 -34769 -528
rect -34896 -608 -34769 -592
rect -34896 -672 -34849 -608
rect -34785 -672 -34769 -608
rect -34896 -688 -34769 -672
rect -34896 -752 -34849 -688
rect -34785 -752 -34769 -688
rect -34896 -768 -34769 -752
rect -34896 -832 -34849 -768
rect -34785 -832 -34769 -768
rect -34896 -848 -34769 -832
rect -34896 -912 -34849 -848
rect -34785 -912 -34769 -848
rect -34896 -928 -34769 -912
rect -34896 -992 -34849 -928
rect -34785 -992 -34769 -928
rect -34896 -1008 -34769 -992
rect -34896 -1072 -34849 -1008
rect -34785 -1072 -34769 -1008
rect -34896 -1088 -34769 -1072
rect -34896 -1152 -34849 -1088
rect -34785 -1152 -34769 -1088
rect -34896 -1168 -34769 -1152
rect -34896 -1232 -34849 -1168
rect -34785 -1232 -34769 -1168
rect -34896 -1248 -34769 -1232
rect -34896 -1312 -34849 -1248
rect -34785 -1312 -34769 -1248
rect -34896 -1328 -34769 -1312
rect -34896 -1392 -34849 -1328
rect -34785 -1392 -34769 -1328
rect -34896 -1408 -34769 -1392
rect -34896 -1472 -34849 -1408
rect -34785 -1472 -34769 -1408
rect -34896 -1488 -34769 -1472
rect -34896 -1552 -34849 -1488
rect -34785 -1552 -34769 -1488
rect -34896 -1568 -34769 -1552
rect -34896 -1632 -34849 -1568
rect -34785 -1632 -34769 -1568
rect -34896 -1648 -34769 -1632
rect -34896 -1712 -34849 -1648
rect -34785 -1712 -34769 -1648
rect -34896 -1728 -34769 -1712
rect -34896 -1792 -34849 -1728
rect -34785 -1792 -34769 -1728
rect -34896 -1808 -34769 -1792
rect -34896 -1872 -34849 -1808
rect -34785 -1872 -34769 -1808
rect -34896 -1888 -34769 -1872
rect -34896 -1952 -34849 -1888
rect -34785 -1952 -34769 -1888
rect -34896 -1968 -34769 -1952
rect -34896 -2032 -34849 -1968
rect -34785 -2032 -34769 -1968
rect -34896 -2048 -34769 -2032
rect -34896 -2112 -34849 -2048
rect -34785 -2112 -34769 -2048
rect -34896 -2128 -34769 -2112
rect -34896 -2192 -34849 -2128
rect -34785 -2192 -34769 -2128
rect -34896 -2208 -34769 -2192
rect -34896 -2272 -34849 -2208
rect -34785 -2272 -34769 -2208
rect -34896 -2288 -34769 -2272
rect -34896 -2352 -34849 -2288
rect -34785 -2352 -34769 -2288
rect -34896 -2368 -34769 -2352
rect -34896 -2432 -34849 -2368
rect -34785 -2432 -34769 -2368
rect -34896 -2448 -34769 -2432
rect -34896 -2512 -34849 -2448
rect -34785 -2512 -34769 -2448
rect -34896 -2528 -34769 -2512
rect -34896 -2592 -34849 -2528
rect -34785 -2592 -34769 -2528
rect -34896 -2608 -34769 -2592
rect -34896 -2672 -34849 -2608
rect -34785 -2672 -34769 -2608
rect -34896 -2688 -34769 -2672
rect -34896 -2752 -34849 -2688
rect -34785 -2752 -34769 -2688
rect -34896 -2768 -34769 -2752
rect -34896 -2832 -34849 -2768
rect -34785 -2832 -34769 -2768
rect -34896 -2848 -34769 -2832
rect -34896 -2912 -34849 -2848
rect -34785 -2912 -34769 -2848
rect -34896 -2928 -34769 -2912
rect -41215 -3008 -41088 -2992
rect -41215 -3072 -41168 -3008
rect -41104 -3072 -41088 -3008
rect -41215 -3088 -41088 -3072
rect -41215 -3212 -41111 -3088
rect -41215 -3228 -41088 -3212
rect -41215 -3292 -41168 -3228
rect -41104 -3292 -41088 -3228
rect -41215 -3308 -41088 -3292
rect -47244 -3348 -41322 -3339
rect -47244 -9252 -47235 -3348
rect -41331 -9252 -41322 -3348
rect -47244 -9261 -41322 -9252
rect -41215 -3372 -41168 -3308
rect -41104 -3372 -41088 -3308
rect -38016 -3339 -37912 -2961
rect -34896 -2992 -34849 -2928
rect -34785 -2992 -34769 -2928
rect -34606 2952 -28684 2961
rect -34606 -2952 -34597 2952
rect -28693 -2952 -28684 2952
rect -34606 -2961 -28684 -2952
rect -28577 2928 -28530 2992
rect -28466 2928 -28450 2992
rect -25378 2961 -25274 3339
rect -22258 3308 -22211 3372
rect -22147 3308 -22131 3372
rect -21968 9252 -16046 9261
rect -21968 3348 -21959 9252
rect -16055 3348 -16046 9252
rect -21968 3339 -16046 3348
rect -15939 9228 -15892 9292
rect -15828 9228 -15812 9292
rect -12740 9261 -12636 9639
rect -9620 9608 -9573 9672
rect -9509 9608 -9493 9672
rect -9330 15552 -3408 15561
rect -9330 9648 -9321 15552
rect -3417 9648 -3408 15552
rect -9330 9639 -3408 9648
rect -3301 15528 -3254 15592
rect -3190 15528 -3174 15592
rect -102 15561 2 15939
rect 3018 15908 3065 15972
rect 3129 15908 3145 15972
rect 3308 21852 9230 21861
rect 3308 15948 3317 21852
rect 9221 15948 9230 21852
rect 3308 15939 9230 15948
rect 9337 21828 9384 21892
rect 9448 21828 9464 21892
rect 12536 21861 12640 22239
rect 15656 22208 15703 22272
rect 15767 22208 15783 22272
rect 15946 28152 21868 28161
rect 15946 22248 15955 28152
rect 21859 22248 21868 28152
rect 15946 22239 21868 22248
rect 21975 28128 22022 28192
rect 22086 28128 22102 28192
rect 25174 28161 25278 28539
rect 28294 28508 28341 28572
rect 28405 28508 28421 28572
rect 28584 34452 34506 34461
rect 28584 28548 28593 34452
rect 34497 28548 34506 34452
rect 28584 28539 34506 28548
rect 34613 34428 34660 34492
rect 34724 34428 34740 34492
rect 37812 34461 37916 34839
rect 40932 34808 40979 34872
rect 41043 34808 41059 34872
rect 41222 40752 47144 40761
rect 41222 34848 41231 40752
rect 47135 34848 47144 40752
rect 41222 34839 47144 34848
rect 47251 40728 47298 40792
rect 47362 40728 47378 40792
rect 47251 40712 47378 40728
rect 47251 40648 47298 40712
rect 47362 40648 47378 40712
rect 47251 40632 47378 40648
rect 47251 40568 47298 40632
rect 47362 40568 47378 40632
rect 47251 40552 47378 40568
rect 47251 40488 47298 40552
rect 47362 40488 47378 40552
rect 47251 40472 47378 40488
rect 47251 40408 47298 40472
rect 47362 40408 47378 40472
rect 47251 40392 47378 40408
rect 47251 40328 47298 40392
rect 47362 40328 47378 40392
rect 47251 40312 47378 40328
rect 47251 40248 47298 40312
rect 47362 40248 47378 40312
rect 47251 40232 47378 40248
rect 47251 40168 47298 40232
rect 47362 40168 47378 40232
rect 47251 40152 47378 40168
rect 47251 40088 47298 40152
rect 47362 40088 47378 40152
rect 47251 40072 47378 40088
rect 47251 40008 47298 40072
rect 47362 40008 47378 40072
rect 47251 39992 47378 40008
rect 47251 39928 47298 39992
rect 47362 39928 47378 39992
rect 47251 39912 47378 39928
rect 47251 39848 47298 39912
rect 47362 39848 47378 39912
rect 47251 39832 47378 39848
rect 47251 39768 47298 39832
rect 47362 39768 47378 39832
rect 47251 39752 47378 39768
rect 47251 39688 47298 39752
rect 47362 39688 47378 39752
rect 47251 39672 47378 39688
rect 47251 39608 47298 39672
rect 47362 39608 47378 39672
rect 47251 39592 47378 39608
rect 47251 39528 47298 39592
rect 47362 39528 47378 39592
rect 47251 39512 47378 39528
rect 47251 39448 47298 39512
rect 47362 39448 47378 39512
rect 47251 39432 47378 39448
rect 47251 39368 47298 39432
rect 47362 39368 47378 39432
rect 47251 39352 47378 39368
rect 47251 39288 47298 39352
rect 47362 39288 47378 39352
rect 47251 39272 47378 39288
rect 47251 39208 47298 39272
rect 47362 39208 47378 39272
rect 47251 39192 47378 39208
rect 47251 39128 47298 39192
rect 47362 39128 47378 39192
rect 47251 39112 47378 39128
rect 47251 39048 47298 39112
rect 47362 39048 47378 39112
rect 47251 39032 47378 39048
rect 47251 38968 47298 39032
rect 47362 38968 47378 39032
rect 47251 38952 47378 38968
rect 47251 38888 47298 38952
rect 47362 38888 47378 38952
rect 47251 38872 47378 38888
rect 47251 38808 47298 38872
rect 47362 38808 47378 38872
rect 47251 38792 47378 38808
rect 47251 38728 47298 38792
rect 47362 38728 47378 38792
rect 47251 38712 47378 38728
rect 47251 38648 47298 38712
rect 47362 38648 47378 38712
rect 47251 38632 47378 38648
rect 47251 38568 47298 38632
rect 47362 38568 47378 38632
rect 47251 38552 47378 38568
rect 47251 38488 47298 38552
rect 47362 38488 47378 38552
rect 47251 38472 47378 38488
rect 47251 38408 47298 38472
rect 47362 38408 47378 38472
rect 47251 38392 47378 38408
rect 47251 38328 47298 38392
rect 47362 38328 47378 38392
rect 47251 38312 47378 38328
rect 47251 38248 47298 38312
rect 47362 38248 47378 38312
rect 47251 38232 47378 38248
rect 47251 38168 47298 38232
rect 47362 38168 47378 38232
rect 47251 38152 47378 38168
rect 47251 38088 47298 38152
rect 47362 38088 47378 38152
rect 47251 38072 47378 38088
rect 47251 38008 47298 38072
rect 47362 38008 47378 38072
rect 47251 37992 47378 38008
rect 47251 37928 47298 37992
rect 47362 37928 47378 37992
rect 47251 37912 47378 37928
rect 47251 37848 47298 37912
rect 47362 37848 47378 37912
rect 47251 37832 47378 37848
rect 47251 37768 47298 37832
rect 47362 37768 47378 37832
rect 47251 37752 47378 37768
rect 47251 37688 47298 37752
rect 47362 37688 47378 37752
rect 47251 37672 47378 37688
rect 47251 37608 47298 37672
rect 47362 37608 47378 37672
rect 47251 37592 47378 37608
rect 47251 37528 47298 37592
rect 47362 37528 47378 37592
rect 47251 37512 47378 37528
rect 47251 37448 47298 37512
rect 47362 37448 47378 37512
rect 47251 37432 47378 37448
rect 47251 37368 47298 37432
rect 47362 37368 47378 37432
rect 47251 37352 47378 37368
rect 47251 37288 47298 37352
rect 47362 37288 47378 37352
rect 47251 37272 47378 37288
rect 47251 37208 47298 37272
rect 47362 37208 47378 37272
rect 47251 37192 47378 37208
rect 47251 37128 47298 37192
rect 47362 37128 47378 37192
rect 47251 37112 47378 37128
rect 47251 37048 47298 37112
rect 47362 37048 47378 37112
rect 47251 37032 47378 37048
rect 47251 36968 47298 37032
rect 47362 36968 47378 37032
rect 47251 36952 47378 36968
rect 47251 36888 47298 36952
rect 47362 36888 47378 36952
rect 47251 36872 47378 36888
rect 47251 36808 47298 36872
rect 47362 36808 47378 36872
rect 47251 36792 47378 36808
rect 47251 36728 47298 36792
rect 47362 36728 47378 36792
rect 47251 36712 47378 36728
rect 47251 36648 47298 36712
rect 47362 36648 47378 36712
rect 47251 36632 47378 36648
rect 47251 36568 47298 36632
rect 47362 36568 47378 36632
rect 47251 36552 47378 36568
rect 47251 36488 47298 36552
rect 47362 36488 47378 36552
rect 47251 36472 47378 36488
rect 47251 36408 47298 36472
rect 47362 36408 47378 36472
rect 47251 36392 47378 36408
rect 47251 36328 47298 36392
rect 47362 36328 47378 36392
rect 47251 36312 47378 36328
rect 47251 36248 47298 36312
rect 47362 36248 47378 36312
rect 47251 36232 47378 36248
rect 47251 36168 47298 36232
rect 47362 36168 47378 36232
rect 47251 36152 47378 36168
rect 47251 36088 47298 36152
rect 47362 36088 47378 36152
rect 47251 36072 47378 36088
rect 47251 36008 47298 36072
rect 47362 36008 47378 36072
rect 47251 35992 47378 36008
rect 47251 35928 47298 35992
rect 47362 35928 47378 35992
rect 47251 35912 47378 35928
rect 47251 35848 47298 35912
rect 47362 35848 47378 35912
rect 47251 35832 47378 35848
rect 47251 35768 47298 35832
rect 47362 35768 47378 35832
rect 47251 35752 47378 35768
rect 47251 35688 47298 35752
rect 47362 35688 47378 35752
rect 47251 35672 47378 35688
rect 47251 35608 47298 35672
rect 47362 35608 47378 35672
rect 47251 35592 47378 35608
rect 47251 35528 47298 35592
rect 47362 35528 47378 35592
rect 47251 35512 47378 35528
rect 47251 35448 47298 35512
rect 47362 35448 47378 35512
rect 47251 35432 47378 35448
rect 47251 35368 47298 35432
rect 47362 35368 47378 35432
rect 47251 35352 47378 35368
rect 47251 35288 47298 35352
rect 47362 35288 47378 35352
rect 47251 35272 47378 35288
rect 47251 35208 47298 35272
rect 47362 35208 47378 35272
rect 47251 35192 47378 35208
rect 47251 35128 47298 35192
rect 47362 35128 47378 35192
rect 47251 35112 47378 35128
rect 47251 35048 47298 35112
rect 47362 35048 47378 35112
rect 47251 35032 47378 35048
rect 47251 34968 47298 35032
rect 47362 34968 47378 35032
rect 47251 34952 47378 34968
rect 47251 34888 47298 34952
rect 47362 34888 47378 34952
rect 47251 34872 47378 34888
rect 40932 34792 41059 34808
rect 40932 34728 40979 34792
rect 41043 34728 41059 34792
rect 40932 34712 41059 34728
rect 40932 34588 41036 34712
rect 40932 34572 41059 34588
rect 40932 34508 40979 34572
rect 41043 34508 41059 34572
rect 40932 34492 41059 34508
rect 34613 34412 34740 34428
rect 34613 34348 34660 34412
rect 34724 34348 34740 34412
rect 34613 34332 34740 34348
rect 34613 34268 34660 34332
rect 34724 34268 34740 34332
rect 34613 34252 34740 34268
rect 34613 34188 34660 34252
rect 34724 34188 34740 34252
rect 34613 34172 34740 34188
rect 34613 34108 34660 34172
rect 34724 34108 34740 34172
rect 34613 34092 34740 34108
rect 34613 34028 34660 34092
rect 34724 34028 34740 34092
rect 34613 34012 34740 34028
rect 34613 33948 34660 34012
rect 34724 33948 34740 34012
rect 34613 33932 34740 33948
rect 34613 33868 34660 33932
rect 34724 33868 34740 33932
rect 34613 33852 34740 33868
rect 34613 33788 34660 33852
rect 34724 33788 34740 33852
rect 34613 33772 34740 33788
rect 34613 33708 34660 33772
rect 34724 33708 34740 33772
rect 34613 33692 34740 33708
rect 34613 33628 34660 33692
rect 34724 33628 34740 33692
rect 34613 33612 34740 33628
rect 34613 33548 34660 33612
rect 34724 33548 34740 33612
rect 34613 33532 34740 33548
rect 34613 33468 34660 33532
rect 34724 33468 34740 33532
rect 34613 33452 34740 33468
rect 34613 33388 34660 33452
rect 34724 33388 34740 33452
rect 34613 33372 34740 33388
rect 34613 33308 34660 33372
rect 34724 33308 34740 33372
rect 34613 33292 34740 33308
rect 34613 33228 34660 33292
rect 34724 33228 34740 33292
rect 34613 33212 34740 33228
rect 34613 33148 34660 33212
rect 34724 33148 34740 33212
rect 34613 33132 34740 33148
rect 34613 33068 34660 33132
rect 34724 33068 34740 33132
rect 34613 33052 34740 33068
rect 34613 32988 34660 33052
rect 34724 32988 34740 33052
rect 34613 32972 34740 32988
rect 34613 32908 34660 32972
rect 34724 32908 34740 32972
rect 34613 32892 34740 32908
rect 34613 32828 34660 32892
rect 34724 32828 34740 32892
rect 34613 32812 34740 32828
rect 34613 32748 34660 32812
rect 34724 32748 34740 32812
rect 34613 32732 34740 32748
rect 34613 32668 34660 32732
rect 34724 32668 34740 32732
rect 34613 32652 34740 32668
rect 34613 32588 34660 32652
rect 34724 32588 34740 32652
rect 34613 32572 34740 32588
rect 34613 32508 34660 32572
rect 34724 32508 34740 32572
rect 34613 32492 34740 32508
rect 34613 32428 34660 32492
rect 34724 32428 34740 32492
rect 34613 32412 34740 32428
rect 34613 32348 34660 32412
rect 34724 32348 34740 32412
rect 34613 32332 34740 32348
rect 34613 32268 34660 32332
rect 34724 32268 34740 32332
rect 34613 32252 34740 32268
rect 34613 32188 34660 32252
rect 34724 32188 34740 32252
rect 34613 32172 34740 32188
rect 34613 32108 34660 32172
rect 34724 32108 34740 32172
rect 34613 32092 34740 32108
rect 34613 32028 34660 32092
rect 34724 32028 34740 32092
rect 34613 32012 34740 32028
rect 34613 31948 34660 32012
rect 34724 31948 34740 32012
rect 34613 31932 34740 31948
rect 34613 31868 34660 31932
rect 34724 31868 34740 31932
rect 34613 31852 34740 31868
rect 34613 31788 34660 31852
rect 34724 31788 34740 31852
rect 34613 31772 34740 31788
rect 34613 31708 34660 31772
rect 34724 31708 34740 31772
rect 34613 31692 34740 31708
rect 34613 31628 34660 31692
rect 34724 31628 34740 31692
rect 34613 31612 34740 31628
rect 34613 31548 34660 31612
rect 34724 31548 34740 31612
rect 34613 31532 34740 31548
rect 34613 31468 34660 31532
rect 34724 31468 34740 31532
rect 34613 31452 34740 31468
rect 34613 31388 34660 31452
rect 34724 31388 34740 31452
rect 34613 31372 34740 31388
rect 34613 31308 34660 31372
rect 34724 31308 34740 31372
rect 34613 31292 34740 31308
rect 34613 31228 34660 31292
rect 34724 31228 34740 31292
rect 34613 31212 34740 31228
rect 34613 31148 34660 31212
rect 34724 31148 34740 31212
rect 34613 31132 34740 31148
rect 34613 31068 34660 31132
rect 34724 31068 34740 31132
rect 34613 31052 34740 31068
rect 34613 30988 34660 31052
rect 34724 30988 34740 31052
rect 34613 30972 34740 30988
rect 34613 30908 34660 30972
rect 34724 30908 34740 30972
rect 34613 30892 34740 30908
rect 34613 30828 34660 30892
rect 34724 30828 34740 30892
rect 34613 30812 34740 30828
rect 34613 30748 34660 30812
rect 34724 30748 34740 30812
rect 34613 30732 34740 30748
rect 34613 30668 34660 30732
rect 34724 30668 34740 30732
rect 34613 30652 34740 30668
rect 34613 30588 34660 30652
rect 34724 30588 34740 30652
rect 34613 30572 34740 30588
rect 34613 30508 34660 30572
rect 34724 30508 34740 30572
rect 34613 30492 34740 30508
rect 34613 30428 34660 30492
rect 34724 30428 34740 30492
rect 34613 30412 34740 30428
rect 34613 30348 34660 30412
rect 34724 30348 34740 30412
rect 34613 30332 34740 30348
rect 34613 30268 34660 30332
rect 34724 30268 34740 30332
rect 34613 30252 34740 30268
rect 34613 30188 34660 30252
rect 34724 30188 34740 30252
rect 34613 30172 34740 30188
rect 34613 30108 34660 30172
rect 34724 30108 34740 30172
rect 34613 30092 34740 30108
rect 34613 30028 34660 30092
rect 34724 30028 34740 30092
rect 34613 30012 34740 30028
rect 34613 29948 34660 30012
rect 34724 29948 34740 30012
rect 34613 29932 34740 29948
rect 34613 29868 34660 29932
rect 34724 29868 34740 29932
rect 34613 29852 34740 29868
rect 34613 29788 34660 29852
rect 34724 29788 34740 29852
rect 34613 29772 34740 29788
rect 34613 29708 34660 29772
rect 34724 29708 34740 29772
rect 34613 29692 34740 29708
rect 34613 29628 34660 29692
rect 34724 29628 34740 29692
rect 34613 29612 34740 29628
rect 34613 29548 34660 29612
rect 34724 29548 34740 29612
rect 34613 29532 34740 29548
rect 34613 29468 34660 29532
rect 34724 29468 34740 29532
rect 34613 29452 34740 29468
rect 34613 29388 34660 29452
rect 34724 29388 34740 29452
rect 34613 29372 34740 29388
rect 34613 29308 34660 29372
rect 34724 29308 34740 29372
rect 34613 29292 34740 29308
rect 34613 29228 34660 29292
rect 34724 29228 34740 29292
rect 34613 29212 34740 29228
rect 34613 29148 34660 29212
rect 34724 29148 34740 29212
rect 34613 29132 34740 29148
rect 34613 29068 34660 29132
rect 34724 29068 34740 29132
rect 34613 29052 34740 29068
rect 34613 28988 34660 29052
rect 34724 28988 34740 29052
rect 34613 28972 34740 28988
rect 34613 28908 34660 28972
rect 34724 28908 34740 28972
rect 34613 28892 34740 28908
rect 34613 28828 34660 28892
rect 34724 28828 34740 28892
rect 34613 28812 34740 28828
rect 34613 28748 34660 28812
rect 34724 28748 34740 28812
rect 34613 28732 34740 28748
rect 34613 28668 34660 28732
rect 34724 28668 34740 28732
rect 34613 28652 34740 28668
rect 34613 28588 34660 28652
rect 34724 28588 34740 28652
rect 34613 28572 34740 28588
rect 28294 28492 28421 28508
rect 28294 28428 28341 28492
rect 28405 28428 28421 28492
rect 28294 28412 28421 28428
rect 28294 28288 28398 28412
rect 28294 28272 28421 28288
rect 28294 28208 28341 28272
rect 28405 28208 28421 28272
rect 28294 28192 28421 28208
rect 21975 28112 22102 28128
rect 21975 28048 22022 28112
rect 22086 28048 22102 28112
rect 21975 28032 22102 28048
rect 21975 27968 22022 28032
rect 22086 27968 22102 28032
rect 21975 27952 22102 27968
rect 21975 27888 22022 27952
rect 22086 27888 22102 27952
rect 21975 27872 22102 27888
rect 21975 27808 22022 27872
rect 22086 27808 22102 27872
rect 21975 27792 22102 27808
rect 21975 27728 22022 27792
rect 22086 27728 22102 27792
rect 21975 27712 22102 27728
rect 21975 27648 22022 27712
rect 22086 27648 22102 27712
rect 21975 27632 22102 27648
rect 21975 27568 22022 27632
rect 22086 27568 22102 27632
rect 21975 27552 22102 27568
rect 21975 27488 22022 27552
rect 22086 27488 22102 27552
rect 21975 27472 22102 27488
rect 21975 27408 22022 27472
rect 22086 27408 22102 27472
rect 21975 27392 22102 27408
rect 21975 27328 22022 27392
rect 22086 27328 22102 27392
rect 21975 27312 22102 27328
rect 21975 27248 22022 27312
rect 22086 27248 22102 27312
rect 21975 27232 22102 27248
rect 21975 27168 22022 27232
rect 22086 27168 22102 27232
rect 21975 27152 22102 27168
rect 21975 27088 22022 27152
rect 22086 27088 22102 27152
rect 21975 27072 22102 27088
rect 21975 27008 22022 27072
rect 22086 27008 22102 27072
rect 21975 26992 22102 27008
rect 21975 26928 22022 26992
rect 22086 26928 22102 26992
rect 21975 26912 22102 26928
rect 21975 26848 22022 26912
rect 22086 26848 22102 26912
rect 21975 26832 22102 26848
rect 21975 26768 22022 26832
rect 22086 26768 22102 26832
rect 21975 26752 22102 26768
rect 21975 26688 22022 26752
rect 22086 26688 22102 26752
rect 21975 26672 22102 26688
rect 21975 26608 22022 26672
rect 22086 26608 22102 26672
rect 21975 26592 22102 26608
rect 21975 26528 22022 26592
rect 22086 26528 22102 26592
rect 21975 26512 22102 26528
rect 21975 26448 22022 26512
rect 22086 26448 22102 26512
rect 21975 26432 22102 26448
rect 21975 26368 22022 26432
rect 22086 26368 22102 26432
rect 21975 26352 22102 26368
rect 21975 26288 22022 26352
rect 22086 26288 22102 26352
rect 21975 26272 22102 26288
rect 21975 26208 22022 26272
rect 22086 26208 22102 26272
rect 21975 26192 22102 26208
rect 21975 26128 22022 26192
rect 22086 26128 22102 26192
rect 21975 26112 22102 26128
rect 21975 26048 22022 26112
rect 22086 26048 22102 26112
rect 21975 26032 22102 26048
rect 21975 25968 22022 26032
rect 22086 25968 22102 26032
rect 21975 25952 22102 25968
rect 21975 25888 22022 25952
rect 22086 25888 22102 25952
rect 21975 25872 22102 25888
rect 21975 25808 22022 25872
rect 22086 25808 22102 25872
rect 21975 25792 22102 25808
rect 21975 25728 22022 25792
rect 22086 25728 22102 25792
rect 21975 25712 22102 25728
rect 21975 25648 22022 25712
rect 22086 25648 22102 25712
rect 21975 25632 22102 25648
rect 21975 25568 22022 25632
rect 22086 25568 22102 25632
rect 21975 25552 22102 25568
rect 21975 25488 22022 25552
rect 22086 25488 22102 25552
rect 21975 25472 22102 25488
rect 21975 25408 22022 25472
rect 22086 25408 22102 25472
rect 21975 25392 22102 25408
rect 21975 25328 22022 25392
rect 22086 25328 22102 25392
rect 21975 25312 22102 25328
rect 21975 25248 22022 25312
rect 22086 25248 22102 25312
rect 21975 25232 22102 25248
rect 21975 25168 22022 25232
rect 22086 25168 22102 25232
rect 21975 25152 22102 25168
rect 21975 25088 22022 25152
rect 22086 25088 22102 25152
rect 21975 25072 22102 25088
rect 21975 25008 22022 25072
rect 22086 25008 22102 25072
rect 21975 24992 22102 25008
rect 21975 24928 22022 24992
rect 22086 24928 22102 24992
rect 21975 24912 22102 24928
rect 21975 24848 22022 24912
rect 22086 24848 22102 24912
rect 21975 24832 22102 24848
rect 21975 24768 22022 24832
rect 22086 24768 22102 24832
rect 21975 24752 22102 24768
rect 21975 24688 22022 24752
rect 22086 24688 22102 24752
rect 21975 24672 22102 24688
rect 21975 24608 22022 24672
rect 22086 24608 22102 24672
rect 21975 24592 22102 24608
rect 21975 24528 22022 24592
rect 22086 24528 22102 24592
rect 21975 24512 22102 24528
rect 21975 24448 22022 24512
rect 22086 24448 22102 24512
rect 21975 24432 22102 24448
rect 21975 24368 22022 24432
rect 22086 24368 22102 24432
rect 21975 24352 22102 24368
rect 21975 24288 22022 24352
rect 22086 24288 22102 24352
rect 21975 24272 22102 24288
rect 21975 24208 22022 24272
rect 22086 24208 22102 24272
rect 21975 24192 22102 24208
rect 21975 24128 22022 24192
rect 22086 24128 22102 24192
rect 21975 24112 22102 24128
rect 21975 24048 22022 24112
rect 22086 24048 22102 24112
rect 21975 24032 22102 24048
rect 21975 23968 22022 24032
rect 22086 23968 22102 24032
rect 21975 23952 22102 23968
rect 21975 23888 22022 23952
rect 22086 23888 22102 23952
rect 21975 23872 22102 23888
rect 21975 23808 22022 23872
rect 22086 23808 22102 23872
rect 21975 23792 22102 23808
rect 21975 23728 22022 23792
rect 22086 23728 22102 23792
rect 21975 23712 22102 23728
rect 21975 23648 22022 23712
rect 22086 23648 22102 23712
rect 21975 23632 22102 23648
rect 21975 23568 22022 23632
rect 22086 23568 22102 23632
rect 21975 23552 22102 23568
rect 21975 23488 22022 23552
rect 22086 23488 22102 23552
rect 21975 23472 22102 23488
rect 21975 23408 22022 23472
rect 22086 23408 22102 23472
rect 21975 23392 22102 23408
rect 21975 23328 22022 23392
rect 22086 23328 22102 23392
rect 21975 23312 22102 23328
rect 21975 23248 22022 23312
rect 22086 23248 22102 23312
rect 21975 23232 22102 23248
rect 21975 23168 22022 23232
rect 22086 23168 22102 23232
rect 21975 23152 22102 23168
rect 21975 23088 22022 23152
rect 22086 23088 22102 23152
rect 21975 23072 22102 23088
rect 21975 23008 22022 23072
rect 22086 23008 22102 23072
rect 21975 22992 22102 23008
rect 21975 22928 22022 22992
rect 22086 22928 22102 22992
rect 21975 22912 22102 22928
rect 21975 22848 22022 22912
rect 22086 22848 22102 22912
rect 21975 22832 22102 22848
rect 21975 22768 22022 22832
rect 22086 22768 22102 22832
rect 21975 22752 22102 22768
rect 21975 22688 22022 22752
rect 22086 22688 22102 22752
rect 21975 22672 22102 22688
rect 21975 22608 22022 22672
rect 22086 22608 22102 22672
rect 21975 22592 22102 22608
rect 21975 22528 22022 22592
rect 22086 22528 22102 22592
rect 21975 22512 22102 22528
rect 21975 22448 22022 22512
rect 22086 22448 22102 22512
rect 21975 22432 22102 22448
rect 21975 22368 22022 22432
rect 22086 22368 22102 22432
rect 21975 22352 22102 22368
rect 21975 22288 22022 22352
rect 22086 22288 22102 22352
rect 21975 22272 22102 22288
rect 15656 22192 15783 22208
rect 15656 22128 15703 22192
rect 15767 22128 15783 22192
rect 15656 22112 15783 22128
rect 15656 21988 15760 22112
rect 15656 21972 15783 21988
rect 15656 21908 15703 21972
rect 15767 21908 15783 21972
rect 15656 21892 15783 21908
rect 9337 21812 9464 21828
rect 9337 21748 9384 21812
rect 9448 21748 9464 21812
rect 9337 21732 9464 21748
rect 9337 21668 9384 21732
rect 9448 21668 9464 21732
rect 9337 21652 9464 21668
rect 9337 21588 9384 21652
rect 9448 21588 9464 21652
rect 9337 21572 9464 21588
rect 9337 21508 9384 21572
rect 9448 21508 9464 21572
rect 9337 21492 9464 21508
rect 9337 21428 9384 21492
rect 9448 21428 9464 21492
rect 9337 21412 9464 21428
rect 9337 21348 9384 21412
rect 9448 21348 9464 21412
rect 9337 21332 9464 21348
rect 9337 21268 9384 21332
rect 9448 21268 9464 21332
rect 9337 21252 9464 21268
rect 9337 21188 9384 21252
rect 9448 21188 9464 21252
rect 9337 21172 9464 21188
rect 9337 21108 9384 21172
rect 9448 21108 9464 21172
rect 9337 21092 9464 21108
rect 9337 21028 9384 21092
rect 9448 21028 9464 21092
rect 9337 21012 9464 21028
rect 9337 20948 9384 21012
rect 9448 20948 9464 21012
rect 9337 20932 9464 20948
rect 9337 20868 9384 20932
rect 9448 20868 9464 20932
rect 9337 20852 9464 20868
rect 9337 20788 9384 20852
rect 9448 20788 9464 20852
rect 9337 20772 9464 20788
rect 9337 20708 9384 20772
rect 9448 20708 9464 20772
rect 9337 20692 9464 20708
rect 9337 20628 9384 20692
rect 9448 20628 9464 20692
rect 9337 20612 9464 20628
rect 9337 20548 9384 20612
rect 9448 20548 9464 20612
rect 9337 20532 9464 20548
rect 9337 20468 9384 20532
rect 9448 20468 9464 20532
rect 9337 20452 9464 20468
rect 9337 20388 9384 20452
rect 9448 20388 9464 20452
rect 9337 20372 9464 20388
rect 9337 20308 9384 20372
rect 9448 20308 9464 20372
rect 9337 20292 9464 20308
rect 9337 20228 9384 20292
rect 9448 20228 9464 20292
rect 9337 20212 9464 20228
rect 9337 20148 9384 20212
rect 9448 20148 9464 20212
rect 9337 20132 9464 20148
rect 9337 20068 9384 20132
rect 9448 20068 9464 20132
rect 9337 20052 9464 20068
rect 9337 19988 9384 20052
rect 9448 19988 9464 20052
rect 9337 19972 9464 19988
rect 9337 19908 9384 19972
rect 9448 19908 9464 19972
rect 9337 19892 9464 19908
rect 9337 19828 9384 19892
rect 9448 19828 9464 19892
rect 9337 19812 9464 19828
rect 9337 19748 9384 19812
rect 9448 19748 9464 19812
rect 9337 19732 9464 19748
rect 9337 19668 9384 19732
rect 9448 19668 9464 19732
rect 9337 19652 9464 19668
rect 9337 19588 9384 19652
rect 9448 19588 9464 19652
rect 9337 19572 9464 19588
rect 9337 19508 9384 19572
rect 9448 19508 9464 19572
rect 9337 19492 9464 19508
rect 9337 19428 9384 19492
rect 9448 19428 9464 19492
rect 9337 19412 9464 19428
rect 9337 19348 9384 19412
rect 9448 19348 9464 19412
rect 9337 19332 9464 19348
rect 9337 19268 9384 19332
rect 9448 19268 9464 19332
rect 9337 19252 9464 19268
rect 9337 19188 9384 19252
rect 9448 19188 9464 19252
rect 9337 19172 9464 19188
rect 9337 19108 9384 19172
rect 9448 19108 9464 19172
rect 9337 19092 9464 19108
rect 9337 19028 9384 19092
rect 9448 19028 9464 19092
rect 9337 19012 9464 19028
rect 9337 18948 9384 19012
rect 9448 18948 9464 19012
rect 9337 18932 9464 18948
rect 9337 18868 9384 18932
rect 9448 18868 9464 18932
rect 9337 18852 9464 18868
rect 9337 18788 9384 18852
rect 9448 18788 9464 18852
rect 9337 18772 9464 18788
rect 9337 18708 9384 18772
rect 9448 18708 9464 18772
rect 9337 18692 9464 18708
rect 9337 18628 9384 18692
rect 9448 18628 9464 18692
rect 9337 18612 9464 18628
rect 9337 18548 9384 18612
rect 9448 18548 9464 18612
rect 9337 18532 9464 18548
rect 9337 18468 9384 18532
rect 9448 18468 9464 18532
rect 9337 18452 9464 18468
rect 9337 18388 9384 18452
rect 9448 18388 9464 18452
rect 9337 18372 9464 18388
rect 9337 18308 9384 18372
rect 9448 18308 9464 18372
rect 9337 18292 9464 18308
rect 9337 18228 9384 18292
rect 9448 18228 9464 18292
rect 9337 18212 9464 18228
rect 9337 18148 9384 18212
rect 9448 18148 9464 18212
rect 9337 18132 9464 18148
rect 9337 18068 9384 18132
rect 9448 18068 9464 18132
rect 9337 18052 9464 18068
rect 9337 17988 9384 18052
rect 9448 17988 9464 18052
rect 9337 17972 9464 17988
rect 9337 17908 9384 17972
rect 9448 17908 9464 17972
rect 9337 17892 9464 17908
rect 9337 17828 9384 17892
rect 9448 17828 9464 17892
rect 9337 17812 9464 17828
rect 9337 17748 9384 17812
rect 9448 17748 9464 17812
rect 9337 17732 9464 17748
rect 9337 17668 9384 17732
rect 9448 17668 9464 17732
rect 9337 17652 9464 17668
rect 9337 17588 9384 17652
rect 9448 17588 9464 17652
rect 9337 17572 9464 17588
rect 9337 17508 9384 17572
rect 9448 17508 9464 17572
rect 9337 17492 9464 17508
rect 9337 17428 9384 17492
rect 9448 17428 9464 17492
rect 9337 17412 9464 17428
rect 9337 17348 9384 17412
rect 9448 17348 9464 17412
rect 9337 17332 9464 17348
rect 9337 17268 9384 17332
rect 9448 17268 9464 17332
rect 9337 17252 9464 17268
rect 9337 17188 9384 17252
rect 9448 17188 9464 17252
rect 9337 17172 9464 17188
rect 9337 17108 9384 17172
rect 9448 17108 9464 17172
rect 9337 17092 9464 17108
rect 9337 17028 9384 17092
rect 9448 17028 9464 17092
rect 9337 17012 9464 17028
rect 9337 16948 9384 17012
rect 9448 16948 9464 17012
rect 9337 16932 9464 16948
rect 9337 16868 9384 16932
rect 9448 16868 9464 16932
rect 9337 16852 9464 16868
rect 9337 16788 9384 16852
rect 9448 16788 9464 16852
rect 9337 16772 9464 16788
rect 9337 16708 9384 16772
rect 9448 16708 9464 16772
rect 9337 16692 9464 16708
rect 9337 16628 9384 16692
rect 9448 16628 9464 16692
rect 9337 16612 9464 16628
rect 9337 16548 9384 16612
rect 9448 16548 9464 16612
rect 9337 16532 9464 16548
rect 9337 16468 9384 16532
rect 9448 16468 9464 16532
rect 9337 16452 9464 16468
rect 9337 16388 9384 16452
rect 9448 16388 9464 16452
rect 9337 16372 9464 16388
rect 9337 16308 9384 16372
rect 9448 16308 9464 16372
rect 9337 16292 9464 16308
rect 9337 16228 9384 16292
rect 9448 16228 9464 16292
rect 9337 16212 9464 16228
rect 9337 16148 9384 16212
rect 9448 16148 9464 16212
rect 9337 16132 9464 16148
rect 9337 16068 9384 16132
rect 9448 16068 9464 16132
rect 9337 16052 9464 16068
rect 9337 15988 9384 16052
rect 9448 15988 9464 16052
rect 9337 15972 9464 15988
rect 3018 15892 3145 15908
rect 3018 15828 3065 15892
rect 3129 15828 3145 15892
rect 3018 15812 3145 15828
rect 3018 15688 3122 15812
rect 3018 15672 3145 15688
rect 3018 15608 3065 15672
rect 3129 15608 3145 15672
rect 3018 15592 3145 15608
rect -3301 15512 -3174 15528
rect -3301 15448 -3254 15512
rect -3190 15448 -3174 15512
rect -3301 15432 -3174 15448
rect -3301 15368 -3254 15432
rect -3190 15368 -3174 15432
rect -3301 15352 -3174 15368
rect -3301 15288 -3254 15352
rect -3190 15288 -3174 15352
rect -3301 15272 -3174 15288
rect -3301 15208 -3254 15272
rect -3190 15208 -3174 15272
rect -3301 15192 -3174 15208
rect -3301 15128 -3254 15192
rect -3190 15128 -3174 15192
rect -3301 15112 -3174 15128
rect -3301 15048 -3254 15112
rect -3190 15048 -3174 15112
rect -3301 15032 -3174 15048
rect -3301 14968 -3254 15032
rect -3190 14968 -3174 15032
rect -3301 14952 -3174 14968
rect -3301 14888 -3254 14952
rect -3190 14888 -3174 14952
rect -3301 14872 -3174 14888
rect -3301 14808 -3254 14872
rect -3190 14808 -3174 14872
rect -3301 14792 -3174 14808
rect -3301 14728 -3254 14792
rect -3190 14728 -3174 14792
rect -3301 14712 -3174 14728
rect -3301 14648 -3254 14712
rect -3190 14648 -3174 14712
rect -3301 14632 -3174 14648
rect -3301 14568 -3254 14632
rect -3190 14568 -3174 14632
rect -3301 14552 -3174 14568
rect -3301 14488 -3254 14552
rect -3190 14488 -3174 14552
rect -3301 14472 -3174 14488
rect -3301 14408 -3254 14472
rect -3190 14408 -3174 14472
rect -3301 14392 -3174 14408
rect -3301 14328 -3254 14392
rect -3190 14328 -3174 14392
rect -3301 14312 -3174 14328
rect -3301 14248 -3254 14312
rect -3190 14248 -3174 14312
rect -3301 14232 -3174 14248
rect -3301 14168 -3254 14232
rect -3190 14168 -3174 14232
rect -3301 14152 -3174 14168
rect -3301 14088 -3254 14152
rect -3190 14088 -3174 14152
rect -3301 14072 -3174 14088
rect -3301 14008 -3254 14072
rect -3190 14008 -3174 14072
rect -3301 13992 -3174 14008
rect -3301 13928 -3254 13992
rect -3190 13928 -3174 13992
rect -3301 13912 -3174 13928
rect -3301 13848 -3254 13912
rect -3190 13848 -3174 13912
rect -3301 13832 -3174 13848
rect -3301 13768 -3254 13832
rect -3190 13768 -3174 13832
rect -3301 13752 -3174 13768
rect -3301 13688 -3254 13752
rect -3190 13688 -3174 13752
rect -3301 13672 -3174 13688
rect -3301 13608 -3254 13672
rect -3190 13608 -3174 13672
rect -3301 13592 -3174 13608
rect -3301 13528 -3254 13592
rect -3190 13528 -3174 13592
rect -3301 13512 -3174 13528
rect -3301 13448 -3254 13512
rect -3190 13448 -3174 13512
rect -3301 13432 -3174 13448
rect -3301 13368 -3254 13432
rect -3190 13368 -3174 13432
rect -3301 13352 -3174 13368
rect -3301 13288 -3254 13352
rect -3190 13288 -3174 13352
rect -3301 13272 -3174 13288
rect -3301 13208 -3254 13272
rect -3190 13208 -3174 13272
rect -3301 13192 -3174 13208
rect -3301 13128 -3254 13192
rect -3190 13128 -3174 13192
rect -3301 13112 -3174 13128
rect -3301 13048 -3254 13112
rect -3190 13048 -3174 13112
rect -3301 13032 -3174 13048
rect -3301 12968 -3254 13032
rect -3190 12968 -3174 13032
rect -3301 12952 -3174 12968
rect -3301 12888 -3254 12952
rect -3190 12888 -3174 12952
rect -3301 12872 -3174 12888
rect -3301 12808 -3254 12872
rect -3190 12808 -3174 12872
rect -3301 12792 -3174 12808
rect -3301 12728 -3254 12792
rect -3190 12728 -3174 12792
rect -3301 12712 -3174 12728
rect -3301 12648 -3254 12712
rect -3190 12648 -3174 12712
rect -3301 12632 -3174 12648
rect -3301 12568 -3254 12632
rect -3190 12568 -3174 12632
rect -3301 12552 -3174 12568
rect -3301 12488 -3254 12552
rect -3190 12488 -3174 12552
rect -3301 12472 -3174 12488
rect -3301 12408 -3254 12472
rect -3190 12408 -3174 12472
rect -3301 12392 -3174 12408
rect -3301 12328 -3254 12392
rect -3190 12328 -3174 12392
rect -3301 12312 -3174 12328
rect -3301 12248 -3254 12312
rect -3190 12248 -3174 12312
rect -3301 12232 -3174 12248
rect -3301 12168 -3254 12232
rect -3190 12168 -3174 12232
rect -3301 12152 -3174 12168
rect -3301 12088 -3254 12152
rect -3190 12088 -3174 12152
rect -3301 12072 -3174 12088
rect -3301 12008 -3254 12072
rect -3190 12008 -3174 12072
rect -3301 11992 -3174 12008
rect -3301 11928 -3254 11992
rect -3190 11928 -3174 11992
rect -3301 11912 -3174 11928
rect -3301 11848 -3254 11912
rect -3190 11848 -3174 11912
rect -3301 11832 -3174 11848
rect -3301 11768 -3254 11832
rect -3190 11768 -3174 11832
rect -3301 11752 -3174 11768
rect -3301 11688 -3254 11752
rect -3190 11688 -3174 11752
rect -3301 11672 -3174 11688
rect -3301 11608 -3254 11672
rect -3190 11608 -3174 11672
rect -3301 11592 -3174 11608
rect -3301 11528 -3254 11592
rect -3190 11528 -3174 11592
rect -3301 11512 -3174 11528
rect -3301 11448 -3254 11512
rect -3190 11448 -3174 11512
rect -3301 11432 -3174 11448
rect -3301 11368 -3254 11432
rect -3190 11368 -3174 11432
rect -3301 11352 -3174 11368
rect -3301 11288 -3254 11352
rect -3190 11288 -3174 11352
rect -3301 11272 -3174 11288
rect -3301 11208 -3254 11272
rect -3190 11208 -3174 11272
rect -3301 11192 -3174 11208
rect -3301 11128 -3254 11192
rect -3190 11128 -3174 11192
rect -3301 11112 -3174 11128
rect -3301 11048 -3254 11112
rect -3190 11048 -3174 11112
rect -3301 11032 -3174 11048
rect -3301 10968 -3254 11032
rect -3190 10968 -3174 11032
rect -3301 10952 -3174 10968
rect -3301 10888 -3254 10952
rect -3190 10888 -3174 10952
rect -3301 10872 -3174 10888
rect -3301 10808 -3254 10872
rect -3190 10808 -3174 10872
rect -3301 10792 -3174 10808
rect -3301 10728 -3254 10792
rect -3190 10728 -3174 10792
rect -3301 10712 -3174 10728
rect -3301 10648 -3254 10712
rect -3190 10648 -3174 10712
rect -3301 10632 -3174 10648
rect -3301 10568 -3254 10632
rect -3190 10568 -3174 10632
rect -3301 10552 -3174 10568
rect -3301 10488 -3254 10552
rect -3190 10488 -3174 10552
rect -3301 10472 -3174 10488
rect -3301 10408 -3254 10472
rect -3190 10408 -3174 10472
rect -3301 10392 -3174 10408
rect -3301 10328 -3254 10392
rect -3190 10328 -3174 10392
rect -3301 10312 -3174 10328
rect -3301 10248 -3254 10312
rect -3190 10248 -3174 10312
rect -3301 10232 -3174 10248
rect -3301 10168 -3254 10232
rect -3190 10168 -3174 10232
rect -3301 10152 -3174 10168
rect -3301 10088 -3254 10152
rect -3190 10088 -3174 10152
rect -3301 10072 -3174 10088
rect -3301 10008 -3254 10072
rect -3190 10008 -3174 10072
rect -3301 9992 -3174 10008
rect -3301 9928 -3254 9992
rect -3190 9928 -3174 9992
rect -3301 9912 -3174 9928
rect -3301 9848 -3254 9912
rect -3190 9848 -3174 9912
rect -3301 9832 -3174 9848
rect -3301 9768 -3254 9832
rect -3190 9768 -3174 9832
rect -3301 9752 -3174 9768
rect -3301 9688 -3254 9752
rect -3190 9688 -3174 9752
rect -3301 9672 -3174 9688
rect -9620 9592 -9493 9608
rect -9620 9528 -9573 9592
rect -9509 9528 -9493 9592
rect -9620 9512 -9493 9528
rect -9620 9388 -9516 9512
rect -9620 9372 -9493 9388
rect -9620 9308 -9573 9372
rect -9509 9308 -9493 9372
rect -9620 9292 -9493 9308
rect -15939 9212 -15812 9228
rect -15939 9148 -15892 9212
rect -15828 9148 -15812 9212
rect -15939 9132 -15812 9148
rect -15939 9068 -15892 9132
rect -15828 9068 -15812 9132
rect -15939 9052 -15812 9068
rect -15939 8988 -15892 9052
rect -15828 8988 -15812 9052
rect -15939 8972 -15812 8988
rect -15939 8908 -15892 8972
rect -15828 8908 -15812 8972
rect -15939 8892 -15812 8908
rect -15939 8828 -15892 8892
rect -15828 8828 -15812 8892
rect -15939 8812 -15812 8828
rect -15939 8748 -15892 8812
rect -15828 8748 -15812 8812
rect -15939 8732 -15812 8748
rect -15939 8668 -15892 8732
rect -15828 8668 -15812 8732
rect -15939 8652 -15812 8668
rect -15939 8588 -15892 8652
rect -15828 8588 -15812 8652
rect -15939 8572 -15812 8588
rect -15939 8508 -15892 8572
rect -15828 8508 -15812 8572
rect -15939 8492 -15812 8508
rect -15939 8428 -15892 8492
rect -15828 8428 -15812 8492
rect -15939 8412 -15812 8428
rect -15939 8348 -15892 8412
rect -15828 8348 -15812 8412
rect -15939 8332 -15812 8348
rect -15939 8268 -15892 8332
rect -15828 8268 -15812 8332
rect -15939 8252 -15812 8268
rect -15939 8188 -15892 8252
rect -15828 8188 -15812 8252
rect -15939 8172 -15812 8188
rect -15939 8108 -15892 8172
rect -15828 8108 -15812 8172
rect -15939 8092 -15812 8108
rect -15939 8028 -15892 8092
rect -15828 8028 -15812 8092
rect -15939 8012 -15812 8028
rect -15939 7948 -15892 8012
rect -15828 7948 -15812 8012
rect -15939 7932 -15812 7948
rect -15939 7868 -15892 7932
rect -15828 7868 -15812 7932
rect -15939 7852 -15812 7868
rect -15939 7788 -15892 7852
rect -15828 7788 -15812 7852
rect -15939 7772 -15812 7788
rect -15939 7708 -15892 7772
rect -15828 7708 -15812 7772
rect -15939 7692 -15812 7708
rect -15939 7628 -15892 7692
rect -15828 7628 -15812 7692
rect -15939 7612 -15812 7628
rect -15939 7548 -15892 7612
rect -15828 7548 -15812 7612
rect -15939 7532 -15812 7548
rect -15939 7468 -15892 7532
rect -15828 7468 -15812 7532
rect -15939 7452 -15812 7468
rect -15939 7388 -15892 7452
rect -15828 7388 -15812 7452
rect -15939 7372 -15812 7388
rect -15939 7308 -15892 7372
rect -15828 7308 -15812 7372
rect -15939 7292 -15812 7308
rect -15939 7228 -15892 7292
rect -15828 7228 -15812 7292
rect -15939 7212 -15812 7228
rect -15939 7148 -15892 7212
rect -15828 7148 -15812 7212
rect -15939 7132 -15812 7148
rect -15939 7068 -15892 7132
rect -15828 7068 -15812 7132
rect -15939 7052 -15812 7068
rect -15939 6988 -15892 7052
rect -15828 6988 -15812 7052
rect -15939 6972 -15812 6988
rect -15939 6908 -15892 6972
rect -15828 6908 -15812 6972
rect -15939 6892 -15812 6908
rect -15939 6828 -15892 6892
rect -15828 6828 -15812 6892
rect -15939 6812 -15812 6828
rect -15939 6748 -15892 6812
rect -15828 6748 -15812 6812
rect -15939 6732 -15812 6748
rect -15939 6668 -15892 6732
rect -15828 6668 -15812 6732
rect -15939 6652 -15812 6668
rect -15939 6588 -15892 6652
rect -15828 6588 -15812 6652
rect -15939 6572 -15812 6588
rect -15939 6508 -15892 6572
rect -15828 6508 -15812 6572
rect -15939 6492 -15812 6508
rect -15939 6428 -15892 6492
rect -15828 6428 -15812 6492
rect -15939 6412 -15812 6428
rect -15939 6348 -15892 6412
rect -15828 6348 -15812 6412
rect -15939 6332 -15812 6348
rect -15939 6268 -15892 6332
rect -15828 6268 -15812 6332
rect -15939 6252 -15812 6268
rect -15939 6188 -15892 6252
rect -15828 6188 -15812 6252
rect -15939 6172 -15812 6188
rect -15939 6108 -15892 6172
rect -15828 6108 -15812 6172
rect -15939 6092 -15812 6108
rect -15939 6028 -15892 6092
rect -15828 6028 -15812 6092
rect -15939 6012 -15812 6028
rect -15939 5948 -15892 6012
rect -15828 5948 -15812 6012
rect -15939 5932 -15812 5948
rect -15939 5868 -15892 5932
rect -15828 5868 -15812 5932
rect -15939 5852 -15812 5868
rect -15939 5788 -15892 5852
rect -15828 5788 -15812 5852
rect -15939 5772 -15812 5788
rect -15939 5708 -15892 5772
rect -15828 5708 -15812 5772
rect -15939 5692 -15812 5708
rect -15939 5628 -15892 5692
rect -15828 5628 -15812 5692
rect -15939 5612 -15812 5628
rect -15939 5548 -15892 5612
rect -15828 5548 -15812 5612
rect -15939 5532 -15812 5548
rect -15939 5468 -15892 5532
rect -15828 5468 -15812 5532
rect -15939 5452 -15812 5468
rect -15939 5388 -15892 5452
rect -15828 5388 -15812 5452
rect -15939 5372 -15812 5388
rect -15939 5308 -15892 5372
rect -15828 5308 -15812 5372
rect -15939 5292 -15812 5308
rect -15939 5228 -15892 5292
rect -15828 5228 -15812 5292
rect -15939 5212 -15812 5228
rect -15939 5148 -15892 5212
rect -15828 5148 -15812 5212
rect -15939 5132 -15812 5148
rect -15939 5068 -15892 5132
rect -15828 5068 -15812 5132
rect -15939 5052 -15812 5068
rect -15939 4988 -15892 5052
rect -15828 4988 -15812 5052
rect -15939 4972 -15812 4988
rect -15939 4908 -15892 4972
rect -15828 4908 -15812 4972
rect -15939 4892 -15812 4908
rect -15939 4828 -15892 4892
rect -15828 4828 -15812 4892
rect -15939 4812 -15812 4828
rect -15939 4748 -15892 4812
rect -15828 4748 -15812 4812
rect -15939 4732 -15812 4748
rect -15939 4668 -15892 4732
rect -15828 4668 -15812 4732
rect -15939 4652 -15812 4668
rect -15939 4588 -15892 4652
rect -15828 4588 -15812 4652
rect -15939 4572 -15812 4588
rect -15939 4508 -15892 4572
rect -15828 4508 -15812 4572
rect -15939 4492 -15812 4508
rect -15939 4428 -15892 4492
rect -15828 4428 -15812 4492
rect -15939 4412 -15812 4428
rect -15939 4348 -15892 4412
rect -15828 4348 -15812 4412
rect -15939 4332 -15812 4348
rect -15939 4268 -15892 4332
rect -15828 4268 -15812 4332
rect -15939 4252 -15812 4268
rect -15939 4188 -15892 4252
rect -15828 4188 -15812 4252
rect -15939 4172 -15812 4188
rect -15939 4108 -15892 4172
rect -15828 4108 -15812 4172
rect -15939 4092 -15812 4108
rect -15939 4028 -15892 4092
rect -15828 4028 -15812 4092
rect -15939 4012 -15812 4028
rect -15939 3948 -15892 4012
rect -15828 3948 -15812 4012
rect -15939 3932 -15812 3948
rect -15939 3868 -15892 3932
rect -15828 3868 -15812 3932
rect -15939 3852 -15812 3868
rect -15939 3788 -15892 3852
rect -15828 3788 -15812 3852
rect -15939 3772 -15812 3788
rect -15939 3708 -15892 3772
rect -15828 3708 -15812 3772
rect -15939 3692 -15812 3708
rect -15939 3628 -15892 3692
rect -15828 3628 -15812 3692
rect -15939 3612 -15812 3628
rect -15939 3548 -15892 3612
rect -15828 3548 -15812 3612
rect -15939 3532 -15812 3548
rect -15939 3468 -15892 3532
rect -15828 3468 -15812 3532
rect -15939 3452 -15812 3468
rect -15939 3388 -15892 3452
rect -15828 3388 -15812 3452
rect -15939 3372 -15812 3388
rect -22258 3292 -22131 3308
rect -22258 3228 -22211 3292
rect -22147 3228 -22131 3292
rect -22258 3212 -22131 3228
rect -22258 3088 -22154 3212
rect -22258 3072 -22131 3088
rect -22258 3008 -22211 3072
rect -22147 3008 -22131 3072
rect -22258 2992 -22131 3008
rect -28577 2912 -28450 2928
rect -28577 2848 -28530 2912
rect -28466 2848 -28450 2912
rect -28577 2832 -28450 2848
rect -28577 2768 -28530 2832
rect -28466 2768 -28450 2832
rect -28577 2752 -28450 2768
rect -28577 2688 -28530 2752
rect -28466 2688 -28450 2752
rect -28577 2672 -28450 2688
rect -28577 2608 -28530 2672
rect -28466 2608 -28450 2672
rect -28577 2592 -28450 2608
rect -28577 2528 -28530 2592
rect -28466 2528 -28450 2592
rect -28577 2512 -28450 2528
rect -28577 2448 -28530 2512
rect -28466 2448 -28450 2512
rect -28577 2432 -28450 2448
rect -28577 2368 -28530 2432
rect -28466 2368 -28450 2432
rect -28577 2352 -28450 2368
rect -28577 2288 -28530 2352
rect -28466 2288 -28450 2352
rect -28577 2272 -28450 2288
rect -28577 2208 -28530 2272
rect -28466 2208 -28450 2272
rect -28577 2192 -28450 2208
rect -28577 2128 -28530 2192
rect -28466 2128 -28450 2192
rect -28577 2112 -28450 2128
rect -28577 2048 -28530 2112
rect -28466 2048 -28450 2112
rect -28577 2032 -28450 2048
rect -28577 1968 -28530 2032
rect -28466 1968 -28450 2032
rect -28577 1952 -28450 1968
rect -28577 1888 -28530 1952
rect -28466 1888 -28450 1952
rect -28577 1872 -28450 1888
rect -28577 1808 -28530 1872
rect -28466 1808 -28450 1872
rect -28577 1792 -28450 1808
rect -28577 1728 -28530 1792
rect -28466 1728 -28450 1792
rect -28577 1712 -28450 1728
rect -28577 1648 -28530 1712
rect -28466 1648 -28450 1712
rect -28577 1632 -28450 1648
rect -28577 1568 -28530 1632
rect -28466 1568 -28450 1632
rect -28577 1552 -28450 1568
rect -28577 1488 -28530 1552
rect -28466 1488 -28450 1552
rect -28577 1472 -28450 1488
rect -28577 1408 -28530 1472
rect -28466 1408 -28450 1472
rect -28577 1392 -28450 1408
rect -28577 1328 -28530 1392
rect -28466 1328 -28450 1392
rect -28577 1312 -28450 1328
rect -28577 1248 -28530 1312
rect -28466 1248 -28450 1312
rect -28577 1232 -28450 1248
rect -28577 1168 -28530 1232
rect -28466 1168 -28450 1232
rect -28577 1152 -28450 1168
rect -28577 1088 -28530 1152
rect -28466 1088 -28450 1152
rect -28577 1072 -28450 1088
rect -28577 1008 -28530 1072
rect -28466 1008 -28450 1072
rect -28577 992 -28450 1008
rect -28577 928 -28530 992
rect -28466 928 -28450 992
rect -28577 912 -28450 928
rect -28577 848 -28530 912
rect -28466 848 -28450 912
rect -28577 832 -28450 848
rect -28577 768 -28530 832
rect -28466 768 -28450 832
rect -28577 752 -28450 768
rect -28577 688 -28530 752
rect -28466 688 -28450 752
rect -28577 672 -28450 688
rect -28577 608 -28530 672
rect -28466 608 -28450 672
rect -28577 592 -28450 608
rect -28577 528 -28530 592
rect -28466 528 -28450 592
rect -28577 512 -28450 528
rect -28577 448 -28530 512
rect -28466 448 -28450 512
rect -28577 432 -28450 448
rect -28577 368 -28530 432
rect -28466 368 -28450 432
rect -28577 352 -28450 368
rect -28577 288 -28530 352
rect -28466 288 -28450 352
rect -28577 272 -28450 288
rect -28577 208 -28530 272
rect -28466 208 -28450 272
rect -28577 192 -28450 208
rect -28577 128 -28530 192
rect -28466 128 -28450 192
rect -28577 112 -28450 128
rect -28577 48 -28530 112
rect -28466 48 -28450 112
rect -28577 32 -28450 48
rect -28577 -32 -28530 32
rect -28466 -32 -28450 32
rect -28577 -48 -28450 -32
rect -28577 -112 -28530 -48
rect -28466 -112 -28450 -48
rect -28577 -128 -28450 -112
rect -28577 -192 -28530 -128
rect -28466 -192 -28450 -128
rect -28577 -208 -28450 -192
rect -28577 -272 -28530 -208
rect -28466 -272 -28450 -208
rect -28577 -288 -28450 -272
rect -28577 -352 -28530 -288
rect -28466 -352 -28450 -288
rect -28577 -368 -28450 -352
rect -28577 -432 -28530 -368
rect -28466 -432 -28450 -368
rect -28577 -448 -28450 -432
rect -28577 -512 -28530 -448
rect -28466 -512 -28450 -448
rect -28577 -528 -28450 -512
rect -28577 -592 -28530 -528
rect -28466 -592 -28450 -528
rect -28577 -608 -28450 -592
rect -28577 -672 -28530 -608
rect -28466 -672 -28450 -608
rect -28577 -688 -28450 -672
rect -28577 -752 -28530 -688
rect -28466 -752 -28450 -688
rect -28577 -768 -28450 -752
rect -28577 -832 -28530 -768
rect -28466 -832 -28450 -768
rect -28577 -848 -28450 -832
rect -28577 -912 -28530 -848
rect -28466 -912 -28450 -848
rect -28577 -928 -28450 -912
rect -28577 -992 -28530 -928
rect -28466 -992 -28450 -928
rect -28577 -1008 -28450 -992
rect -28577 -1072 -28530 -1008
rect -28466 -1072 -28450 -1008
rect -28577 -1088 -28450 -1072
rect -28577 -1152 -28530 -1088
rect -28466 -1152 -28450 -1088
rect -28577 -1168 -28450 -1152
rect -28577 -1232 -28530 -1168
rect -28466 -1232 -28450 -1168
rect -28577 -1248 -28450 -1232
rect -28577 -1312 -28530 -1248
rect -28466 -1312 -28450 -1248
rect -28577 -1328 -28450 -1312
rect -28577 -1392 -28530 -1328
rect -28466 -1392 -28450 -1328
rect -28577 -1408 -28450 -1392
rect -28577 -1472 -28530 -1408
rect -28466 -1472 -28450 -1408
rect -28577 -1488 -28450 -1472
rect -28577 -1552 -28530 -1488
rect -28466 -1552 -28450 -1488
rect -28577 -1568 -28450 -1552
rect -28577 -1632 -28530 -1568
rect -28466 -1632 -28450 -1568
rect -28577 -1648 -28450 -1632
rect -28577 -1712 -28530 -1648
rect -28466 -1712 -28450 -1648
rect -28577 -1728 -28450 -1712
rect -28577 -1792 -28530 -1728
rect -28466 -1792 -28450 -1728
rect -28577 -1808 -28450 -1792
rect -28577 -1872 -28530 -1808
rect -28466 -1872 -28450 -1808
rect -28577 -1888 -28450 -1872
rect -28577 -1952 -28530 -1888
rect -28466 -1952 -28450 -1888
rect -28577 -1968 -28450 -1952
rect -28577 -2032 -28530 -1968
rect -28466 -2032 -28450 -1968
rect -28577 -2048 -28450 -2032
rect -28577 -2112 -28530 -2048
rect -28466 -2112 -28450 -2048
rect -28577 -2128 -28450 -2112
rect -28577 -2192 -28530 -2128
rect -28466 -2192 -28450 -2128
rect -28577 -2208 -28450 -2192
rect -28577 -2272 -28530 -2208
rect -28466 -2272 -28450 -2208
rect -28577 -2288 -28450 -2272
rect -28577 -2352 -28530 -2288
rect -28466 -2352 -28450 -2288
rect -28577 -2368 -28450 -2352
rect -28577 -2432 -28530 -2368
rect -28466 -2432 -28450 -2368
rect -28577 -2448 -28450 -2432
rect -28577 -2512 -28530 -2448
rect -28466 -2512 -28450 -2448
rect -28577 -2528 -28450 -2512
rect -28577 -2592 -28530 -2528
rect -28466 -2592 -28450 -2528
rect -28577 -2608 -28450 -2592
rect -28577 -2672 -28530 -2608
rect -28466 -2672 -28450 -2608
rect -28577 -2688 -28450 -2672
rect -28577 -2752 -28530 -2688
rect -28466 -2752 -28450 -2688
rect -28577 -2768 -28450 -2752
rect -28577 -2832 -28530 -2768
rect -28466 -2832 -28450 -2768
rect -28577 -2848 -28450 -2832
rect -28577 -2912 -28530 -2848
rect -28466 -2912 -28450 -2848
rect -28577 -2928 -28450 -2912
rect -34896 -3008 -34769 -2992
rect -34896 -3072 -34849 -3008
rect -34785 -3072 -34769 -3008
rect -34896 -3088 -34769 -3072
rect -34896 -3212 -34792 -3088
rect -34896 -3228 -34769 -3212
rect -34896 -3292 -34849 -3228
rect -34785 -3292 -34769 -3228
rect -34896 -3308 -34769 -3292
rect -41215 -3388 -41088 -3372
rect -41215 -3452 -41168 -3388
rect -41104 -3452 -41088 -3388
rect -41215 -3468 -41088 -3452
rect -41215 -3532 -41168 -3468
rect -41104 -3532 -41088 -3468
rect -41215 -3548 -41088 -3532
rect -41215 -3612 -41168 -3548
rect -41104 -3612 -41088 -3548
rect -41215 -3628 -41088 -3612
rect -41215 -3692 -41168 -3628
rect -41104 -3692 -41088 -3628
rect -41215 -3708 -41088 -3692
rect -41215 -3772 -41168 -3708
rect -41104 -3772 -41088 -3708
rect -41215 -3788 -41088 -3772
rect -41215 -3852 -41168 -3788
rect -41104 -3852 -41088 -3788
rect -41215 -3868 -41088 -3852
rect -41215 -3932 -41168 -3868
rect -41104 -3932 -41088 -3868
rect -41215 -3948 -41088 -3932
rect -41215 -4012 -41168 -3948
rect -41104 -4012 -41088 -3948
rect -41215 -4028 -41088 -4012
rect -41215 -4092 -41168 -4028
rect -41104 -4092 -41088 -4028
rect -41215 -4108 -41088 -4092
rect -41215 -4172 -41168 -4108
rect -41104 -4172 -41088 -4108
rect -41215 -4188 -41088 -4172
rect -41215 -4252 -41168 -4188
rect -41104 -4252 -41088 -4188
rect -41215 -4268 -41088 -4252
rect -41215 -4332 -41168 -4268
rect -41104 -4332 -41088 -4268
rect -41215 -4348 -41088 -4332
rect -41215 -4412 -41168 -4348
rect -41104 -4412 -41088 -4348
rect -41215 -4428 -41088 -4412
rect -41215 -4492 -41168 -4428
rect -41104 -4492 -41088 -4428
rect -41215 -4508 -41088 -4492
rect -41215 -4572 -41168 -4508
rect -41104 -4572 -41088 -4508
rect -41215 -4588 -41088 -4572
rect -41215 -4652 -41168 -4588
rect -41104 -4652 -41088 -4588
rect -41215 -4668 -41088 -4652
rect -41215 -4732 -41168 -4668
rect -41104 -4732 -41088 -4668
rect -41215 -4748 -41088 -4732
rect -41215 -4812 -41168 -4748
rect -41104 -4812 -41088 -4748
rect -41215 -4828 -41088 -4812
rect -41215 -4892 -41168 -4828
rect -41104 -4892 -41088 -4828
rect -41215 -4908 -41088 -4892
rect -41215 -4972 -41168 -4908
rect -41104 -4972 -41088 -4908
rect -41215 -4988 -41088 -4972
rect -41215 -5052 -41168 -4988
rect -41104 -5052 -41088 -4988
rect -41215 -5068 -41088 -5052
rect -41215 -5132 -41168 -5068
rect -41104 -5132 -41088 -5068
rect -41215 -5148 -41088 -5132
rect -41215 -5212 -41168 -5148
rect -41104 -5212 -41088 -5148
rect -41215 -5228 -41088 -5212
rect -41215 -5292 -41168 -5228
rect -41104 -5292 -41088 -5228
rect -41215 -5308 -41088 -5292
rect -41215 -5372 -41168 -5308
rect -41104 -5372 -41088 -5308
rect -41215 -5388 -41088 -5372
rect -41215 -5452 -41168 -5388
rect -41104 -5452 -41088 -5388
rect -41215 -5468 -41088 -5452
rect -41215 -5532 -41168 -5468
rect -41104 -5532 -41088 -5468
rect -41215 -5548 -41088 -5532
rect -41215 -5612 -41168 -5548
rect -41104 -5612 -41088 -5548
rect -41215 -5628 -41088 -5612
rect -41215 -5692 -41168 -5628
rect -41104 -5692 -41088 -5628
rect -41215 -5708 -41088 -5692
rect -41215 -5772 -41168 -5708
rect -41104 -5772 -41088 -5708
rect -41215 -5788 -41088 -5772
rect -41215 -5852 -41168 -5788
rect -41104 -5852 -41088 -5788
rect -41215 -5868 -41088 -5852
rect -41215 -5932 -41168 -5868
rect -41104 -5932 -41088 -5868
rect -41215 -5948 -41088 -5932
rect -41215 -6012 -41168 -5948
rect -41104 -6012 -41088 -5948
rect -41215 -6028 -41088 -6012
rect -41215 -6092 -41168 -6028
rect -41104 -6092 -41088 -6028
rect -41215 -6108 -41088 -6092
rect -41215 -6172 -41168 -6108
rect -41104 -6172 -41088 -6108
rect -41215 -6188 -41088 -6172
rect -41215 -6252 -41168 -6188
rect -41104 -6252 -41088 -6188
rect -41215 -6268 -41088 -6252
rect -41215 -6332 -41168 -6268
rect -41104 -6332 -41088 -6268
rect -41215 -6348 -41088 -6332
rect -41215 -6412 -41168 -6348
rect -41104 -6412 -41088 -6348
rect -41215 -6428 -41088 -6412
rect -41215 -6492 -41168 -6428
rect -41104 -6492 -41088 -6428
rect -41215 -6508 -41088 -6492
rect -41215 -6572 -41168 -6508
rect -41104 -6572 -41088 -6508
rect -41215 -6588 -41088 -6572
rect -41215 -6652 -41168 -6588
rect -41104 -6652 -41088 -6588
rect -41215 -6668 -41088 -6652
rect -41215 -6732 -41168 -6668
rect -41104 -6732 -41088 -6668
rect -41215 -6748 -41088 -6732
rect -41215 -6812 -41168 -6748
rect -41104 -6812 -41088 -6748
rect -41215 -6828 -41088 -6812
rect -41215 -6892 -41168 -6828
rect -41104 -6892 -41088 -6828
rect -41215 -6908 -41088 -6892
rect -41215 -6972 -41168 -6908
rect -41104 -6972 -41088 -6908
rect -41215 -6988 -41088 -6972
rect -41215 -7052 -41168 -6988
rect -41104 -7052 -41088 -6988
rect -41215 -7068 -41088 -7052
rect -41215 -7132 -41168 -7068
rect -41104 -7132 -41088 -7068
rect -41215 -7148 -41088 -7132
rect -41215 -7212 -41168 -7148
rect -41104 -7212 -41088 -7148
rect -41215 -7228 -41088 -7212
rect -41215 -7292 -41168 -7228
rect -41104 -7292 -41088 -7228
rect -41215 -7308 -41088 -7292
rect -41215 -7372 -41168 -7308
rect -41104 -7372 -41088 -7308
rect -41215 -7388 -41088 -7372
rect -41215 -7452 -41168 -7388
rect -41104 -7452 -41088 -7388
rect -41215 -7468 -41088 -7452
rect -41215 -7532 -41168 -7468
rect -41104 -7532 -41088 -7468
rect -41215 -7548 -41088 -7532
rect -41215 -7612 -41168 -7548
rect -41104 -7612 -41088 -7548
rect -41215 -7628 -41088 -7612
rect -41215 -7692 -41168 -7628
rect -41104 -7692 -41088 -7628
rect -41215 -7708 -41088 -7692
rect -41215 -7772 -41168 -7708
rect -41104 -7772 -41088 -7708
rect -41215 -7788 -41088 -7772
rect -41215 -7852 -41168 -7788
rect -41104 -7852 -41088 -7788
rect -41215 -7868 -41088 -7852
rect -41215 -7932 -41168 -7868
rect -41104 -7932 -41088 -7868
rect -41215 -7948 -41088 -7932
rect -41215 -8012 -41168 -7948
rect -41104 -8012 -41088 -7948
rect -41215 -8028 -41088 -8012
rect -41215 -8092 -41168 -8028
rect -41104 -8092 -41088 -8028
rect -41215 -8108 -41088 -8092
rect -41215 -8172 -41168 -8108
rect -41104 -8172 -41088 -8108
rect -41215 -8188 -41088 -8172
rect -41215 -8252 -41168 -8188
rect -41104 -8252 -41088 -8188
rect -41215 -8268 -41088 -8252
rect -41215 -8332 -41168 -8268
rect -41104 -8332 -41088 -8268
rect -41215 -8348 -41088 -8332
rect -41215 -8412 -41168 -8348
rect -41104 -8412 -41088 -8348
rect -41215 -8428 -41088 -8412
rect -41215 -8492 -41168 -8428
rect -41104 -8492 -41088 -8428
rect -41215 -8508 -41088 -8492
rect -41215 -8572 -41168 -8508
rect -41104 -8572 -41088 -8508
rect -41215 -8588 -41088 -8572
rect -41215 -8652 -41168 -8588
rect -41104 -8652 -41088 -8588
rect -41215 -8668 -41088 -8652
rect -41215 -8732 -41168 -8668
rect -41104 -8732 -41088 -8668
rect -41215 -8748 -41088 -8732
rect -41215 -8812 -41168 -8748
rect -41104 -8812 -41088 -8748
rect -41215 -8828 -41088 -8812
rect -41215 -8892 -41168 -8828
rect -41104 -8892 -41088 -8828
rect -41215 -8908 -41088 -8892
rect -41215 -8972 -41168 -8908
rect -41104 -8972 -41088 -8908
rect -41215 -8988 -41088 -8972
rect -41215 -9052 -41168 -8988
rect -41104 -9052 -41088 -8988
rect -41215 -9068 -41088 -9052
rect -41215 -9132 -41168 -9068
rect -41104 -9132 -41088 -9068
rect -41215 -9148 -41088 -9132
rect -41215 -9212 -41168 -9148
rect -41104 -9212 -41088 -9148
rect -41215 -9228 -41088 -9212
rect -44335 -9639 -44231 -9261
rect -41215 -9292 -41168 -9228
rect -41104 -9292 -41088 -9228
rect -40925 -3348 -35003 -3339
rect -40925 -9252 -40916 -3348
rect -35012 -9252 -35003 -3348
rect -40925 -9261 -35003 -9252
rect -34896 -3372 -34849 -3308
rect -34785 -3372 -34769 -3308
rect -31697 -3339 -31593 -2961
rect -28577 -2992 -28530 -2928
rect -28466 -2992 -28450 -2928
rect -28287 2952 -22365 2961
rect -28287 -2952 -28278 2952
rect -22374 -2952 -22365 2952
rect -28287 -2961 -22365 -2952
rect -22258 2928 -22211 2992
rect -22147 2928 -22131 2992
rect -19059 2961 -18955 3339
rect -15939 3308 -15892 3372
rect -15828 3308 -15812 3372
rect -15649 9252 -9727 9261
rect -15649 3348 -15640 9252
rect -9736 3348 -9727 9252
rect -15649 3339 -9727 3348
rect -9620 9228 -9573 9292
rect -9509 9228 -9493 9292
rect -6421 9261 -6317 9639
rect -3301 9608 -3254 9672
rect -3190 9608 -3174 9672
rect -3011 15552 2911 15561
rect -3011 9648 -3002 15552
rect 2902 9648 2911 15552
rect -3011 9639 2911 9648
rect 3018 15528 3065 15592
rect 3129 15528 3145 15592
rect 6217 15561 6321 15939
rect 9337 15908 9384 15972
rect 9448 15908 9464 15972
rect 9627 21852 15549 21861
rect 9627 15948 9636 21852
rect 15540 15948 15549 21852
rect 9627 15939 15549 15948
rect 15656 21828 15703 21892
rect 15767 21828 15783 21892
rect 18855 21861 18959 22239
rect 21975 22208 22022 22272
rect 22086 22208 22102 22272
rect 22265 28152 28187 28161
rect 22265 22248 22274 28152
rect 28178 22248 28187 28152
rect 22265 22239 28187 22248
rect 28294 28128 28341 28192
rect 28405 28128 28421 28192
rect 31493 28161 31597 28539
rect 34613 28508 34660 28572
rect 34724 28508 34740 28572
rect 34903 34452 40825 34461
rect 34903 28548 34912 34452
rect 40816 28548 40825 34452
rect 34903 28539 40825 28548
rect 40932 34428 40979 34492
rect 41043 34428 41059 34492
rect 44131 34461 44235 34839
rect 47251 34808 47298 34872
rect 47362 34808 47378 34872
rect 47251 34792 47378 34808
rect 47251 34728 47298 34792
rect 47362 34728 47378 34792
rect 47251 34712 47378 34728
rect 47251 34588 47355 34712
rect 47251 34572 47378 34588
rect 47251 34508 47298 34572
rect 47362 34508 47378 34572
rect 47251 34492 47378 34508
rect 40932 34412 41059 34428
rect 40932 34348 40979 34412
rect 41043 34348 41059 34412
rect 40932 34332 41059 34348
rect 40932 34268 40979 34332
rect 41043 34268 41059 34332
rect 40932 34252 41059 34268
rect 40932 34188 40979 34252
rect 41043 34188 41059 34252
rect 40932 34172 41059 34188
rect 40932 34108 40979 34172
rect 41043 34108 41059 34172
rect 40932 34092 41059 34108
rect 40932 34028 40979 34092
rect 41043 34028 41059 34092
rect 40932 34012 41059 34028
rect 40932 33948 40979 34012
rect 41043 33948 41059 34012
rect 40932 33932 41059 33948
rect 40932 33868 40979 33932
rect 41043 33868 41059 33932
rect 40932 33852 41059 33868
rect 40932 33788 40979 33852
rect 41043 33788 41059 33852
rect 40932 33772 41059 33788
rect 40932 33708 40979 33772
rect 41043 33708 41059 33772
rect 40932 33692 41059 33708
rect 40932 33628 40979 33692
rect 41043 33628 41059 33692
rect 40932 33612 41059 33628
rect 40932 33548 40979 33612
rect 41043 33548 41059 33612
rect 40932 33532 41059 33548
rect 40932 33468 40979 33532
rect 41043 33468 41059 33532
rect 40932 33452 41059 33468
rect 40932 33388 40979 33452
rect 41043 33388 41059 33452
rect 40932 33372 41059 33388
rect 40932 33308 40979 33372
rect 41043 33308 41059 33372
rect 40932 33292 41059 33308
rect 40932 33228 40979 33292
rect 41043 33228 41059 33292
rect 40932 33212 41059 33228
rect 40932 33148 40979 33212
rect 41043 33148 41059 33212
rect 40932 33132 41059 33148
rect 40932 33068 40979 33132
rect 41043 33068 41059 33132
rect 40932 33052 41059 33068
rect 40932 32988 40979 33052
rect 41043 32988 41059 33052
rect 40932 32972 41059 32988
rect 40932 32908 40979 32972
rect 41043 32908 41059 32972
rect 40932 32892 41059 32908
rect 40932 32828 40979 32892
rect 41043 32828 41059 32892
rect 40932 32812 41059 32828
rect 40932 32748 40979 32812
rect 41043 32748 41059 32812
rect 40932 32732 41059 32748
rect 40932 32668 40979 32732
rect 41043 32668 41059 32732
rect 40932 32652 41059 32668
rect 40932 32588 40979 32652
rect 41043 32588 41059 32652
rect 40932 32572 41059 32588
rect 40932 32508 40979 32572
rect 41043 32508 41059 32572
rect 40932 32492 41059 32508
rect 40932 32428 40979 32492
rect 41043 32428 41059 32492
rect 40932 32412 41059 32428
rect 40932 32348 40979 32412
rect 41043 32348 41059 32412
rect 40932 32332 41059 32348
rect 40932 32268 40979 32332
rect 41043 32268 41059 32332
rect 40932 32252 41059 32268
rect 40932 32188 40979 32252
rect 41043 32188 41059 32252
rect 40932 32172 41059 32188
rect 40932 32108 40979 32172
rect 41043 32108 41059 32172
rect 40932 32092 41059 32108
rect 40932 32028 40979 32092
rect 41043 32028 41059 32092
rect 40932 32012 41059 32028
rect 40932 31948 40979 32012
rect 41043 31948 41059 32012
rect 40932 31932 41059 31948
rect 40932 31868 40979 31932
rect 41043 31868 41059 31932
rect 40932 31852 41059 31868
rect 40932 31788 40979 31852
rect 41043 31788 41059 31852
rect 40932 31772 41059 31788
rect 40932 31708 40979 31772
rect 41043 31708 41059 31772
rect 40932 31692 41059 31708
rect 40932 31628 40979 31692
rect 41043 31628 41059 31692
rect 40932 31612 41059 31628
rect 40932 31548 40979 31612
rect 41043 31548 41059 31612
rect 40932 31532 41059 31548
rect 40932 31468 40979 31532
rect 41043 31468 41059 31532
rect 40932 31452 41059 31468
rect 40932 31388 40979 31452
rect 41043 31388 41059 31452
rect 40932 31372 41059 31388
rect 40932 31308 40979 31372
rect 41043 31308 41059 31372
rect 40932 31292 41059 31308
rect 40932 31228 40979 31292
rect 41043 31228 41059 31292
rect 40932 31212 41059 31228
rect 40932 31148 40979 31212
rect 41043 31148 41059 31212
rect 40932 31132 41059 31148
rect 40932 31068 40979 31132
rect 41043 31068 41059 31132
rect 40932 31052 41059 31068
rect 40932 30988 40979 31052
rect 41043 30988 41059 31052
rect 40932 30972 41059 30988
rect 40932 30908 40979 30972
rect 41043 30908 41059 30972
rect 40932 30892 41059 30908
rect 40932 30828 40979 30892
rect 41043 30828 41059 30892
rect 40932 30812 41059 30828
rect 40932 30748 40979 30812
rect 41043 30748 41059 30812
rect 40932 30732 41059 30748
rect 40932 30668 40979 30732
rect 41043 30668 41059 30732
rect 40932 30652 41059 30668
rect 40932 30588 40979 30652
rect 41043 30588 41059 30652
rect 40932 30572 41059 30588
rect 40932 30508 40979 30572
rect 41043 30508 41059 30572
rect 40932 30492 41059 30508
rect 40932 30428 40979 30492
rect 41043 30428 41059 30492
rect 40932 30412 41059 30428
rect 40932 30348 40979 30412
rect 41043 30348 41059 30412
rect 40932 30332 41059 30348
rect 40932 30268 40979 30332
rect 41043 30268 41059 30332
rect 40932 30252 41059 30268
rect 40932 30188 40979 30252
rect 41043 30188 41059 30252
rect 40932 30172 41059 30188
rect 40932 30108 40979 30172
rect 41043 30108 41059 30172
rect 40932 30092 41059 30108
rect 40932 30028 40979 30092
rect 41043 30028 41059 30092
rect 40932 30012 41059 30028
rect 40932 29948 40979 30012
rect 41043 29948 41059 30012
rect 40932 29932 41059 29948
rect 40932 29868 40979 29932
rect 41043 29868 41059 29932
rect 40932 29852 41059 29868
rect 40932 29788 40979 29852
rect 41043 29788 41059 29852
rect 40932 29772 41059 29788
rect 40932 29708 40979 29772
rect 41043 29708 41059 29772
rect 40932 29692 41059 29708
rect 40932 29628 40979 29692
rect 41043 29628 41059 29692
rect 40932 29612 41059 29628
rect 40932 29548 40979 29612
rect 41043 29548 41059 29612
rect 40932 29532 41059 29548
rect 40932 29468 40979 29532
rect 41043 29468 41059 29532
rect 40932 29452 41059 29468
rect 40932 29388 40979 29452
rect 41043 29388 41059 29452
rect 40932 29372 41059 29388
rect 40932 29308 40979 29372
rect 41043 29308 41059 29372
rect 40932 29292 41059 29308
rect 40932 29228 40979 29292
rect 41043 29228 41059 29292
rect 40932 29212 41059 29228
rect 40932 29148 40979 29212
rect 41043 29148 41059 29212
rect 40932 29132 41059 29148
rect 40932 29068 40979 29132
rect 41043 29068 41059 29132
rect 40932 29052 41059 29068
rect 40932 28988 40979 29052
rect 41043 28988 41059 29052
rect 40932 28972 41059 28988
rect 40932 28908 40979 28972
rect 41043 28908 41059 28972
rect 40932 28892 41059 28908
rect 40932 28828 40979 28892
rect 41043 28828 41059 28892
rect 40932 28812 41059 28828
rect 40932 28748 40979 28812
rect 41043 28748 41059 28812
rect 40932 28732 41059 28748
rect 40932 28668 40979 28732
rect 41043 28668 41059 28732
rect 40932 28652 41059 28668
rect 40932 28588 40979 28652
rect 41043 28588 41059 28652
rect 40932 28572 41059 28588
rect 34613 28492 34740 28508
rect 34613 28428 34660 28492
rect 34724 28428 34740 28492
rect 34613 28412 34740 28428
rect 34613 28288 34717 28412
rect 34613 28272 34740 28288
rect 34613 28208 34660 28272
rect 34724 28208 34740 28272
rect 34613 28192 34740 28208
rect 28294 28112 28421 28128
rect 28294 28048 28341 28112
rect 28405 28048 28421 28112
rect 28294 28032 28421 28048
rect 28294 27968 28341 28032
rect 28405 27968 28421 28032
rect 28294 27952 28421 27968
rect 28294 27888 28341 27952
rect 28405 27888 28421 27952
rect 28294 27872 28421 27888
rect 28294 27808 28341 27872
rect 28405 27808 28421 27872
rect 28294 27792 28421 27808
rect 28294 27728 28341 27792
rect 28405 27728 28421 27792
rect 28294 27712 28421 27728
rect 28294 27648 28341 27712
rect 28405 27648 28421 27712
rect 28294 27632 28421 27648
rect 28294 27568 28341 27632
rect 28405 27568 28421 27632
rect 28294 27552 28421 27568
rect 28294 27488 28341 27552
rect 28405 27488 28421 27552
rect 28294 27472 28421 27488
rect 28294 27408 28341 27472
rect 28405 27408 28421 27472
rect 28294 27392 28421 27408
rect 28294 27328 28341 27392
rect 28405 27328 28421 27392
rect 28294 27312 28421 27328
rect 28294 27248 28341 27312
rect 28405 27248 28421 27312
rect 28294 27232 28421 27248
rect 28294 27168 28341 27232
rect 28405 27168 28421 27232
rect 28294 27152 28421 27168
rect 28294 27088 28341 27152
rect 28405 27088 28421 27152
rect 28294 27072 28421 27088
rect 28294 27008 28341 27072
rect 28405 27008 28421 27072
rect 28294 26992 28421 27008
rect 28294 26928 28341 26992
rect 28405 26928 28421 26992
rect 28294 26912 28421 26928
rect 28294 26848 28341 26912
rect 28405 26848 28421 26912
rect 28294 26832 28421 26848
rect 28294 26768 28341 26832
rect 28405 26768 28421 26832
rect 28294 26752 28421 26768
rect 28294 26688 28341 26752
rect 28405 26688 28421 26752
rect 28294 26672 28421 26688
rect 28294 26608 28341 26672
rect 28405 26608 28421 26672
rect 28294 26592 28421 26608
rect 28294 26528 28341 26592
rect 28405 26528 28421 26592
rect 28294 26512 28421 26528
rect 28294 26448 28341 26512
rect 28405 26448 28421 26512
rect 28294 26432 28421 26448
rect 28294 26368 28341 26432
rect 28405 26368 28421 26432
rect 28294 26352 28421 26368
rect 28294 26288 28341 26352
rect 28405 26288 28421 26352
rect 28294 26272 28421 26288
rect 28294 26208 28341 26272
rect 28405 26208 28421 26272
rect 28294 26192 28421 26208
rect 28294 26128 28341 26192
rect 28405 26128 28421 26192
rect 28294 26112 28421 26128
rect 28294 26048 28341 26112
rect 28405 26048 28421 26112
rect 28294 26032 28421 26048
rect 28294 25968 28341 26032
rect 28405 25968 28421 26032
rect 28294 25952 28421 25968
rect 28294 25888 28341 25952
rect 28405 25888 28421 25952
rect 28294 25872 28421 25888
rect 28294 25808 28341 25872
rect 28405 25808 28421 25872
rect 28294 25792 28421 25808
rect 28294 25728 28341 25792
rect 28405 25728 28421 25792
rect 28294 25712 28421 25728
rect 28294 25648 28341 25712
rect 28405 25648 28421 25712
rect 28294 25632 28421 25648
rect 28294 25568 28341 25632
rect 28405 25568 28421 25632
rect 28294 25552 28421 25568
rect 28294 25488 28341 25552
rect 28405 25488 28421 25552
rect 28294 25472 28421 25488
rect 28294 25408 28341 25472
rect 28405 25408 28421 25472
rect 28294 25392 28421 25408
rect 28294 25328 28341 25392
rect 28405 25328 28421 25392
rect 28294 25312 28421 25328
rect 28294 25248 28341 25312
rect 28405 25248 28421 25312
rect 28294 25232 28421 25248
rect 28294 25168 28341 25232
rect 28405 25168 28421 25232
rect 28294 25152 28421 25168
rect 28294 25088 28341 25152
rect 28405 25088 28421 25152
rect 28294 25072 28421 25088
rect 28294 25008 28341 25072
rect 28405 25008 28421 25072
rect 28294 24992 28421 25008
rect 28294 24928 28341 24992
rect 28405 24928 28421 24992
rect 28294 24912 28421 24928
rect 28294 24848 28341 24912
rect 28405 24848 28421 24912
rect 28294 24832 28421 24848
rect 28294 24768 28341 24832
rect 28405 24768 28421 24832
rect 28294 24752 28421 24768
rect 28294 24688 28341 24752
rect 28405 24688 28421 24752
rect 28294 24672 28421 24688
rect 28294 24608 28341 24672
rect 28405 24608 28421 24672
rect 28294 24592 28421 24608
rect 28294 24528 28341 24592
rect 28405 24528 28421 24592
rect 28294 24512 28421 24528
rect 28294 24448 28341 24512
rect 28405 24448 28421 24512
rect 28294 24432 28421 24448
rect 28294 24368 28341 24432
rect 28405 24368 28421 24432
rect 28294 24352 28421 24368
rect 28294 24288 28341 24352
rect 28405 24288 28421 24352
rect 28294 24272 28421 24288
rect 28294 24208 28341 24272
rect 28405 24208 28421 24272
rect 28294 24192 28421 24208
rect 28294 24128 28341 24192
rect 28405 24128 28421 24192
rect 28294 24112 28421 24128
rect 28294 24048 28341 24112
rect 28405 24048 28421 24112
rect 28294 24032 28421 24048
rect 28294 23968 28341 24032
rect 28405 23968 28421 24032
rect 28294 23952 28421 23968
rect 28294 23888 28341 23952
rect 28405 23888 28421 23952
rect 28294 23872 28421 23888
rect 28294 23808 28341 23872
rect 28405 23808 28421 23872
rect 28294 23792 28421 23808
rect 28294 23728 28341 23792
rect 28405 23728 28421 23792
rect 28294 23712 28421 23728
rect 28294 23648 28341 23712
rect 28405 23648 28421 23712
rect 28294 23632 28421 23648
rect 28294 23568 28341 23632
rect 28405 23568 28421 23632
rect 28294 23552 28421 23568
rect 28294 23488 28341 23552
rect 28405 23488 28421 23552
rect 28294 23472 28421 23488
rect 28294 23408 28341 23472
rect 28405 23408 28421 23472
rect 28294 23392 28421 23408
rect 28294 23328 28341 23392
rect 28405 23328 28421 23392
rect 28294 23312 28421 23328
rect 28294 23248 28341 23312
rect 28405 23248 28421 23312
rect 28294 23232 28421 23248
rect 28294 23168 28341 23232
rect 28405 23168 28421 23232
rect 28294 23152 28421 23168
rect 28294 23088 28341 23152
rect 28405 23088 28421 23152
rect 28294 23072 28421 23088
rect 28294 23008 28341 23072
rect 28405 23008 28421 23072
rect 28294 22992 28421 23008
rect 28294 22928 28341 22992
rect 28405 22928 28421 22992
rect 28294 22912 28421 22928
rect 28294 22848 28341 22912
rect 28405 22848 28421 22912
rect 28294 22832 28421 22848
rect 28294 22768 28341 22832
rect 28405 22768 28421 22832
rect 28294 22752 28421 22768
rect 28294 22688 28341 22752
rect 28405 22688 28421 22752
rect 28294 22672 28421 22688
rect 28294 22608 28341 22672
rect 28405 22608 28421 22672
rect 28294 22592 28421 22608
rect 28294 22528 28341 22592
rect 28405 22528 28421 22592
rect 28294 22512 28421 22528
rect 28294 22448 28341 22512
rect 28405 22448 28421 22512
rect 28294 22432 28421 22448
rect 28294 22368 28341 22432
rect 28405 22368 28421 22432
rect 28294 22352 28421 22368
rect 28294 22288 28341 22352
rect 28405 22288 28421 22352
rect 28294 22272 28421 22288
rect 21975 22192 22102 22208
rect 21975 22128 22022 22192
rect 22086 22128 22102 22192
rect 21975 22112 22102 22128
rect 21975 21988 22079 22112
rect 21975 21972 22102 21988
rect 21975 21908 22022 21972
rect 22086 21908 22102 21972
rect 21975 21892 22102 21908
rect 15656 21812 15783 21828
rect 15656 21748 15703 21812
rect 15767 21748 15783 21812
rect 15656 21732 15783 21748
rect 15656 21668 15703 21732
rect 15767 21668 15783 21732
rect 15656 21652 15783 21668
rect 15656 21588 15703 21652
rect 15767 21588 15783 21652
rect 15656 21572 15783 21588
rect 15656 21508 15703 21572
rect 15767 21508 15783 21572
rect 15656 21492 15783 21508
rect 15656 21428 15703 21492
rect 15767 21428 15783 21492
rect 15656 21412 15783 21428
rect 15656 21348 15703 21412
rect 15767 21348 15783 21412
rect 15656 21332 15783 21348
rect 15656 21268 15703 21332
rect 15767 21268 15783 21332
rect 15656 21252 15783 21268
rect 15656 21188 15703 21252
rect 15767 21188 15783 21252
rect 15656 21172 15783 21188
rect 15656 21108 15703 21172
rect 15767 21108 15783 21172
rect 15656 21092 15783 21108
rect 15656 21028 15703 21092
rect 15767 21028 15783 21092
rect 15656 21012 15783 21028
rect 15656 20948 15703 21012
rect 15767 20948 15783 21012
rect 15656 20932 15783 20948
rect 15656 20868 15703 20932
rect 15767 20868 15783 20932
rect 15656 20852 15783 20868
rect 15656 20788 15703 20852
rect 15767 20788 15783 20852
rect 15656 20772 15783 20788
rect 15656 20708 15703 20772
rect 15767 20708 15783 20772
rect 15656 20692 15783 20708
rect 15656 20628 15703 20692
rect 15767 20628 15783 20692
rect 15656 20612 15783 20628
rect 15656 20548 15703 20612
rect 15767 20548 15783 20612
rect 15656 20532 15783 20548
rect 15656 20468 15703 20532
rect 15767 20468 15783 20532
rect 15656 20452 15783 20468
rect 15656 20388 15703 20452
rect 15767 20388 15783 20452
rect 15656 20372 15783 20388
rect 15656 20308 15703 20372
rect 15767 20308 15783 20372
rect 15656 20292 15783 20308
rect 15656 20228 15703 20292
rect 15767 20228 15783 20292
rect 15656 20212 15783 20228
rect 15656 20148 15703 20212
rect 15767 20148 15783 20212
rect 15656 20132 15783 20148
rect 15656 20068 15703 20132
rect 15767 20068 15783 20132
rect 15656 20052 15783 20068
rect 15656 19988 15703 20052
rect 15767 19988 15783 20052
rect 15656 19972 15783 19988
rect 15656 19908 15703 19972
rect 15767 19908 15783 19972
rect 15656 19892 15783 19908
rect 15656 19828 15703 19892
rect 15767 19828 15783 19892
rect 15656 19812 15783 19828
rect 15656 19748 15703 19812
rect 15767 19748 15783 19812
rect 15656 19732 15783 19748
rect 15656 19668 15703 19732
rect 15767 19668 15783 19732
rect 15656 19652 15783 19668
rect 15656 19588 15703 19652
rect 15767 19588 15783 19652
rect 15656 19572 15783 19588
rect 15656 19508 15703 19572
rect 15767 19508 15783 19572
rect 15656 19492 15783 19508
rect 15656 19428 15703 19492
rect 15767 19428 15783 19492
rect 15656 19412 15783 19428
rect 15656 19348 15703 19412
rect 15767 19348 15783 19412
rect 15656 19332 15783 19348
rect 15656 19268 15703 19332
rect 15767 19268 15783 19332
rect 15656 19252 15783 19268
rect 15656 19188 15703 19252
rect 15767 19188 15783 19252
rect 15656 19172 15783 19188
rect 15656 19108 15703 19172
rect 15767 19108 15783 19172
rect 15656 19092 15783 19108
rect 15656 19028 15703 19092
rect 15767 19028 15783 19092
rect 15656 19012 15783 19028
rect 15656 18948 15703 19012
rect 15767 18948 15783 19012
rect 15656 18932 15783 18948
rect 15656 18868 15703 18932
rect 15767 18868 15783 18932
rect 15656 18852 15783 18868
rect 15656 18788 15703 18852
rect 15767 18788 15783 18852
rect 15656 18772 15783 18788
rect 15656 18708 15703 18772
rect 15767 18708 15783 18772
rect 15656 18692 15783 18708
rect 15656 18628 15703 18692
rect 15767 18628 15783 18692
rect 15656 18612 15783 18628
rect 15656 18548 15703 18612
rect 15767 18548 15783 18612
rect 15656 18532 15783 18548
rect 15656 18468 15703 18532
rect 15767 18468 15783 18532
rect 15656 18452 15783 18468
rect 15656 18388 15703 18452
rect 15767 18388 15783 18452
rect 15656 18372 15783 18388
rect 15656 18308 15703 18372
rect 15767 18308 15783 18372
rect 15656 18292 15783 18308
rect 15656 18228 15703 18292
rect 15767 18228 15783 18292
rect 15656 18212 15783 18228
rect 15656 18148 15703 18212
rect 15767 18148 15783 18212
rect 15656 18132 15783 18148
rect 15656 18068 15703 18132
rect 15767 18068 15783 18132
rect 15656 18052 15783 18068
rect 15656 17988 15703 18052
rect 15767 17988 15783 18052
rect 15656 17972 15783 17988
rect 15656 17908 15703 17972
rect 15767 17908 15783 17972
rect 15656 17892 15783 17908
rect 15656 17828 15703 17892
rect 15767 17828 15783 17892
rect 15656 17812 15783 17828
rect 15656 17748 15703 17812
rect 15767 17748 15783 17812
rect 15656 17732 15783 17748
rect 15656 17668 15703 17732
rect 15767 17668 15783 17732
rect 15656 17652 15783 17668
rect 15656 17588 15703 17652
rect 15767 17588 15783 17652
rect 15656 17572 15783 17588
rect 15656 17508 15703 17572
rect 15767 17508 15783 17572
rect 15656 17492 15783 17508
rect 15656 17428 15703 17492
rect 15767 17428 15783 17492
rect 15656 17412 15783 17428
rect 15656 17348 15703 17412
rect 15767 17348 15783 17412
rect 15656 17332 15783 17348
rect 15656 17268 15703 17332
rect 15767 17268 15783 17332
rect 15656 17252 15783 17268
rect 15656 17188 15703 17252
rect 15767 17188 15783 17252
rect 15656 17172 15783 17188
rect 15656 17108 15703 17172
rect 15767 17108 15783 17172
rect 15656 17092 15783 17108
rect 15656 17028 15703 17092
rect 15767 17028 15783 17092
rect 15656 17012 15783 17028
rect 15656 16948 15703 17012
rect 15767 16948 15783 17012
rect 15656 16932 15783 16948
rect 15656 16868 15703 16932
rect 15767 16868 15783 16932
rect 15656 16852 15783 16868
rect 15656 16788 15703 16852
rect 15767 16788 15783 16852
rect 15656 16772 15783 16788
rect 15656 16708 15703 16772
rect 15767 16708 15783 16772
rect 15656 16692 15783 16708
rect 15656 16628 15703 16692
rect 15767 16628 15783 16692
rect 15656 16612 15783 16628
rect 15656 16548 15703 16612
rect 15767 16548 15783 16612
rect 15656 16532 15783 16548
rect 15656 16468 15703 16532
rect 15767 16468 15783 16532
rect 15656 16452 15783 16468
rect 15656 16388 15703 16452
rect 15767 16388 15783 16452
rect 15656 16372 15783 16388
rect 15656 16308 15703 16372
rect 15767 16308 15783 16372
rect 15656 16292 15783 16308
rect 15656 16228 15703 16292
rect 15767 16228 15783 16292
rect 15656 16212 15783 16228
rect 15656 16148 15703 16212
rect 15767 16148 15783 16212
rect 15656 16132 15783 16148
rect 15656 16068 15703 16132
rect 15767 16068 15783 16132
rect 15656 16052 15783 16068
rect 15656 15988 15703 16052
rect 15767 15988 15783 16052
rect 15656 15972 15783 15988
rect 9337 15892 9464 15908
rect 9337 15828 9384 15892
rect 9448 15828 9464 15892
rect 9337 15812 9464 15828
rect 9337 15688 9441 15812
rect 9337 15672 9464 15688
rect 9337 15608 9384 15672
rect 9448 15608 9464 15672
rect 9337 15592 9464 15608
rect 3018 15512 3145 15528
rect 3018 15448 3065 15512
rect 3129 15448 3145 15512
rect 3018 15432 3145 15448
rect 3018 15368 3065 15432
rect 3129 15368 3145 15432
rect 3018 15352 3145 15368
rect 3018 15288 3065 15352
rect 3129 15288 3145 15352
rect 3018 15272 3145 15288
rect 3018 15208 3065 15272
rect 3129 15208 3145 15272
rect 3018 15192 3145 15208
rect 3018 15128 3065 15192
rect 3129 15128 3145 15192
rect 3018 15112 3145 15128
rect 3018 15048 3065 15112
rect 3129 15048 3145 15112
rect 3018 15032 3145 15048
rect 3018 14968 3065 15032
rect 3129 14968 3145 15032
rect 3018 14952 3145 14968
rect 3018 14888 3065 14952
rect 3129 14888 3145 14952
rect 3018 14872 3145 14888
rect 3018 14808 3065 14872
rect 3129 14808 3145 14872
rect 3018 14792 3145 14808
rect 3018 14728 3065 14792
rect 3129 14728 3145 14792
rect 3018 14712 3145 14728
rect 3018 14648 3065 14712
rect 3129 14648 3145 14712
rect 3018 14632 3145 14648
rect 3018 14568 3065 14632
rect 3129 14568 3145 14632
rect 3018 14552 3145 14568
rect 3018 14488 3065 14552
rect 3129 14488 3145 14552
rect 3018 14472 3145 14488
rect 3018 14408 3065 14472
rect 3129 14408 3145 14472
rect 3018 14392 3145 14408
rect 3018 14328 3065 14392
rect 3129 14328 3145 14392
rect 3018 14312 3145 14328
rect 3018 14248 3065 14312
rect 3129 14248 3145 14312
rect 3018 14232 3145 14248
rect 3018 14168 3065 14232
rect 3129 14168 3145 14232
rect 3018 14152 3145 14168
rect 3018 14088 3065 14152
rect 3129 14088 3145 14152
rect 3018 14072 3145 14088
rect 3018 14008 3065 14072
rect 3129 14008 3145 14072
rect 3018 13992 3145 14008
rect 3018 13928 3065 13992
rect 3129 13928 3145 13992
rect 3018 13912 3145 13928
rect 3018 13848 3065 13912
rect 3129 13848 3145 13912
rect 3018 13832 3145 13848
rect 3018 13768 3065 13832
rect 3129 13768 3145 13832
rect 3018 13752 3145 13768
rect 3018 13688 3065 13752
rect 3129 13688 3145 13752
rect 3018 13672 3145 13688
rect 3018 13608 3065 13672
rect 3129 13608 3145 13672
rect 3018 13592 3145 13608
rect 3018 13528 3065 13592
rect 3129 13528 3145 13592
rect 3018 13512 3145 13528
rect 3018 13448 3065 13512
rect 3129 13448 3145 13512
rect 3018 13432 3145 13448
rect 3018 13368 3065 13432
rect 3129 13368 3145 13432
rect 3018 13352 3145 13368
rect 3018 13288 3065 13352
rect 3129 13288 3145 13352
rect 3018 13272 3145 13288
rect 3018 13208 3065 13272
rect 3129 13208 3145 13272
rect 3018 13192 3145 13208
rect 3018 13128 3065 13192
rect 3129 13128 3145 13192
rect 3018 13112 3145 13128
rect 3018 13048 3065 13112
rect 3129 13048 3145 13112
rect 3018 13032 3145 13048
rect 3018 12968 3065 13032
rect 3129 12968 3145 13032
rect 3018 12952 3145 12968
rect 3018 12888 3065 12952
rect 3129 12888 3145 12952
rect 3018 12872 3145 12888
rect 3018 12808 3065 12872
rect 3129 12808 3145 12872
rect 3018 12792 3145 12808
rect 3018 12728 3065 12792
rect 3129 12728 3145 12792
rect 3018 12712 3145 12728
rect 3018 12648 3065 12712
rect 3129 12648 3145 12712
rect 3018 12632 3145 12648
rect 3018 12568 3065 12632
rect 3129 12568 3145 12632
rect 3018 12552 3145 12568
rect 3018 12488 3065 12552
rect 3129 12488 3145 12552
rect 3018 12472 3145 12488
rect 3018 12408 3065 12472
rect 3129 12408 3145 12472
rect 3018 12392 3145 12408
rect 3018 12328 3065 12392
rect 3129 12328 3145 12392
rect 3018 12312 3145 12328
rect 3018 12248 3065 12312
rect 3129 12248 3145 12312
rect 3018 12232 3145 12248
rect 3018 12168 3065 12232
rect 3129 12168 3145 12232
rect 3018 12152 3145 12168
rect 3018 12088 3065 12152
rect 3129 12088 3145 12152
rect 3018 12072 3145 12088
rect 3018 12008 3065 12072
rect 3129 12008 3145 12072
rect 3018 11992 3145 12008
rect 3018 11928 3065 11992
rect 3129 11928 3145 11992
rect 3018 11912 3145 11928
rect 3018 11848 3065 11912
rect 3129 11848 3145 11912
rect 3018 11832 3145 11848
rect 3018 11768 3065 11832
rect 3129 11768 3145 11832
rect 3018 11752 3145 11768
rect 3018 11688 3065 11752
rect 3129 11688 3145 11752
rect 3018 11672 3145 11688
rect 3018 11608 3065 11672
rect 3129 11608 3145 11672
rect 3018 11592 3145 11608
rect 3018 11528 3065 11592
rect 3129 11528 3145 11592
rect 3018 11512 3145 11528
rect 3018 11448 3065 11512
rect 3129 11448 3145 11512
rect 3018 11432 3145 11448
rect 3018 11368 3065 11432
rect 3129 11368 3145 11432
rect 3018 11352 3145 11368
rect 3018 11288 3065 11352
rect 3129 11288 3145 11352
rect 3018 11272 3145 11288
rect 3018 11208 3065 11272
rect 3129 11208 3145 11272
rect 3018 11192 3145 11208
rect 3018 11128 3065 11192
rect 3129 11128 3145 11192
rect 3018 11112 3145 11128
rect 3018 11048 3065 11112
rect 3129 11048 3145 11112
rect 3018 11032 3145 11048
rect 3018 10968 3065 11032
rect 3129 10968 3145 11032
rect 3018 10952 3145 10968
rect 3018 10888 3065 10952
rect 3129 10888 3145 10952
rect 3018 10872 3145 10888
rect 3018 10808 3065 10872
rect 3129 10808 3145 10872
rect 3018 10792 3145 10808
rect 3018 10728 3065 10792
rect 3129 10728 3145 10792
rect 3018 10712 3145 10728
rect 3018 10648 3065 10712
rect 3129 10648 3145 10712
rect 3018 10632 3145 10648
rect 3018 10568 3065 10632
rect 3129 10568 3145 10632
rect 3018 10552 3145 10568
rect 3018 10488 3065 10552
rect 3129 10488 3145 10552
rect 3018 10472 3145 10488
rect 3018 10408 3065 10472
rect 3129 10408 3145 10472
rect 3018 10392 3145 10408
rect 3018 10328 3065 10392
rect 3129 10328 3145 10392
rect 3018 10312 3145 10328
rect 3018 10248 3065 10312
rect 3129 10248 3145 10312
rect 3018 10232 3145 10248
rect 3018 10168 3065 10232
rect 3129 10168 3145 10232
rect 3018 10152 3145 10168
rect 3018 10088 3065 10152
rect 3129 10088 3145 10152
rect 3018 10072 3145 10088
rect 3018 10008 3065 10072
rect 3129 10008 3145 10072
rect 3018 9992 3145 10008
rect 3018 9928 3065 9992
rect 3129 9928 3145 9992
rect 3018 9912 3145 9928
rect 3018 9848 3065 9912
rect 3129 9848 3145 9912
rect 3018 9832 3145 9848
rect 3018 9768 3065 9832
rect 3129 9768 3145 9832
rect 3018 9752 3145 9768
rect 3018 9688 3065 9752
rect 3129 9688 3145 9752
rect 3018 9672 3145 9688
rect -3301 9592 -3174 9608
rect -3301 9528 -3254 9592
rect -3190 9528 -3174 9592
rect -3301 9512 -3174 9528
rect -3301 9388 -3197 9512
rect -3301 9372 -3174 9388
rect -3301 9308 -3254 9372
rect -3190 9308 -3174 9372
rect -3301 9292 -3174 9308
rect -9620 9212 -9493 9228
rect -9620 9148 -9573 9212
rect -9509 9148 -9493 9212
rect -9620 9132 -9493 9148
rect -9620 9068 -9573 9132
rect -9509 9068 -9493 9132
rect -9620 9052 -9493 9068
rect -9620 8988 -9573 9052
rect -9509 8988 -9493 9052
rect -9620 8972 -9493 8988
rect -9620 8908 -9573 8972
rect -9509 8908 -9493 8972
rect -9620 8892 -9493 8908
rect -9620 8828 -9573 8892
rect -9509 8828 -9493 8892
rect -9620 8812 -9493 8828
rect -9620 8748 -9573 8812
rect -9509 8748 -9493 8812
rect -9620 8732 -9493 8748
rect -9620 8668 -9573 8732
rect -9509 8668 -9493 8732
rect -9620 8652 -9493 8668
rect -9620 8588 -9573 8652
rect -9509 8588 -9493 8652
rect -9620 8572 -9493 8588
rect -9620 8508 -9573 8572
rect -9509 8508 -9493 8572
rect -9620 8492 -9493 8508
rect -9620 8428 -9573 8492
rect -9509 8428 -9493 8492
rect -9620 8412 -9493 8428
rect -9620 8348 -9573 8412
rect -9509 8348 -9493 8412
rect -9620 8332 -9493 8348
rect -9620 8268 -9573 8332
rect -9509 8268 -9493 8332
rect -9620 8252 -9493 8268
rect -9620 8188 -9573 8252
rect -9509 8188 -9493 8252
rect -9620 8172 -9493 8188
rect -9620 8108 -9573 8172
rect -9509 8108 -9493 8172
rect -9620 8092 -9493 8108
rect -9620 8028 -9573 8092
rect -9509 8028 -9493 8092
rect -9620 8012 -9493 8028
rect -9620 7948 -9573 8012
rect -9509 7948 -9493 8012
rect -9620 7932 -9493 7948
rect -9620 7868 -9573 7932
rect -9509 7868 -9493 7932
rect -9620 7852 -9493 7868
rect -9620 7788 -9573 7852
rect -9509 7788 -9493 7852
rect -9620 7772 -9493 7788
rect -9620 7708 -9573 7772
rect -9509 7708 -9493 7772
rect -9620 7692 -9493 7708
rect -9620 7628 -9573 7692
rect -9509 7628 -9493 7692
rect -9620 7612 -9493 7628
rect -9620 7548 -9573 7612
rect -9509 7548 -9493 7612
rect -9620 7532 -9493 7548
rect -9620 7468 -9573 7532
rect -9509 7468 -9493 7532
rect -9620 7452 -9493 7468
rect -9620 7388 -9573 7452
rect -9509 7388 -9493 7452
rect -9620 7372 -9493 7388
rect -9620 7308 -9573 7372
rect -9509 7308 -9493 7372
rect -9620 7292 -9493 7308
rect -9620 7228 -9573 7292
rect -9509 7228 -9493 7292
rect -9620 7212 -9493 7228
rect -9620 7148 -9573 7212
rect -9509 7148 -9493 7212
rect -9620 7132 -9493 7148
rect -9620 7068 -9573 7132
rect -9509 7068 -9493 7132
rect -9620 7052 -9493 7068
rect -9620 6988 -9573 7052
rect -9509 6988 -9493 7052
rect -9620 6972 -9493 6988
rect -9620 6908 -9573 6972
rect -9509 6908 -9493 6972
rect -9620 6892 -9493 6908
rect -9620 6828 -9573 6892
rect -9509 6828 -9493 6892
rect -9620 6812 -9493 6828
rect -9620 6748 -9573 6812
rect -9509 6748 -9493 6812
rect -9620 6732 -9493 6748
rect -9620 6668 -9573 6732
rect -9509 6668 -9493 6732
rect -9620 6652 -9493 6668
rect -9620 6588 -9573 6652
rect -9509 6588 -9493 6652
rect -9620 6572 -9493 6588
rect -9620 6508 -9573 6572
rect -9509 6508 -9493 6572
rect -9620 6492 -9493 6508
rect -9620 6428 -9573 6492
rect -9509 6428 -9493 6492
rect -9620 6412 -9493 6428
rect -9620 6348 -9573 6412
rect -9509 6348 -9493 6412
rect -9620 6332 -9493 6348
rect -9620 6268 -9573 6332
rect -9509 6268 -9493 6332
rect -9620 6252 -9493 6268
rect -9620 6188 -9573 6252
rect -9509 6188 -9493 6252
rect -9620 6172 -9493 6188
rect -9620 6108 -9573 6172
rect -9509 6108 -9493 6172
rect -9620 6092 -9493 6108
rect -9620 6028 -9573 6092
rect -9509 6028 -9493 6092
rect -9620 6012 -9493 6028
rect -9620 5948 -9573 6012
rect -9509 5948 -9493 6012
rect -9620 5932 -9493 5948
rect -9620 5868 -9573 5932
rect -9509 5868 -9493 5932
rect -9620 5852 -9493 5868
rect -9620 5788 -9573 5852
rect -9509 5788 -9493 5852
rect -9620 5772 -9493 5788
rect -9620 5708 -9573 5772
rect -9509 5708 -9493 5772
rect -9620 5692 -9493 5708
rect -9620 5628 -9573 5692
rect -9509 5628 -9493 5692
rect -9620 5612 -9493 5628
rect -9620 5548 -9573 5612
rect -9509 5548 -9493 5612
rect -9620 5532 -9493 5548
rect -9620 5468 -9573 5532
rect -9509 5468 -9493 5532
rect -9620 5452 -9493 5468
rect -9620 5388 -9573 5452
rect -9509 5388 -9493 5452
rect -9620 5372 -9493 5388
rect -9620 5308 -9573 5372
rect -9509 5308 -9493 5372
rect -9620 5292 -9493 5308
rect -9620 5228 -9573 5292
rect -9509 5228 -9493 5292
rect -9620 5212 -9493 5228
rect -9620 5148 -9573 5212
rect -9509 5148 -9493 5212
rect -9620 5132 -9493 5148
rect -9620 5068 -9573 5132
rect -9509 5068 -9493 5132
rect -9620 5052 -9493 5068
rect -9620 4988 -9573 5052
rect -9509 4988 -9493 5052
rect -9620 4972 -9493 4988
rect -9620 4908 -9573 4972
rect -9509 4908 -9493 4972
rect -9620 4892 -9493 4908
rect -9620 4828 -9573 4892
rect -9509 4828 -9493 4892
rect -9620 4812 -9493 4828
rect -9620 4748 -9573 4812
rect -9509 4748 -9493 4812
rect -9620 4732 -9493 4748
rect -9620 4668 -9573 4732
rect -9509 4668 -9493 4732
rect -9620 4652 -9493 4668
rect -9620 4588 -9573 4652
rect -9509 4588 -9493 4652
rect -9620 4572 -9493 4588
rect -9620 4508 -9573 4572
rect -9509 4508 -9493 4572
rect -9620 4492 -9493 4508
rect -9620 4428 -9573 4492
rect -9509 4428 -9493 4492
rect -9620 4412 -9493 4428
rect -9620 4348 -9573 4412
rect -9509 4348 -9493 4412
rect -9620 4332 -9493 4348
rect -9620 4268 -9573 4332
rect -9509 4268 -9493 4332
rect -9620 4252 -9493 4268
rect -9620 4188 -9573 4252
rect -9509 4188 -9493 4252
rect -9620 4172 -9493 4188
rect -9620 4108 -9573 4172
rect -9509 4108 -9493 4172
rect -9620 4092 -9493 4108
rect -9620 4028 -9573 4092
rect -9509 4028 -9493 4092
rect -9620 4012 -9493 4028
rect -9620 3948 -9573 4012
rect -9509 3948 -9493 4012
rect -9620 3932 -9493 3948
rect -9620 3868 -9573 3932
rect -9509 3868 -9493 3932
rect -9620 3852 -9493 3868
rect -9620 3788 -9573 3852
rect -9509 3788 -9493 3852
rect -9620 3772 -9493 3788
rect -9620 3708 -9573 3772
rect -9509 3708 -9493 3772
rect -9620 3692 -9493 3708
rect -9620 3628 -9573 3692
rect -9509 3628 -9493 3692
rect -9620 3612 -9493 3628
rect -9620 3548 -9573 3612
rect -9509 3548 -9493 3612
rect -9620 3532 -9493 3548
rect -9620 3468 -9573 3532
rect -9509 3468 -9493 3532
rect -9620 3452 -9493 3468
rect -9620 3388 -9573 3452
rect -9509 3388 -9493 3452
rect -9620 3372 -9493 3388
rect -15939 3292 -15812 3308
rect -15939 3228 -15892 3292
rect -15828 3228 -15812 3292
rect -15939 3212 -15812 3228
rect -15939 3088 -15835 3212
rect -15939 3072 -15812 3088
rect -15939 3008 -15892 3072
rect -15828 3008 -15812 3072
rect -15939 2992 -15812 3008
rect -22258 2912 -22131 2928
rect -22258 2848 -22211 2912
rect -22147 2848 -22131 2912
rect -22258 2832 -22131 2848
rect -22258 2768 -22211 2832
rect -22147 2768 -22131 2832
rect -22258 2752 -22131 2768
rect -22258 2688 -22211 2752
rect -22147 2688 -22131 2752
rect -22258 2672 -22131 2688
rect -22258 2608 -22211 2672
rect -22147 2608 -22131 2672
rect -22258 2592 -22131 2608
rect -22258 2528 -22211 2592
rect -22147 2528 -22131 2592
rect -22258 2512 -22131 2528
rect -22258 2448 -22211 2512
rect -22147 2448 -22131 2512
rect -22258 2432 -22131 2448
rect -22258 2368 -22211 2432
rect -22147 2368 -22131 2432
rect -22258 2352 -22131 2368
rect -22258 2288 -22211 2352
rect -22147 2288 -22131 2352
rect -22258 2272 -22131 2288
rect -22258 2208 -22211 2272
rect -22147 2208 -22131 2272
rect -22258 2192 -22131 2208
rect -22258 2128 -22211 2192
rect -22147 2128 -22131 2192
rect -22258 2112 -22131 2128
rect -22258 2048 -22211 2112
rect -22147 2048 -22131 2112
rect -22258 2032 -22131 2048
rect -22258 1968 -22211 2032
rect -22147 1968 -22131 2032
rect -22258 1952 -22131 1968
rect -22258 1888 -22211 1952
rect -22147 1888 -22131 1952
rect -22258 1872 -22131 1888
rect -22258 1808 -22211 1872
rect -22147 1808 -22131 1872
rect -22258 1792 -22131 1808
rect -22258 1728 -22211 1792
rect -22147 1728 -22131 1792
rect -22258 1712 -22131 1728
rect -22258 1648 -22211 1712
rect -22147 1648 -22131 1712
rect -22258 1632 -22131 1648
rect -22258 1568 -22211 1632
rect -22147 1568 -22131 1632
rect -22258 1552 -22131 1568
rect -22258 1488 -22211 1552
rect -22147 1488 -22131 1552
rect -22258 1472 -22131 1488
rect -22258 1408 -22211 1472
rect -22147 1408 -22131 1472
rect -22258 1392 -22131 1408
rect -22258 1328 -22211 1392
rect -22147 1328 -22131 1392
rect -22258 1312 -22131 1328
rect -22258 1248 -22211 1312
rect -22147 1248 -22131 1312
rect -22258 1232 -22131 1248
rect -22258 1168 -22211 1232
rect -22147 1168 -22131 1232
rect -22258 1152 -22131 1168
rect -22258 1088 -22211 1152
rect -22147 1088 -22131 1152
rect -22258 1072 -22131 1088
rect -22258 1008 -22211 1072
rect -22147 1008 -22131 1072
rect -22258 992 -22131 1008
rect -22258 928 -22211 992
rect -22147 928 -22131 992
rect -22258 912 -22131 928
rect -22258 848 -22211 912
rect -22147 848 -22131 912
rect -22258 832 -22131 848
rect -22258 768 -22211 832
rect -22147 768 -22131 832
rect -22258 752 -22131 768
rect -22258 688 -22211 752
rect -22147 688 -22131 752
rect -22258 672 -22131 688
rect -22258 608 -22211 672
rect -22147 608 -22131 672
rect -22258 592 -22131 608
rect -22258 528 -22211 592
rect -22147 528 -22131 592
rect -22258 512 -22131 528
rect -22258 448 -22211 512
rect -22147 448 -22131 512
rect -22258 432 -22131 448
rect -22258 368 -22211 432
rect -22147 368 -22131 432
rect -22258 352 -22131 368
rect -22258 288 -22211 352
rect -22147 288 -22131 352
rect -22258 272 -22131 288
rect -22258 208 -22211 272
rect -22147 208 -22131 272
rect -22258 192 -22131 208
rect -22258 128 -22211 192
rect -22147 128 -22131 192
rect -22258 112 -22131 128
rect -22258 48 -22211 112
rect -22147 48 -22131 112
rect -22258 32 -22131 48
rect -22258 -32 -22211 32
rect -22147 -32 -22131 32
rect -22258 -48 -22131 -32
rect -22258 -112 -22211 -48
rect -22147 -112 -22131 -48
rect -22258 -128 -22131 -112
rect -22258 -192 -22211 -128
rect -22147 -192 -22131 -128
rect -22258 -208 -22131 -192
rect -22258 -272 -22211 -208
rect -22147 -272 -22131 -208
rect -22258 -288 -22131 -272
rect -22258 -352 -22211 -288
rect -22147 -352 -22131 -288
rect -22258 -368 -22131 -352
rect -22258 -432 -22211 -368
rect -22147 -432 -22131 -368
rect -22258 -448 -22131 -432
rect -22258 -512 -22211 -448
rect -22147 -512 -22131 -448
rect -22258 -528 -22131 -512
rect -22258 -592 -22211 -528
rect -22147 -592 -22131 -528
rect -22258 -608 -22131 -592
rect -22258 -672 -22211 -608
rect -22147 -672 -22131 -608
rect -22258 -688 -22131 -672
rect -22258 -752 -22211 -688
rect -22147 -752 -22131 -688
rect -22258 -768 -22131 -752
rect -22258 -832 -22211 -768
rect -22147 -832 -22131 -768
rect -22258 -848 -22131 -832
rect -22258 -912 -22211 -848
rect -22147 -912 -22131 -848
rect -22258 -928 -22131 -912
rect -22258 -992 -22211 -928
rect -22147 -992 -22131 -928
rect -22258 -1008 -22131 -992
rect -22258 -1072 -22211 -1008
rect -22147 -1072 -22131 -1008
rect -22258 -1088 -22131 -1072
rect -22258 -1152 -22211 -1088
rect -22147 -1152 -22131 -1088
rect -22258 -1168 -22131 -1152
rect -22258 -1232 -22211 -1168
rect -22147 -1232 -22131 -1168
rect -22258 -1248 -22131 -1232
rect -22258 -1312 -22211 -1248
rect -22147 -1312 -22131 -1248
rect -22258 -1328 -22131 -1312
rect -22258 -1392 -22211 -1328
rect -22147 -1392 -22131 -1328
rect -22258 -1408 -22131 -1392
rect -22258 -1472 -22211 -1408
rect -22147 -1472 -22131 -1408
rect -22258 -1488 -22131 -1472
rect -22258 -1552 -22211 -1488
rect -22147 -1552 -22131 -1488
rect -22258 -1568 -22131 -1552
rect -22258 -1632 -22211 -1568
rect -22147 -1632 -22131 -1568
rect -22258 -1648 -22131 -1632
rect -22258 -1712 -22211 -1648
rect -22147 -1712 -22131 -1648
rect -22258 -1728 -22131 -1712
rect -22258 -1792 -22211 -1728
rect -22147 -1792 -22131 -1728
rect -22258 -1808 -22131 -1792
rect -22258 -1872 -22211 -1808
rect -22147 -1872 -22131 -1808
rect -22258 -1888 -22131 -1872
rect -22258 -1952 -22211 -1888
rect -22147 -1952 -22131 -1888
rect -22258 -1968 -22131 -1952
rect -22258 -2032 -22211 -1968
rect -22147 -2032 -22131 -1968
rect -22258 -2048 -22131 -2032
rect -22258 -2112 -22211 -2048
rect -22147 -2112 -22131 -2048
rect -22258 -2128 -22131 -2112
rect -22258 -2192 -22211 -2128
rect -22147 -2192 -22131 -2128
rect -22258 -2208 -22131 -2192
rect -22258 -2272 -22211 -2208
rect -22147 -2272 -22131 -2208
rect -22258 -2288 -22131 -2272
rect -22258 -2352 -22211 -2288
rect -22147 -2352 -22131 -2288
rect -22258 -2368 -22131 -2352
rect -22258 -2432 -22211 -2368
rect -22147 -2432 -22131 -2368
rect -22258 -2448 -22131 -2432
rect -22258 -2512 -22211 -2448
rect -22147 -2512 -22131 -2448
rect -22258 -2528 -22131 -2512
rect -22258 -2592 -22211 -2528
rect -22147 -2592 -22131 -2528
rect -22258 -2608 -22131 -2592
rect -22258 -2672 -22211 -2608
rect -22147 -2672 -22131 -2608
rect -22258 -2688 -22131 -2672
rect -22258 -2752 -22211 -2688
rect -22147 -2752 -22131 -2688
rect -22258 -2768 -22131 -2752
rect -22258 -2832 -22211 -2768
rect -22147 -2832 -22131 -2768
rect -22258 -2848 -22131 -2832
rect -22258 -2912 -22211 -2848
rect -22147 -2912 -22131 -2848
rect -22258 -2928 -22131 -2912
rect -28577 -3008 -28450 -2992
rect -28577 -3072 -28530 -3008
rect -28466 -3072 -28450 -3008
rect -28577 -3088 -28450 -3072
rect -28577 -3212 -28473 -3088
rect -28577 -3228 -28450 -3212
rect -28577 -3292 -28530 -3228
rect -28466 -3292 -28450 -3228
rect -28577 -3308 -28450 -3292
rect -34896 -3388 -34769 -3372
rect -34896 -3452 -34849 -3388
rect -34785 -3452 -34769 -3388
rect -34896 -3468 -34769 -3452
rect -34896 -3532 -34849 -3468
rect -34785 -3532 -34769 -3468
rect -34896 -3548 -34769 -3532
rect -34896 -3612 -34849 -3548
rect -34785 -3612 -34769 -3548
rect -34896 -3628 -34769 -3612
rect -34896 -3692 -34849 -3628
rect -34785 -3692 -34769 -3628
rect -34896 -3708 -34769 -3692
rect -34896 -3772 -34849 -3708
rect -34785 -3772 -34769 -3708
rect -34896 -3788 -34769 -3772
rect -34896 -3852 -34849 -3788
rect -34785 -3852 -34769 -3788
rect -34896 -3868 -34769 -3852
rect -34896 -3932 -34849 -3868
rect -34785 -3932 -34769 -3868
rect -34896 -3948 -34769 -3932
rect -34896 -4012 -34849 -3948
rect -34785 -4012 -34769 -3948
rect -34896 -4028 -34769 -4012
rect -34896 -4092 -34849 -4028
rect -34785 -4092 -34769 -4028
rect -34896 -4108 -34769 -4092
rect -34896 -4172 -34849 -4108
rect -34785 -4172 -34769 -4108
rect -34896 -4188 -34769 -4172
rect -34896 -4252 -34849 -4188
rect -34785 -4252 -34769 -4188
rect -34896 -4268 -34769 -4252
rect -34896 -4332 -34849 -4268
rect -34785 -4332 -34769 -4268
rect -34896 -4348 -34769 -4332
rect -34896 -4412 -34849 -4348
rect -34785 -4412 -34769 -4348
rect -34896 -4428 -34769 -4412
rect -34896 -4492 -34849 -4428
rect -34785 -4492 -34769 -4428
rect -34896 -4508 -34769 -4492
rect -34896 -4572 -34849 -4508
rect -34785 -4572 -34769 -4508
rect -34896 -4588 -34769 -4572
rect -34896 -4652 -34849 -4588
rect -34785 -4652 -34769 -4588
rect -34896 -4668 -34769 -4652
rect -34896 -4732 -34849 -4668
rect -34785 -4732 -34769 -4668
rect -34896 -4748 -34769 -4732
rect -34896 -4812 -34849 -4748
rect -34785 -4812 -34769 -4748
rect -34896 -4828 -34769 -4812
rect -34896 -4892 -34849 -4828
rect -34785 -4892 -34769 -4828
rect -34896 -4908 -34769 -4892
rect -34896 -4972 -34849 -4908
rect -34785 -4972 -34769 -4908
rect -34896 -4988 -34769 -4972
rect -34896 -5052 -34849 -4988
rect -34785 -5052 -34769 -4988
rect -34896 -5068 -34769 -5052
rect -34896 -5132 -34849 -5068
rect -34785 -5132 -34769 -5068
rect -34896 -5148 -34769 -5132
rect -34896 -5212 -34849 -5148
rect -34785 -5212 -34769 -5148
rect -34896 -5228 -34769 -5212
rect -34896 -5292 -34849 -5228
rect -34785 -5292 -34769 -5228
rect -34896 -5308 -34769 -5292
rect -34896 -5372 -34849 -5308
rect -34785 -5372 -34769 -5308
rect -34896 -5388 -34769 -5372
rect -34896 -5452 -34849 -5388
rect -34785 -5452 -34769 -5388
rect -34896 -5468 -34769 -5452
rect -34896 -5532 -34849 -5468
rect -34785 -5532 -34769 -5468
rect -34896 -5548 -34769 -5532
rect -34896 -5612 -34849 -5548
rect -34785 -5612 -34769 -5548
rect -34896 -5628 -34769 -5612
rect -34896 -5692 -34849 -5628
rect -34785 -5692 -34769 -5628
rect -34896 -5708 -34769 -5692
rect -34896 -5772 -34849 -5708
rect -34785 -5772 -34769 -5708
rect -34896 -5788 -34769 -5772
rect -34896 -5852 -34849 -5788
rect -34785 -5852 -34769 -5788
rect -34896 -5868 -34769 -5852
rect -34896 -5932 -34849 -5868
rect -34785 -5932 -34769 -5868
rect -34896 -5948 -34769 -5932
rect -34896 -6012 -34849 -5948
rect -34785 -6012 -34769 -5948
rect -34896 -6028 -34769 -6012
rect -34896 -6092 -34849 -6028
rect -34785 -6092 -34769 -6028
rect -34896 -6108 -34769 -6092
rect -34896 -6172 -34849 -6108
rect -34785 -6172 -34769 -6108
rect -34896 -6188 -34769 -6172
rect -34896 -6252 -34849 -6188
rect -34785 -6252 -34769 -6188
rect -34896 -6268 -34769 -6252
rect -34896 -6332 -34849 -6268
rect -34785 -6332 -34769 -6268
rect -34896 -6348 -34769 -6332
rect -34896 -6412 -34849 -6348
rect -34785 -6412 -34769 -6348
rect -34896 -6428 -34769 -6412
rect -34896 -6492 -34849 -6428
rect -34785 -6492 -34769 -6428
rect -34896 -6508 -34769 -6492
rect -34896 -6572 -34849 -6508
rect -34785 -6572 -34769 -6508
rect -34896 -6588 -34769 -6572
rect -34896 -6652 -34849 -6588
rect -34785 -6652 -34769 -6588
rect -34896 -6668 -34769 -6652
rect -34896 -6732 -34849 -6668
rect -34785 -6732 -34769 -6668
rect -34896 -6748 -34769 -6732
rect -34896 -6812 -34849 -6748
rect -34785 -6812 -34769 -6748
rect -34896 -6828 -34769 -6812
rect -34896 -6892 -34849 -6828
rect -34785 -6892 -34769 -6828
rect -34896 -6908 -34769 -6892
rect -34896 -6972 -34849 -6908
rect -34785 -6972 -34769 -6908
rect -34896 -6988 -34769 -6972
rect -34896 -7052 -34849 -6988
rect -34785 -7052 -34769 -6988
rect -34896 -7068 -34769 -7052
rect -34896 -7132 -34849 -7068
rect -34785 -7132 -34769 -7068
rect -34896 -7148 -34769 -7132
rect -34896 -7212 -34849 -7148
rect -34785 -7212 -34769 -7148
rect -34896 -7228 -34769 -7212
rect -34896 -7292 -34849 -7228
rect -34785 -7292 -34769 -7228
rect -34896 -7308 -34769 -7292
rect -34896 -7372 -34849 -7308
rect -34785 -7372 -34769 -7308
rect -34896 -7388 -34769 -7372
rect -34896 -7452 -34849 -7388
rect -34785 -7452 -34769 -7388
rect -34896 -7468 -34769 -7452
rect -34896 -7532 -34849 -7468
rect -34785 -7532 -34769 -7468
rect -34896 -7548 -34769 -7532
rect -34896 -7612 -34849 -7548
rect -34785 -7612 -34769 -7548
rect -34896 -7628 -34769 -7612
rect -34896 -7692 -34849 -7628
rect -34785 -7692 -34769 -7628
rect -34896 -7708 -34769 -7692
rect -34896 -7772 -34849 -7708
rect -34785 -7772 -34769 -7708
rect -34896 -7788 -34769 -7772
rect -34896 -7852 -34849 -7788
rect -34785 -7852 -34769 -7788
rect -34896 -7868 -34769 -7852
rect -34896 -7932 -34849 -7868
rect -34785 -7932 -34769 -7868
rect -34896 -7948 -34769 -7932
rect -34896 -8012 -34849 -7948
rect -34785 -8012 -34769 -7948
rect -34896 -8028 -34769 -8012
rect -34896 -8092 -34849 -8028
rect -34785 -8092 -34769 -8028
rect -34896 -8108 -34769 -8092
rect -34896 -8172 -34849 -8108
rect -34785 -8172 -34769 -8108
rect -34896 -8188 -34769 -8172
rect -34896 -8252 -34849 -8188
rect -34785 -8252 -34769 -8188
rect -34896 -8268 -34769 -8252
rect -34896 -8332 -34849 -8268
rect -34785 -8332 -34769 -8268
rect -34896 -8348 -34769 -8332
rect -34896 -8412 -34849 -8348
rect -34785 -8412 -34769 -8348
rect -34896 -8428 -34769 -8412
rect -34896 -8492 -34849 -8428
rect -34785 -8492 -34769 -8428
rect -34896 -8508 -34769 -8492
rect -34896 -8572 -34849 -8508
rect -34785 -8572 -34769 -8508
rect -34896 -8588 -34769 -8572
rect -34896 -8652 -34849 -8588
rect -34785 -8652 -34769 -8588
rect -34896 -8668 -34769 -8652
rect -34896 -8732 -34849 -8668
rect -34785 -8732 -34769 -8668
rect -34896 -8748 -34769 -8732
rect -34896 -8812 -34849 -8748
rect -34785 -8812 -34769 -8748
rect -34896 -8828 -34769 -8812
rect -34896 -8892 -34849 -8828
rect -34785 -8892 -34769 -8828
rect -34896 -8908 -34769 -8892
rect -34896 -8972 -34849 -8908
rect -34785 -8972 -34769 -8908
rect -34896 -8988 -34769 -8972
rect -34896 -9052 -34849 -8988
rect -34785 -9052 -34769 -8988
rect -34896 -9068 -34769 -9052
rect -34896 -9132 -34849 -9068
rect -34785 -9132 -34769 -9068
rect -34896 -9148 -34769 -9132
rect -34896 -9212 -34849 -9148
rect -34785 -9212 -34769 -9148
rect -34896 -9228 -34769 -9212
rect -41215 -9308 -41088 -9292
rect -41215 -9372 -41168 -9308
rect -41104 -9372 -41088 -9308
rect -41215 -9388 -41088 -9372
rect -41215 -9512 -41111 -9388
rect -41215 -9528 -41088 -9512
rect -41215 -9592 -41168 -9528
rect -41104 -9592 -41088 -9528
rect -41215 -9608 -41088 -9592
rect -47244 -9648 -41322 -9639
rect -47244 -15552 -47235 -9648
rect -41331 -15552 -41322 -9648
rect -47244 -15561 -41322 -15552
rect -41215 -9672 -41168 -9608
rect -41104 -9672 -41088 -9608
rect -38016 -9639 -37912 -9261
rect -34896 -9292 -34849 -9228
rect -34785 -9292 -34769 -9228
rect -34606 -3348 -28684 -3339
rect -34606 -9252 -34597 -3348
rect -28693 -9252 -28684 -3348
rect -34606 -9261 -28684 -9252
rect -28577 -3372 -28530 -3308
rect -28466 -3372 -28450 -3308
rect -25378 -3339 -25274 -2961
rect -22258 -2992 -22211 -2928
rect -22147 -2992 -22131 -2928
rect -21968 2952 -16046 2961
rect -21968 -2952 -21959 2952
rect -16055 -2952 -16046 2952
rect -21968 -2961 -16046 -2952
rect -15939 2928 -15892 2992
rect -15828 2928 -15812 2992
rect -12740 2961 -12636 3339
rect -9620 3308 -9573 3372
rect -9509 3308 -9493 3372
rect -9330 9252 -3408 9261
rect -9330 3348 -9321 9252
rect -3417 3348 -3408 9252
rect -9330 3339 -3408 3348
rect -3301 9228 -3254 9292
rect -3190 9228 -3174 9292
rect -102 9261 2 9639
rect 3018 9608 3065 9672
rect 3129 9608 3145 9672
rect 3308 15552 9230 15561
rect 3308 9648 3317 15552
rect 9221 9648 9230 15552
rect 3308 9639 9230 9648
rect 9337 15528 9384 15592
rect 9448 15528 9464 15592
rect 12536 15561 12640 15939
rect 15656 15908 15703 15972
rect 15767 15908 15783 15972
rect 15946 21852 21868 21861
rect 15946 15948 15955 21852
rect 21859 15948 21868 21852
rect 15946 15939 21868 15948
rect 21975 21828 22022 21892
rect 22086 21828 22102 21892
rect 25174 21861 25278 22239
rect 28294 22208 28341 22272
rect 28405 22208 28421 22272
rect 28584 28152 34506 28161
rect 28584 22248 28593 28152
rect 34497 22248 34506 28152
rect 28584 22239 34506 22248
rect 34613 28128 34660 28192
rect 34724 28128 34740 28192
rect 37812 28161 37916 28539
rect 40932 28508 40979 28572
rect 41043 28508 41059 28572
rect 41222 34452 47144 34461
rect 41222 28548 41231 34452
rect 47135 28548 47144 34452
rect 41222 28539 47144 28548
rect 47251 34428 47298 34492
rect 47362 34428 47378 34492
rect 47251 34412 47378 34428
rect 47251 34348 47298 34412
rect 47362 34348 47378 34412
rect 47251 34332 47378 34348
rect 47251 34268 47298 34332
rect 47362 34268 47378 34332
rect 47251 34252 47378 34268
rect 47251 34188 47298 34252
rect 47362 34188 47378 34252
rect 47251 34172 47378 34188
rect 47251 34108 47298 34172
rect 47362 34108 47378 34172
rect 47251 34092 47378 34108
rect 47251 34028 47298 34092
rect 47362 34028 47378 34092
rect 47251 34012 47378 34028
rect 47251 33948 47298 34012
rect 47362 33948 47378 34012
rect 47251 33932 47378 33948
rect 47251 33868 47298 33932
rect 47362 33868 47378 33932
rect 47251 33852 47378 33868
rect 47251 33788 47298 33852
rect 47362 33788 47378 33852
rect 47251 33772 47378 33788
rect 47251 33708 47298 33772
rect 47362 33708 47378 33772
rect 47251 33692 47378 33708
rect 47251 33628 47298 33692
rect 47362 33628 47378 33692
rect 47251 33612 47378 33628
rect 47251 33548 47298 33612
rect 47362 33548 47378 33612
rect 47251 33532 47378 33548
rect 47251 33468 47298 33532
rect 47362 33468 47378 33532
rect 47251 33452 47378 33468
rect 47251 33388 47298 33452
rect 47362 33388 47378 33452
rect 47251 33372 47378 33388
rect 47251 33308 47298 33372
rect 47362 33308 47378 33372
rect 47251 33292 47378 33308
rect 47251 33228 47298 33292
rect 47362 33228 47378 33292
rect 47251 33212 47378 33228
rect 47251 33148 47298 33212
rect 47362 33148 47378 33212
rect 47251 33132 47378 33148
rect 47251 33068 47298 33132
rect 47362 33068 47378 33132
rect 47251 33052 47378 33068
rect 47251 32988 47298 33052
rect 47362 32988 47378 33052
rect 47251 32972 47378 32988
rect 47251 32908 47298 32972
rect 47362 32908 47378 32972
rect 47251 32892 47378 32908
rect 47251 32828 47298 32892
rect 47362 32828 47378 32892
rect 47251 32812 47378 32828
rect 47251 32748 47298 32812
rect 47362 32748 47378 32812
rect 47251 32732 47378 32748
rect 47251 32668 47298 32732
rect 47362 32668 47378 32732
rect 47251 32652 47378 32668
rect 47251 32588 47298 32652
rect 47362 32588 47378 32652
rect 47251 32572 47378 32588
rect 47251 32508 47298 32572
rect 47362 32508 47378 32572
rect 47251 32492 47378 32508
rect 47251 32428 47298 32492
rect 47362 32428 47378 32492
rect 47251 32412 47378 32428
rect 47251 32348 47298 32412
rect 47362 32348 47378 32412
rect 47251 32332 47378 32348
rect 47251 32268 47298 32332
rect 47362 32268 47378 32332
rect 47251 32252 47378 32268
rect 47251 32188 47298 32252
rect 47362 32188 47378 32252
rect 47251 32172 47378 32188
rect 47251 32108 47298 32172
rect 47362 32108 47378 32172
rect 47251 32092 47378 32108
rect 47251 32028 47298 32092
rect 47362 32028 47378 32092
rect 47251 32012 47378 32028
rect 47251 31948 47298 32012
rect 47362 31948 47378 32012
rect 47251 31932 47378 31948
rect 47251 31868 47298 31932
rect 47362 31868 47378 31932
rect 47251 31852 47378 31868
rect 47251 31788 47298 31852
rect 47362 31788 47378 31852
rect 47251 31772 47378 31788
rect 47251 31708 47298 31772
rect 47362 31708 47378 31772
rect 47251 31692 47378 31708
rect 47251 31628 47298 31692
rect 47362 31628 47378 31692
rect 47251 31612 47378 31628
rect 47251 31548 47298 31612
rect 47362 31548 47378 31612
rect 47251 31532 47378 31548
rect 47251 31468 47298 31532
rect 47362 31468 47378 31532
rect 47251 31452 47378 31468
rect 47251 31388 47298 31452
rect 47362 31388 47378 31452
rect 47251 31372 47378 31388
rect 47251 31308 47298 31372
rect 47362 31308 47378 31372
rect 47251 31292 47378 31308
rect 47251 31228 47298 31292
rect 47362 31228 47378 31292
rect 47251 31212 47378 31228
rect 47251 31148 47298 31212
rect 47362 31148 47378 31212
rect 47251 31132 47378 31148
rect 47251 31068 47298 31132
rect 47362 31068 47378 31132
rect 47251 31052 47378 31068
rect 47251 30988 47298 31052
rect 47362 30988 47378 31052
rect 47251 30972 47378 30988
rect 47251 30908 47298 30972
rect 47362 30908 47378 30972
rect 47251 30892 47378 30908
rect 47251 30828 47298 30892
rect 47362 30828 47378 30892
rect 47251 30812 47378 30828
rect 47251 30748 47298 30812
rect 47362 30748 47378 30812
rect 47251 30732 47378 30748
rect 47251 30668 47298 30732
rect 47362 30668 47378 30732
rect 47251 30652 47378 30668
rect 47251 30588 47298 30652
rect 47362 30588 47378 30652
rect 47251 30572 47378 30588
rect 47251 30508 47298 30572
rect 47362 30508 47378 30572
rect 47251 30492 47378 30508
rect 47251 30428 47298 30492
rect 47362 30428 47378 30492
rect 47251 30412 47378 30428
rect 47251 30348 47298 30412
rect 47362 30348 47378 30412
rect 47251 30332 47378 30348
rect 47251 30268 47298 30332
rect 47362 30268 47378 30332
rect 47251 30252 47378 30268
rect 47251 30188 47298 30252
rect 47362 30188 47378 30252
rect 47251 30172 47378 30188
rect 47251 30108 47298 30172
rect 47362 30108 47378 30172
rect 47251 30092 47378 30108
rect 47251 30028 47298 30092
rect 47362 30028 47378 30092
rect 47251 30012 47378 30028
rect 47251 29948 47298 30012
rect 47362 29948 47378 30012
rect 47251 29932 47378 29948
rect 47251 29868 47298 29932
rect 47362 29868 47378 29932
rect 47251 29852 47378 29868
rect 47251 29788 47298 29852
rect 47362 29788 47378 29852
rect 47251 29772 47378 29788
rect 47251 29708 47298 29772
rect 47362 29708 47378 29772
rect 47251 29692 47378 29708
rect 47251 29628 47298 29692
rect 47362 29628 47378 29692
rect 47251 29612 47378 29628
rect 47251 29548 47298 29612
rect 47362 29548 47378 29612
rect 47251 29532 47378 29548
rect 47251 29468 47298 29532
rect 47362 29468 47378 29532
rect 47251 29452 47378 29468
rect 47251 29388 47298 29452
rect 47362 29388 47378 29452
rect 47251 29372 47378 29388
rect 47251 29308 47298 29372
rect 47362 29308 47378 29372
rect 47251 29292 47378 29308
rect 47251 29228 47298 29292
rect 47362 29228 47378 29292
rect 47251 29212 47378 29228
rect 47251 29148 47298 29212
rect 47362 29148 47378 29212
rect 47251 29132 47378 29148
rect 47251 29068 47298 29132
rect 47362 29068 47378 29132
rect 47251 29052 47378 29068
rect 47251 28988 47298 29052
rect 47362 28988 47378 29052
rect 47251 28972 47378 28988
rect 47251 28908 47298 28972
rect 47362 28908 47378 28972
rect 47251 28892 47378 28908
rect 47251 28828 47298 28892
rect 47362 28828 47378 28892
rect 47251 28812 47378 28828
rect 47251 28748 47298 28812
rect 47362 28748 47378 28812
rect 47251 28732 47378 28748
rect 47251 28668 47298 28732
rect 47362 28668 47378 28732
rect 47251 28652 47378 28668
rect 47251 28588 47298 28652
rect 47362 28588 47378 28652
rect 47251 28572 47378 28588
rect 40932 28492 41059 28508
rect 40932 28428 40979 28492
rect 41043 28428 41059 28492
rect 40932 28412 41059 28428
rect 40932 28288 41036 28412
rect 40932 28272 41059 28288
rect 40932 28208 40979 28272
rect 41043 28208 41059 28272
rect 40932 28192 41059 28208
rect 34613 28112 34740 28128
rect 34613 28048 34660 28112
rect 34724 28048 34740 28112
rect 34613 28032 34740 28048
rect 34613 27968 34660 28032
rect 34724 27968 34740 28032
rect 34613 27952 34740 27968
rect 34613 27888 34660 27952
rect 34724 27888 34740 27952
rect 34613 27872 34740 27888
rect 34613 27808 34660 27872
rect 34724 27808 34740 27872
rect 34613 27792 34740 27808
rect 34613 27728 34660 27792
rect 34724 27728 34740 27792
rect 34613 27712 34740 27728
rect 34613 27648 34660 27712
rect 34724 27648 34740 27712
rect 34613 27632 34740 27648
rect 34613 27568 34660 27632
rect 34724 27568 34740 27632
rect 34613 27552 34740 27568
rect 34613 27488 34660 27552
rect 34724 27488 34740 27552
rect 34613 27472 34740 27488
rect 34613 27408 34660 27472
rect 34724 27408 34740 27472
rect 34613 27392 34740 27408
rect 34613 27328 34660 27392
rect 34724 27328 34740 27392
rect 34613 27312 34740 27328
rect 34613 27248 34660 27312
rect 34724 27248 34740 27312
rect 34613 27232 34740 27248
rect 34613 27168 34660 27232
rect 34724 27168 34740 27232
rect 34613 27152 34740 27168
rect 34613 27088 34660 27152
rect 34724 27088 34740 27152
rect 34613 27072 34740 27088
rect 34613 27008 34660 27072
rect 34724 27008 34740 27072
rect 34613 26992 34740 27008
rect 34613 26928 34660 26992
rect 34724 26928 34740 26992
rect 34613 26912 34740 26928
rect 34613 26848 34660 26912
rect 34724 26848 34740 26912
rect 34613 26832 34740 26848
rect 34613 26768 34660 26832
rect 34724 26768 34740 26832
rect 34613 26752 34740 26768
rect 34613 26688 34660 26752
rect 34724 26688 34740 26752
rect 34613 26672 34740 26688
rect 34613 26608 34660 26672
rect 34724 26608 34740 26672
rect 34613 26592 34740 26608
rect 34613 26528 34660 26592
rect 34724 26528 34740 26592
rect 34613 26512 34740 26528
rect 34613 26448 34660 26512
rect 34724 26448 34740 26512
rect 34613 26432 34740 26448
rect 34613 26368 34660 26432
rect 34724 26368 34740 26432
rect 34613 26352 34740 26368
rect 34613 26288 34660 26352
rect 34724 26288 34740 26352
rect 34613 26272 34740 26288
rect 34613 26208 34660 26272
rect 34724 26208 34740 26272
rect 34613 26192 34740 26208
rect 34613 26128 34660 26192
rect 34724 26128 34740 26192
rect 34613 26112 34740 26128
rect 34613 26048 34660 26112
rect 34724 26048 34740 26112
rect 34613 26032 34740 26048
rect 34613 25968 34660 26032
rect 34724 25968 34740 26032
rect 34613 25952 34740 25968
rect 34613 25888 34660 25952
rect 34724 25888 34740 25952
rect 34613 25872 34740 25888
rect 34613 25808 34660 25872
rect 34724 25808 34740 25872
rect 34613 25792 34740 25808
rect 34613 25728 34660 25792
rect 34724 25728 34740 25792
rect 34613 25712 34740 25728
rect 34613 25648 34660 25712
rect 34724 25648 34740 25712
rect 34613 25632 34740 25648
rect 34613 25568 34660 25632
rect 34724 25568 34740 25632
rect 34613 25552 34740 25568
rect 34613 25488 34660 25552
rect 34724 25488 34740 25552
rect 34613 25472 34740 25488
rect 34613 25408 34660 25472
rect 34724 25408 34740 25472
rect 34613 25392 34740 25408
rect 34613 25328 34660 25392
rect 34724 25328 34740 25392
rect 34613 25312 34740 25328
rect 34613 25248 34660 25312
rect 34724 25248 34740 25312
rect 34613 25232 34740 25248
rect 34613 25168 34660 25232
rect 34724 25168 34740 25232
rect 34613 25152 34740 25168
rect 34613 25088 34660 25152
rect 34724 25088 34740 25152
rect 34613 25072 34740 25088
rect 34613 25008 34660 25072
rect 34724 25008 34740 25072
rect 34613 24992 34740 25008
rect 34613 24928 34660 24992
rect 34724 24928 34740 24992
rect 34613 24912 34740 24928
rect 34613 24848 34660 24912
rect 34724 24848 34740 24912
rect 34613 24832 34740 24848
rect 34613 24768 34660 24832
rect 34724 24768 34740 24832
rect 34613 24752 34740 24768
rect 34613 24688 34660 24752
rect 34724 24688 34740 24752
rect 34613 24672 34740 24688
rect 34613 24608 34660 24672
rect 34724 24608 34740 24672
rect 34613 24592 34740 24608
rect 34613 24528 34660 24592
rect 34724 24528 34740 24592
rect 34613 24512 34740 24528
rect 34613 24448 34660 24512
rect 34724 24448 34740 24512
rect 34613 24432 34740 24448
rect 34613 24368 34660 24432
rect 34724 24368 34740 24432
rect 34613 24352 34740 24368
rect 34613 24288 34660 24352
rect 34724 24288 34740 24352
rect 34613 24272 34740 24288
rect 34613 24208 34660 24272
rect 34724 24208 34740 24272
rect 34613 24192 34740 24208
rect 34613 24128 34660 24192
rect 34724 24128 34740 24192
rect 34613 24112 34740 24128
rect 34613 24048 34660 24112
rect 34724 24048 34740 24112
rect 34613 24032 34740 24048
rect 34613 23968 34660 24032
rect 34724 23968 34740 24032
rect 34613 23952 34740 23968
rect 34613 23888 34660 23952
rect 34724 23888 34740 23952
rect 34613 23872 34740 23888
rect 34613 23808 34660 23872
rect 34724 23808 34740 23872
rect 34613 23792 34740 23808
rect 34613 23728 34660 23792
rect 34724 23728 34740 23792
rect 34613 23712 34740 23728
rect 34613 23648 34660 23712
rect 34724 23648 34740 23712
rect 34613 23632 34740 23648
rect 34613 23568 34660 23632
rect 34724 23568 34740 23632
rect 34613 23552 34740 23568
rect 34613 23488 34660 23552
rect 34724 23488 34740 23552
rect 34613 23472 34740 23488
rect 34613 23408 34660 23472
rect 34724 23408 34740 23472
rect 34613 23392 34740 23408
rect 34613 23328 34660 23392
rect 34724 23328 34740 23392
rect 34613 23312 34740 23328
rect 34613 23248 34660 23312
rect 34724 23248 34740 23312
rect 34613 23232 34740 23248
rect 34613 23168 34660 23232
rect 34724 23168 34740 23232
rect 34613 23152 34740 23168
rect 34613 23088 34660 23152
rect 34724 23088 34740 23152
rect 34613 23072 34740 23088
rect 34613 23008 34660 23072
rect 34724 23008 34740 23072
rect 34613 22992 34740 23008
rect 34613 22928 34660 22992
rect 34724 22928 34740 22992
rect 34613 22912 34740 22928
rect 34613 22848 34660 22912
rect 34724 22848 34740 22912
rect 34613 22832 34740 22848
rect 34613 22768 34660 22832
rect 34724 22768 34740 22832
rect 34613 22752 34740 22768
rect 34613 22688 34660 22752
rect 34724 22688 34740 22752
rect 34613 22672 34740 22688
rect 34613 22608 34660 22672
rect 34724 22608 34740 22672
rect 34613 22592 34740 22608
rect 34613 22528 34660 22592
rect 34724 22528 34740 22592
rect 34613 22512 34740 22528
rect 34613 22448 34660 22512
rect 34724 22448 34740 22512
rect 34613 22432 34740 22448
rect 34613 22368 34660 22432
rect 34724 22368 34740 22432
rect 34613 22352 34740 22368
rect 34613 22288 34660 22352
rect 34724 22288 34740 22352
rect 34613 22272 34740 22288
rect 28294 22192 28421 22208
rect 28294 22128 28341 22192
rect 28405 22128 28421 22192
rect 28294 22112 28421 22128
rect 28294 21988 28398 22112
rect 28294 21972 28421 21988
rect 28294 21908 28341 21972
rect 28405 21908 28421 21972
rect 28294 21892 28421 21908
rect 21975 21812 22102 21828
rect 21975 21748 22022 21812
rect 22086 21748 22102 21812
rect 21975 21732 22102 21748
rect 21975 21668 22022 21732
rect 22086 21668 22102 21732
rect 21975 21652 22102 21668
rect 21975 21588 22022 21652
rect 22086 21588 22102 21652
rect 21975 21572 22102 21588
rect 21975 21508 22022 21572
rect 22086 21508 22102 21572
rect 21975 21492 22102 21508
rect 21975 21428 22022 21492
rect 22086 21428 22102 21492
rect 21975 21412 22102 21428
rect 21975 21348 22022 21412
rect 22086 21348 22102 21412
rect 21975 21332 22102 21348
rect 21975 21268 22022 21332
rect 22086 21268 22102 21332
rect 21975 21252 22102 21268
rect 21975 21188 22022 21252
rect 22086 21188 22102 21252
rect 21975 21172 22102 21188
rect 21975 21108 22022 21172
rect 22086 21108 22102 21172
rect 21975 21092 22102 21108
rect 21975 21028 22022 21092
rect 22086 21028 22102 21092
rect 21975 21012 22102 21028
rect 21975 20948 22022 21012
rect 22086 20948 22102 21012
rect 21975 20932 22102 20948
rect 21975 20868 22022 20932
rect 22086 20868 22102 20932
rect 21975 20852 22102 20868
rect 21975 20788 22022 20852
rect 22086 20788 22102 20852
rect 21975 20772 22102 20788
rect 21975 20708 22022 20772
rect 22086 20708 22102 20772
rect 21975 20692 22102 20708
rect 21975 20628 22022 20692
rect 22086 20628 22102 20692
rect 21975 20612 22102 20628
rect 21975 20548 22022 20612
rect 22086 20548 22102 20612
rect 21975 20532 22102 20548
rect 21975 20468 22022 20532
rect 22086 20468 22102 20532
rect 21975 20452 22102 20468
rect 21975 20388 22022 20452
rect 22086 20388 22102 20452
rect 21975 20372 22102 20388
rect 21975 20308 22022 20372
rect 22086 20308 22102 20372
rect 21975 20292 22102 20308
rect 21975 20228 22022 20292
rect 22086 20228 22102 20292
rect 21975 20212 22102 20228
rect 21975 20148 22022 20212
rect 22086 20148 22102 20212
rect 21975 20132 22102 20148
rect 21975 20068 22022 20132
rect 22086 20068 22102 20132
rect 21975 20052 22102 20068
rect 21975 19988 22022 20052
rect 22086 19988 22102 20052
rect 21975 19972 22102 19988
rect 21975 19908 22022 19972
rect 22086 19908 22102 19972
rect 21975 19892 22102 19908
rect 21975 19828 22022 19892
rect 22086 19828 22102 19892
rect 21975 19812 22102 19828
rect 21975 19748 22022 19812
rect 22086 19748 22102 19812
rect 21975 19732 22102 19748
rect 21975 19668 22022 19732
rect 22086 19668 22102 19732
rect 21975 19652 22102 19668
rect 21975 19588 22022 19652
rect 22086 19588 22102 19652
rect 21975 19572 22102 19588
rect 21975 19508 22022 19572
rect 22086 19508 22102 19572
rect 21975 19492 22102 19508
rect 21975 19428 22022 19492
rect 22086 19428 22102 19492
rect 21975 19412 22102 19428
rect 21975 19348 22022 19412
rect 22086 19348 22102 19412
rect 21975 19332 22102 19348
rect 21975 19268 22022 19332
rect 22086 19268 22102 19332
rect 21975 19252 22102 19268
rect 21975 19188 22022 19252
rect 22086 19188 22102 19252
rect 21975 19172 22102 19188
rect 21975 19108 22022 19172
rect 22086 19108 22102 19172
rect 21975 19092 22102 19108
rect 21975 19028 22022 19092
rect 22086 19028 22102 19092
rect 21975 19012 22102 19028
rect 21975 18948 22022 19012
rect 22086 18948 22102 19012
rect 21975 18932 22102 18948
rect 21975 18868 22022 18932
rect 22086 18868 22102 18932
rect 21975 18852 22102 18868
rect 21975 18788 22022 18852
rect 22086 18788 22102 18852
rect 21975 18772 22102 18788
rect 21975 18708 22022 18772
rect 22086 18708 22102 18772
rect 21975 18692 22102 18708
rect 21975 18628 22022 18692
rect 22086 18628 22102 18692
rect 21975 18612 22102 18628
rect 21975 18548 22022 18612
rect 22086 18548 22102 18612
rect 21975 18532 22102 18548
rect 21975 18468 22022 18532
rect 22086 18468 22102 18532
rect 21975 18452 22102 18468
rect 21975 18388 22022 18452
rect 22086 18388 22102 18452
rect 21975 18372 22102 18388
rect 21975 18308 22022 18372
rect 22086 18308 22102 18372
rect 21975 18292 22102 18308
rect 21975 18228 22022 18292
rect 22086 18228 22102 18292
rect 21975 18212 22102 18228
rect 21975 18148 22022 18212
rect 22086 18148 22102 18212
rect 21975 18132 22102 18148
rect 21975 18068 22022 18132
rect 22086 18068 22102 18132
rect 21975 18052 22102 18068
rect 21975 17988 22022 18052
rect 22086 17988 22102 18052
rect 21975 17972 22102 17988
rect 21975 17908 22022 17972
rect 22086 17908 22102 17972
rect 21975 17892 22102 17908
rect 21975 17828 22022 17892
rect 22086 17828 22102 17892
rect 21975 17812 22102 17828
rect 21975 17748 22022 17812
rect 22086 17748 22102 17812
rect 21975 17732 22102 17748
rect 21975 17668 22022 17732
rect 22086 17668 22102 17732
rect 21975 17652 22102 17668
rect 21975 17588 22022 17652
rect 22086 17588 22102 17652
rect 21975 17572 22102 17588
rect 21975 17508 22022 17572
rect 22086 17508 22102 17572
rect 21975 17492 22102 17508
rect 21975 17428 22022 17492
rect 22086 17428 22102 17492
rect 21975 17412 22102 17428
rect 21975 17348 22022 17412
rect 22086 17348 22102 17412
rect 21975 17332 22102 17348
rect 21975 17268 22022 17332
rect 22086 17268 22102 17332
rect 21975 17252 22102 17268
rect 21975 17188 22022 17252
rect 22086 17188 22102 17252
rect 21975 17172 22102 17188
rect 21975 17108 22022 17172
rect 22086 17108 22102 17172
rect 21975 17092 22102 17108
rect 21975 17028 22022 17092
rect 22086 17028 22102 17092
rect 21975 17012 22102 17028
rect 21975 16948 22022 17012
rect 22086 16948 22102 17012
rect 21975 16932 22102 16948
rect 21975 16868 22022 16932
rect 22086 16868 22102 16932
rect 21975 16852 22102 16868
rect 21975 16788 22022 16852
rect 22086 16788 22102 16852
rect 21975 16772 22102 16788
rect 21975 16708 22022 16772
rect 22086 16708 22102 16772
rect 21975 16692 22102 16708
rect 21975 16628 22022 16692
rect 22086 16628 22102 16692
rect 21975 16612 22102 16628
rect 21975 16548 22022 16612
rect 22086 16548 22102 16612
rect 21975 16532 22102 16548
rect 21975 16468 22022 16532
rect 22086 16468 22102 16532
rect 21975 16452 22102 16468
rect 21975 16388 22022 16452
rect 22086 16388 22102 16452
rect 21975 16372 22102 16388
rect 21975 16308 22022 16372
rect 22086 16308 22102 16372
rect 21975 16292 22102 16308
rect 21975 16228 22022 16292
rect 22086 16228 22102 16292
rect 21975 16212 22102 16228
rect 21975 16148 22022 16212
rect 22086 16148 22102 16212
rect 21975 16132 22102 16148
rect 21975 16068 22022 16132
rect 22086 16068 22102 16132
rect 21975 16052 22102 16068
rect 21975 15988 22022 16052
rect 22086 15988 22102 16052
rect 21975 15972 22102 15988
rect 15656 15892 15783 15908
rect 15656 15828 15703 15892
rect 15767 15828 15783 15892
rect 15656 15812 15783 15828
rect 15656 15688 15760 15812
rect 15656 15672 15783 15688
rect 15656 15608 15703 15672
rect 15767 15608 15783 15672
rect 15656 15592 15783 15608
rect 9337 15512 9464 15528
rect 9337 15448 9384 15512
rect 9448 15448 9464 15512
rect 9337 15432 9464 15448
rect 9337 15368 9384 15432
rect 9448 15368 9464 15432
rect 9337 15352 9464 15368
rect 9337 15288 9384 15352
rect 9448 15288 9464 15352
rect 9337 15272 9464 15288
rect 9337 15208 9384 15272
rect 9448 15208 9464 15272
rect 9337 15192 9464 15208
rect 9337 15128 9384 15192
rect 9448 15128 9464 15192
rect 9337 15112 9464 15128
rect 9337 15048 9384 15112
rect 9448 15048 9464 15112
rect 9337 15032 9464 15048
rect 9337 14968 9384 15032
rect 9448 14968 9464 15032
rect 9337 14952 9464 14968
rect 9337 14888 9384 14952
rect 9448 14888 9464 14952
rect 9337 14872 9464 14888
rect 9337 14808 9384 14872
rect 9448 14808 9464 14872
rect 9337 14792 9464 14808
rect 9337 14728 9384 14792
rect 9448 14728 9464 14792
rect 9337 14712 9464 14728
rect 9337 14648 9384 14712
rect 9448 14648 9464 14712
rect 9337 14632 9464 14648
rect 9337 14568 9384 14632
rect 9448 14568 9464 14632
rect 9337 14552 9464 14568
rect 9337 14488 9384 14552
rect 9448 14488 9464 14552
rect 9337 14472 9464 14488
rect 9337 14408 9384 14472
rect 9448 14408 9464 14472
rect 9337 14392 9464 14408
rect 9337 14328 9384 14392
rect 9448 14328 9464 14392
rect 9337 14312 9464 14328
rect 9337 14248 9384 14312
rect 9448 14248 9464 14312
rect 9337 14232 9464 14248
rect 9337 14168 9384 14232
rect 9448 14168 9464 14232
rect 9337 14152 9464 14168
rect 9337 14088 9384 14152
rect 9448 14088 9464 14152
rect 9337 14072 9464 14088
rect 9337 14008 9384 14072
rect 9448 14008 9464 14072
rect 9337 13992 9464 14008
rect 9337 13928 9384 13992
rect 9448 13928 9464 13992
rect 9337 13912 9464 13928
rect 9337 13848 9384 13912
rect 9448 13848 9464 13912
rect 9337 13832 9464 13848
rect 9337 13768 9384 13832
rect 9448 13768 9464 13832
rect 9337 13752 9464 13768
rect 9337 13688 9384 13752
rect 9448 13688 9464 13752
rect 9337 13672 9464 13688
rect 9337 13608 9384 13672
rect 9448 13608 9464 13672
rect 9337 13592 9464 13608
rect 9337 13528 9384 13592
rect 9448 13528 9464 13592
rect 9337 13512 9464 13528
rect 9337 13448 9384 13512
rect 9448 13448 9464 13512
rect 9337 13432 9464 13448
rect 9337 13368 9384 13432
rect 9448 13368 9464 13432
rect 9337 13352 9464 13368
rect 9337 13288 9384 13352
rect 9448 13288 9464 13352
rect 9337 13272 9464 13288
rect 9337 13208 9384 13272
rect 9448 13208 9464 13272
rect 9337 13192 9464 13208
rect 9337 13128 9384 13192
rect 9448 13128 9464 13192
rect 9337 13112 9464 13128
rect 9337 13048 9384 13112
rect 9448 13048 9464 13112
rect 9337 13032 9464 13048
rect 9337 12968 9384 13032
rect 9448 12968 9464 13032
rect 9337 12952 9464 12968
rect 9337 12888 9384 12952
rect 9448 12888 9464 12952
rect 9337 12872 9464 12888
rect 9337 12808 9384 12872
rect 9448 12808 9464 12872
rect 9337 12792 9464 12808
rect 9337 12728 9384 12792
rect 9448 12728 9464 12792
rect 9337 12712 9464 12728
rect 9337 12648 9384 12712
rect 9448 12648 9464 12712
rect 9337 12632 9464 12648
rect 9337 12568 9384 12632
rect 9448 12568 9464 12632
rect 9337 12552 9464 12568
rect 9337 12488 9384 12552
rect 9448 12488 9464 12552
rect 9337 12472 9464 12488
rect 9337 12408 9384 12472
rect 9448 12408 9464 12472
rect 9337 12392 9464 12408
rect 9337 12328 9384 12392
rect 9448 12328 9464 12392
rect 9337 12312 9464 12328
rect 9337 12248 9384 12312
rect 9448 12248 9464 12312
rect 9337 12232 9464 12248
rect 9337 12168 9384 12232
rect 9448 12168 9464 12232
rect 9337 12152 9464 12168
rect 9337 12088 9384 12152
rect 9448 12088 9464 12152
rect 9337 12072 9464 12088
rect 9337 12008 9384 12072
rect 9448 12008 9464 12072
rect 9337 11992 9464 12008
rect 9337 11928 9384 11992
rect 9448 11928 9464 11992
rect 9337 11912 9464 11928
rect 9337 11848 9384 11912
rect 9448 11848 9464 11912
rect 9337 11832 9464 11848
rect 9337 11768 9384 11832
rect 9448 11768 9464 11832
rect 9337 11752 9464 11768
rect 9337 11688 9384 11752
rect 9448 11688 9464 11752
rect 9337 11672 9464 11688
rect 9337 11608 9384 11672
rect 9448 11608 9464 11672
rect 9337 11592 9464 11608
rect 9337 11528 9384 11592
rect 9448 11528 9464 11592
rect 9337 11512 9464 11528
rect 9337 11448 9384 11512
rect 9448 11448 9464 11512
rect 9337 11432 9464 11448
rect 9337 11368 9384 11432
rect 9448 11368 9464 11432
rect 9337 11352 9464 11368
rect 9337 11288 9384 11352
rect 9448 11288 9464 11352
rect 9337 11272 9464 11288
rect 9337 11208 9384 11272
rect 9448 11208 9464 11272
rect 9337 11192 9464 11208
rect 9337 11128 9384 11192
rect 9448 11128 9464 11192
rect 9337 11112 9464 11128
rect 9337 11048 9384 11112
rect 9448 11048 9464 11112
rect 9337 11032 9464 11048
rect 9337 10968 9384 11032
rect 9448 10968 9464 11032
rect 9337 10952 9464 10968
rect 9337 10888 9384 10952
rect 9448 10888 9464 10952
rect 9337 10872 9464 10888
rect 9337 10808 9384 10872
rect 9448 10808 9464 10872
rect 9337 10792 9464 10808
rect 9337 10728 9384 10792
rect 9448 10728 9464 10792
rect 9337 10712 9464 10728
rect 9337 10648 9384 10712
rect 9448 10648 9464 10712
rect 9337 10632 9464 10648
rect 9337 10568 9384 10632
rect 9448 10568 9464 10632
rect 9337 10552 9464 10568
rect 9337 10488 9384 10552
rect 9448 10488 9464 10552
rect 9337 10472 9464 10488
rect 9337 10408 9384 10472
rect 9448 10408 9464 10472
rect 9337 10392 9464 10408
rect 9337 10328 9384 10392
rect 9448 10328 9464 10392
rect 9337 10312 9464 10328
rect 9337 10248 9384 10312
rect 9448 10248 9464 10312
rect 9337 10232 9464 10248
rect 9337 10168 9384 10232
rect 9448 10168 9464 10232
rect 9337 10152 9464 10168
rect 9337 10088 9384 10152
rect 9448 10088 9464 10152
rect 9337 10072 9464 10088
rect 9337 10008 9384 10072
rect 9448 10008 9464 10072
rect 9337 9992 9464 10008
rect 9337 9928 9384 9992
rect 9448 9928 9464 9992
rect 9337 9912 9464 9928
rect 9337 9848 9384 9912
rect 9448 9848 9464 9912
rect 9337 9832 9464 9848
rect 9337 9768 9384 9832
rect 9448 9768 9464 9832
rect 9337 9752 9464 9768
rect 9337 9688 9384 9752
rect 9448 9688 9464 9752
rect 9337 9672 9464 9688
rect 3018 9592 3145 9608
rect 3018 9528 3065 9592
rect 3129 9528 3145 9592
rect 3018 9512 3145 9528
rect 3018 9388 3122 9512
rect 3018 9372 3145 9388
rect 3018 9308 3065 9372
rect 3129 9308 3145 9372
rect 3018 9292 3145 9308
rect -3301 9212 -3174 9228
rect -3301 9148 -3254 9212
rect -3190 9148 -3174 9212
rect -3301 9132 -3174 9148
rect -3301 9068 -3254 9132
rect -3190 9068 -3174 9132
rect -3301 9052 -3174 9068
rect -3301 8988 -3254 9052
rect -3190 8988 -3174 9052
rect -3301 8972 -3174 8988
rect -3301 8908 -3254 8972
rect -3190 8908 -3174 8972
rect -3301 8892 -3174 8908
rect -3301 8828 -3254 8892
rect -3190 8828 -3174 8892
rect -3301 8812 -3174 8828
rect -3301 8748 -3254 8812
rect -3190 8748 -3174 8812
rect -3301 8732 -3174 8748
rect -3301 8668 -3254 8732
rect -3190 8668 -3174 8732
rect -3301 8652 -3174 8668
rect -3301 8588 -3254 8652
rect -3190 8588 -3174 8652
rect -3301 8572 -3174 8588
rect -3301 8508 -3254 8572
rect -3190 8508 -3174 8572
rect -3301 8492 -3174 8508
rect -3301 8428 -3254 8492
rect -3190 8428 -3174 8492
rect -3301 8412 -3174 8428
rect -3301 8348 -3254 8412
rect -3190 8348 -3174 8412
rect -3301 8332 -3174 8348
rect -3301 8268 -3254 8332
rect -3190 8268 -3174 8332
rect -3301 8252 -3174 8268
rect -3301 8188 -3254 8252
rect -3190 8188 -3174 8252
rect -3301 8172 -3174 8188
rect -3301 8108 -3254 8172
rect -3190 8108 -3174 8172
rect -3301 8092 -3174 8108
rect -3301 8028 -3254 8092
rect -3190 8028 -3174 8092
rect -3301 8012 -3174 8028
rect -3301 7948 -3254 8012
rect -3190 7948 -3174 8012
rect -3301 7932 -3174 7948
rect -3301 7868 -3254 7932
rect -3190 7868 -3174 7932
rect -3301 7852 -3174 7868
rect -3301 7788 -3254 7852
rect -3190 7788 -3174 7852
rect -3301 7772 -3174 7788
rect -3301 7708 -3254 7772
rect -3190 7708 -3174 7772
rect -3301 7692 -3174 7708
rect -3301 7628 -3254 7692
rect -3190 7628 -3174 7692
rect -3301 7612 -3174 7628
rect -3301 7548 -3254 7612
rect -3190 7548 -3174 7612
rect -3301 7532 -3174 7548
rect -3301 7468 -3254 7532
rect -3190 7468 -3174 7532
rect -3301 7452 -3174 7468
rect -3301 7388 -3254 7452
rect -3190 7388 -3174 7452
rect -3301 7372 -3174 7388
rect -3301 7308 -3254 7372
rect -3190 7308 -3174 7372
rect -3301 7292 -3174 7308
rect -3301 7228 -3254 7292
rect -3190 7228 -3174 7292
rect -3301 7212 -3174 7228
rect -3301 7148 -3254 7212
rect -3190 7148 -3174 7212
rect -3301 7132 -3174 7148
rect -3301 7068 -3254 7132
rect -3190 7068 -3174 7132
rect -3301 7052 -3174 7068
rect -3301 6988 -3254 7052
rect -3190 6988 -3174 7052
rect -3301 6972 -3174 6988
rect -3301 6908 -3254 6972
rect -3190 6908 -3174 6972
rect -3301 6892 -3174 6908
rect -3301 6828 -3254 6892
rect -3190 6828 -3174 6892
rect -3301 6812 -3174 6828
rect -3301 6748 -3254 6812
rect -3190 6748 -3174 6812
rect -3301 6732 -3174 6748
rect -3301 6668 -3254 6732
rect -3190 6668 -3174 6732
rect -3301 6652 -3174 6668
rect -3301 6588 -3254 6652
rect -3190 6588 -3174 6652
rect -3301 6572 -3174 6588
rect -3301 6508 -3254 6572
rect -3190 6508 -3174 6572
rect -3301 6492 -3174 6508
rect -3301 6428 -3254 6492
rect -3190 6428 -3174 6492
rect -3301 6412 -3174 6428
rect -3301 6348 -3254 6412
rect -3190 6348 -3174 6412
rect -3301 6332 -3174 6348
rect -3301 6268 -3254 6332
rect -3190 6268 -3174 6332
rect -3301 6252 -3174 6268
rect -3301 6188 -3254 6252
rect -3190 6188 -3174 6252
rect -3301 6172 -3174 6188
rect -3301 6108 -3254 6172
rect -3190 6108 -3174 6172
rect -3301 6092 -3174 6108
rect -3301 6028 -3254 6092
rect -3190 6028 -3174 6092
rect -3301 6012 -3174 6028
rect -3301 5948 -3254 6012
rect -3190 5948 -3174 6012
rect -3301 5932 -3174 5948
rect -3301 5868 -3254 5932
rect -3190 5868 -3174 5932
rect -3301 5852 -3174 5868
rect -3301 5788 -3254 5852
rect -3190 5788 -3174 5852
rect -3301 5772 -3174 5788
rect -3301 5708 -3254 5772
rect -3190 5708 -3174 5772
rect -3301 5692 -3174 5708
rect -3301 5628 -3254 5692
rect -3190 5628 -3174 5692
rect -3301 5612 -3174 5628
rect -3301 5548 -3254 5612
rect -3190 5548 -3174 5612
rect -3301 5532 -3174 5548
rect -3301 5468 -3254 5532
rect -3190 5468 -3174 5532
rect -3301 5452 -3174 5468
rect -3301 5388 -3254 5452
rect -3190 5388 -3174 5452
rect -3301 5372 -3174 5388
rect -3301 5308 -3254 5372
rect -3190 5308 -3174 5372
rect -3301 5292 -3174 5308
rect -3301 5228 -3254 5292
rect -3190 5228 -3174 5292
rect -3301 5212 -3174 5228
rect -3301 5148 -3254 5212
rect -3190 5148 -3174 5212
rect -3301 5132 -3174 5148
rect -3301 5068 -3254 5132
rect -3190 5068 -3174 5132
rect -3301 5052 -3174 5068
rect -3301 4988 -3254 5052
rect -3190 4988 -3174 5052
rect -3301 4972 -3174 4988
rect -3301 4908 -3254 4972
rect -3190 4908 -3174 4972
rect -3301 4892 -3174 4908
rect -3301 4828 -3254 4892
rect -3190 4828 -3174 4892
rect -3301 4812 -3174 4828
rect -3301 4748 -3254 4812
rect -3190 4748 -3174 4812
rect -3301 4732 -3174 4748
rect -3301 4668 -3254 4732
rect -3190 4668 -3174 4732
rect -3301 4652 -3174 4668
rect -3301 4588 -3254 4652
rect -3190 4588 -3174 4652
rect -3301 4572 -3174 4588
rect -3301 4508 -3254 4572
rect -3190 4508 -3174 4572
rect -3301 4492 -3174 4508
rect -3301 4428 -3254 4492
rect -3190 4428 -3174 4492
rect -3301 4412 -3174 4428
rect -3301 4348 -3254 4412
rect -3190 4348 -3174 4412
rect -3301 4332 -3174 4348
rect -3301 4268 -3254 4332
rect -3190 4268 -3174 4332
rect -3301 4252 -3174 4268
rect -3301 4188 -3254 4252
rect -3190 4188 -3174 4252
rect -3301 4172 -3174 4188
rect -3301 4108 -3254 4172
rect -3190 4108 -3174 4172
rect -3301 4092 -3174 4108
rect -3301 4028 -3254 4092
rect -3190 4028 -3174 4092
rect -3301 4012 -3174 4028
rect -3301 3948 -3254 4012
rect -3190 3948 -3174 4012
rect -3301 3932 -3174 3948
rect -3301 3868 -3254 3932
rect -3190 3868 -3174 3932
rect -3301 3852 -3174 3868
rect -3301 3788 -3254 3852
rect -3190 3788 -3174 3852
rect -3301 3772 -3174 3788
rect -3301 3708 -3254 3772
rect -3190 3708 -3174 3772
rect -3301 3692 -3174 3708
rect -3301 3628 -3254 3692
rect -3190 3628 -3174 3692
rect -3301 3612 -3174 3628
rect -3301 3548 -3254 3612
rect -3190 3548 -3174 3612
rect -3301 3532 -3174 3548
rect -3301 3468 -3254 3532
rect -3190 3468 -3174 3532
rect -3301 3452 -3174 3468
rect -3301 3388 -3254 3452
rect -3190 3388 -3174 3452
rect -3301 3372 -3174 3388
rect -9620 3292 -9493 3308
rect -9620 3228 -9573 3292
rect -9509 3228 -9493 3292
rect -9620 3212 -9493 3228
rect -9620 3088 -9516 3212
rect -9620 3072 -9493 3088
rect -9620 3008 -9573 3072
rect -9509 3008 -9493 3072
rect -9620 2992 -9493 3008
rect -15939 2912 -15812 2928
rect -15939 2848 -15892 2912
rect -15828 2848 -15812 2912
rect -15939 2832 -15812 2848
rect -15939 2768 -15892 2832
rect -15828 2768 -15812 2832
rect -15939 2752 -15812 2768
rect -15939 2688 -15892 2752
rect -15828 2688 -15812 2752
rect -15939 2672 -15812 2688
rect -15939 2608 -15892 2672
rect -15828 2608 -15812 2672
rect -15939 2592 -15812 2608
rect -15939 2528 -15892 2592
rect -15828 2528 -15812 2592
rect -15939 2512 -15812 2528
rect -15939 2448 -15892 2512
rect -15828 2448 -15812 2512
rect -15939 2432 -15812 2448
rect -15939 2368 -15892 2432
rect -15828 2368 -15812 2432
rect -15939 2352 -15812 2368
rect -15939 2288 -15892 2352
rect -15828 2288 -15812 2352
rect -15939 2272 -15812 2288
rect -15939 2208 -15892 2272
rect -15828 2208 -15812 2272
rect -15939 2192 -15812 2208
rect -15939 2128 -15892 2192
rect -15828 2128 -15812 2192
rect -15939 2112 -15812 2128
rect -15939 2048 -15892 2112
rect -15828 2048 -15812 2112
rect -15939 2032 -15812 2048
rect -15939 1968 -15892 2032
rect -15828 1968 -15812 2032
rect -15939 1952 -15812 1968
rect -15939 1888 -15892 1952
rect -15828 1888 -15812 1952
rect -15939 1872 -15812 1888
rect -15939 1808 -15892 1872
rect -15828 1808 -15812 1872
rect -15939 1792 -15812 1808
rect -15939 1728 -15892 1792
rect -15828 1728 -15812 1792
rect -15939 1712 -15812 1728
rect -15939 1648 -15892 1712
rect -15828 1648 -15812 1712
rect -15939 1632 -15812 1648
rect -15939 1568 -15892 1632
rect -15828 1568 -15812 1632
rect -15939 1552 -15812 1568
rect -15939 1488 -15892 1552
rect -15828 1488 -15812 1552
rect -15939 1472 -15812 1488
rect -15939 1408 -15892 1472
rect -15828 1408 -15812 1472
rect -15939 1392 -15812 1408
rect -15939 1328 -15892 1392
rect -15828 1328 -15812 1392
rect -15939 1312 -15812 1328
rect -15939 1248 -15892 1312
rect -15828 1248 -15812 1312
rect -15939 1232 -15812 1248
rect -15939 1168 -15892 1232
rect -15828 1168 -15812 1232
rect -15939 1152 -15812 1168
rect -15939 1088 -15892 1152
rect -15828 1088 -15812 1152
rect -15939 1072 -15812 1088
rect -15939 1008 -15892 1072
rect -15828 1008 -15812 1072
rect -15939 992 -15812 1008
rect -15939 928 -15892 992
rect -15828 928 -15812 992
rect -15939 912 -15812 928
rect -15939 848 -15892 912
rect -15828 848 -15812 912
rect -15939 832 -15812 848
rect -15939 768 -15892 832
rect -15828 768 -15812 832
rect -15939 752 -15812 768
rect -15939 688 -15892 752
rect -15828 688 -15812 752
rect -15939 672 -15812 688
rect -15939 608 -15892 672
rect -15828 608 -15812 672
rect -15939 592 -15812 608
rect -15939 528 -15892 592
rect -15828 528 -15812 592
rect -15939 512 -15812 528
rect -15939 448 -15892 512
rect -15828 448 -15812 512
rect -15939 432 -15812 448
rect -15939 368 -15892 432
rect -15828 368 -15812 432
rect -15939 352 -15812 368
rect -15939 288 -15892 352
rect -15828 288 -15812 352
rect -15939 272 -15812 288
rect -15939 208 -15892 272
rect -15828 208 -15812 272
rect -15939 192 -15812 208
rect -15939 128 -15892 192
rect -15828 128 -15812 192
rect -15939 112 -15812 128
rect -15939 48 -15892 112
rect -15828 48 -15812 112
rect -15939 32 -15812 48
rect -15939 -32 -15892 32
rect -15828 -32 -15812 32
rect -15939 -48 -15812 -32
rect -15939 -112 -15892 -48
rect -15828 -112 -15812 -48
rect -15939 -128 -15812 -112
rect -15939 -192 -15892 -128
rect -15828 -192 -15812 -128
rect -15939 -208 -15812 -192
rect -15939 -272 -15892 -208
rect -15828 -272 -15812 -208
rect -15939 -288 -15812 -272
rect -15939 -352 -15892 -288
rect -15828 -352 -15812 -288
rect -15939 -368 -15812 -352
rect -15939 -432 -15892 -368
rect -15828 -432 -15812 -368
rect -15939 -448 -15812 -432
rect -15939 -512 -15892 -448
rect -15828 -512 -15812 -448
rect -15939 -528 -15812 -512
rect -15939 -592 -15892 -528
rect -15828 -592 -15812 -528
rect -15939 -608 -15812 -592
rect -15939 -672 -15892 -608
rect -15828 -672 -15812 -608
rect -15939 -688 -15812 -672
rect -15939 -752 -15892 -688
rect -15828 -752 -15812 -688
rect -15939 -768 -15812 -752
rect -15939 -832 -15892 -768
rect -15828 -832 -15812 -768
rect -15939 -848 -15812 -832
rect -15939 -912 -15892 -848
rect -15828 -912 -15812 -848
rect -15939 -928 -15812 -912
rect -15939 -992 -15892 -928
rect -15828 -992 -15812 -928
rect -15939 -1008 -15812 -992
rect -15939 -1072 -15892 -1008
rect -15828 -1072 -15812 -1008
rect -15939 -1088 -15812 -1072
rect -15939 -1152 -15892 -1088
rect -15828 -1152 -15812 -1088
rect -15939 -1168 -15812 -1152
rect -15939 -1232 -15892 -1168
rect -15828 -1232 -15812 -1168
rect -15939 -1248 -15812 -1232
rect -15939 -1312 -15892 -1248
rect -15828 -1312 -15812 -1248
rect -15939 -1328 -15812 -1312
rect -15939 -1392 -15892 -1328
rect -15828 -1392 -15812 -1328
rect -15939 -1408 -15812 -1392
rect -15939 -1472 -15892 -1408
rect -15828 -1472 -15812 -1408
rect -15939 -1488 -15812 -1472
rect -15939 -1552 -15892 -1488
rect -15828 -1552 -15812 -1488
rect -15939 -1568 -15812 -1552
rect -15939 -1632 -15892 -1568
rect -15828 -1632 -15812 -1568
rect -15939 -1648 -15812 -1632
rect -15939 -1712 -15892 -1648
rect -15828 -1712 -15812 -1648
rect -15939 -1728 -15812 -1712
rect -15939 -1792 -15892 -1728
rect -15828 -1792 -15812 -1728
rect -15939 -1808 -15812 -1792
rect -15939 -1872 -15892 -1808
rect -15828 -1872 -15812 -1808
rect -15939 -1888 -15812 -1872
rect -15939 -1952 -15892 -1888
rect -15828 -1952 -15812 -1888
rect -15939 -1968 -15812 -1952
rect -15939 -2032 -15892 -1968
rect -15828 -2032 -15812 -1968
rect -15939 -2048 -15812 -2032
rect -15939 -2112 -15892 -2048
rect -15828 -2112 -15812 -2048
rect -15939 -2128 -15812 -2112
rect -15939 -2192 -15892 -2128
rect -15828 -2192 -15812 -2128
rect -15939 -2208 -15812 -2192
rect -15939 -2272 -15892 -2208
rect -15828 -2272 -15812 -2208
rect -15939 -2288 -15812 -2272
rect -15939 -2352 -15892 -2288
rect -15828 -2352 -15812 -2288
rect -15939 -2368 -15812 -2352
rect -15939 -2432 -15892 -2368
rect -15828 -2432 -15812 -2368
rect -15939 -2448 -15812 -2432
rect -15939 -2512 -15892 -2448
rect -15828 -2512 -15812 -2448
rect -15939 -2528 -15812 -2512
rect -15939 -2592 -15892 -2528
rect -15828 -2592 -15812 -2528
rect -15939 -2608 -15812 -2592
rect -15939 -2672 -15892 -2608
rect -15828 -2672 -15812 -2608
rect -15939 -2688 -15812 -2672
rect -15939 -2752 -15892 -2688
rect -15828 -2752 -15812 -2688
rect -15939 -2768 -15812 -2752
rect -15939 -2832 -15892 -2768
rect -15828 -2832 -15812 -2768
rect -15939 -2848 -15812 -2832
rect -15939 -2912 -15892 -2848
rect -15828 -2912 -15812 -2848
rect -15939 -2928 -15812 -2912
rect -22258 -3008 -22131 -2992
rect -22258 -3072 -22211 -3008
rect -22147 -3072 -22131 -3008
rect -22258 -3088 -22131 -3072
rect -22258 -3212 -22154 -3088
rect -22258 -3228 -22131 -3212
rect -22258 -3292 -22211 -3228
rect -22147 -3292 -22131 -3228
rect -22258 -3308 -22131 -3292
rect -28577 -3388 -28450 -3372
rect -28577 -3452 -28530 -3388
rect -28466 -3452 -28450 -3388
rect -28577 -3468 -28450 -3452
rect -28577 -3532 -28530 -3468
rect -28466 -3532 -28450 -3468
rect -28577 -3548 -28450 -3532
rect -28577 -3612 -28530 -3548
rect -28466 -3612 -28450 -3548
rect -28577 -3628 -28450 -3612
rect -28577 -3692 -28530 -3628
rect -28466 -3692 -28450 -3628
rect -28577 -3708 -28450 -3692
rect -28577 -3772 -28530 -3708
rect -28466 -3772 -28450 -3708
rect -28577 -3788 -28450 -3772
rect -28577 -3852 -28530 -3788
rect -28466 -3852 -28450 -3788
rect -28577 -3868 -28450 -3852
rect -28577 -3932 -28530 -3868
rect -28466 -3932 -28450 -3868
rect -28577 -3948 -28450 -3932
rect -28577 -4012 -28530 -3948
rect -28466 -4012 -28450 -3948
rect -28577 -4028 -28450 -4012
rect -28577 -4092 -28530 -4028
rect -28466 -4092 -28450 -4028
rect -28577 -4108 -28450 -4092
rect -28577 -4172 -28530 -4108
rect -28466 -4172 -28450 -4108
rect -28577 -4188 -28450 -4172
rect -28577 -4252 -28530 -4188
rect -28466 -4252 -28450 -4188
rect -28577 -4268 -28450 -4252
rect -28577 -4332 -28530 -4268
rect -28466 -4332 -28450 -4268
rect -28577 -4348 -28450 -4332
rect -28577 -4412 -28530 -4348
rect -28466 -4412 -28450 -4348
rect -28577 -4428 -28450 -4412
rect -28577 -4492 -28530 -4428
rect -28466 -4492 -28450 -4428
rect -28577 -4508 -28450 -4492
rect -28577 -4572 -28530 -4508
rect -28466 -4572 -28450 -4508
rect -28577 -4588 -28450 -4572
rect -28577 -4652 -28530 -4588
rect -28466 -4652 -28450 -4588
rect -28577 -4668 -28450 -4652
rect -28577 -4732 -28530 -4668
rect -28466 -4732 -28450 -4668
rect -28577 -4748 -28450 -4732
rect -28577 -4812 -28530 -4748
rect -28466 -4812 -28450 -4748
rect -28577 -4828 -28450 -4812
rect -28577 -4892 -28530 -4828
rect -28466 -4892 -28450 -4828
rect -28577 -4908 -28450 -4892
rect -28577 -4972 -28530 -4908
rect -28466 -4972 -28450 -4908
rect -28577 -4988 -28450 -4972
rect -28577 -5052 -28530 -4988
rect -28466 -5052 -28450 -4988
rect -28577 -5068 -28450 -5052
rect -28577 -5132 -28530 -5068
rect -28466 -5132 -28450 -5068
rect -28577 -5148 -28450 -5132
rect -28577 -5212 -28530 -5148
rect -28466 -5212 -28450 -5148
rect -28577 -5228 -28450 -5212
rect -28577 -5292 -28530 -5228
rect -28466 -5292 -28450 -5228
rect -28577 -5308 -28450 -5292
rect -28577 -5372 -28530 -5308
rect -28466 -5372 -28450 -5308
rect -28577 -5388 -28450 -5372
rect -28577 -5452 -28530 -5388
rect -28466 -5452 -28450 -5388
rect -28577 -5468 -28450 -5452
rect -28577 -5532 -28530 -5468
rect -28466 -5532 -28450 -5468
rect -28577 -5548 -28450 -5532
rect -28577 -5612 -28530 -5548
rect -28466 -5612 -28450 -5548
rect -28577 -5628 -28450 -5612
rect -28577 -5692 -28530 -5628
rect -28466 -5692 -28450 -5628
rect -28577 -5708 -28450 -5692
rect -28577 -5772 -28530 -5708
rect -28466 -5772 -28450 -5708
rect -28577 -5788 -28450 -5772
rect -28577 -5852 -28530 -5788
rect -28466 -5852 -28450 -5788
rect -28577 -5868 -28450 -5852
rect -28577 -5932 -28530 -5868
rect -28466 -5932 -28450 -5868
rect -28577 -5948 -28450 -5932
rect -28577 -6012 -28530 -5948
rect -28466 -6012 -28450 -5948
rect -28577 -6028 -28450 -6012
rect -28577 -6092 -28530 -6028
rect -28466 -6092 -28450 -6028
rect -28577 -6108 -28450 -6092
rect -28577 -6172 -28530 -6108
rect -28466 -6172 -28450 -6108
rect -28577 -6188 -28450 -6172
rect -28577 -6252 -28530 -6188
rect -28466 -6252 -28450 -6188
rect -28577 -6268 -28450 -6252
rect -28577 -6332 -28530 -6268
rect -28466 -6332 -28450 -6268
rect -28577 -6348 -28450 -6332
rect -28577 -6412 -28530 -6348
rect -28466 -6412 -28450 -6348
rect -28577 -6428 -28450 -6412
rect -28577 -6492 -28530 -6428
rect -28466 -6492 -28450 -6428
rect -28577 -6508 -28450 -6492
rect -28577 -6572 -28530 -6508
rect -28466 -6572 -28450 -6508
rect -28577 -6588 -28450 -6572
rect -28577 -6652 -28530 -6588
rect -28466 -6652 -28450 -6588
rect -28577 -6668 -28450 -6652
rect -28577 -6732 -28530 -6668
rect -28466 -6732 -28450 -6668
rect -28577 -6748 -28450 -6732
rect -28577 -6812 -28530 -6748
rect -28466 -6812 -28450 -6748
rect -28577 -6828 -28450 -6812
rect -28577 -6892 -28530 -6828
rect -28466 -6892 -28450 -6828
rect -28577 -6908 -28450 -6892
rect -28577 -6972 -28530 -6908
rect -28466 -6972 -28450 -6908
rect -28577 -6988 -28450 -6972
rect -28577 -7052 -28530 -6988
rect -28466 -7052 -28450 -6988
rect -28577 -7068 -28450 -7052
rect -28577 -7132 -28530 -7068
rect -28466 -7132 -28450 -7068
rect -28577 -7148 -28450 -7132
rect -28577 -7212 -28530 -7148
rect -28466 -7212 -28450 -7148
rect -28577 -7228 -28450 -7212
rect -28577 -7292 -28530 -7228
rect -28466 -7292 -28450 -7228
rect -28577 -7308 -28450 -7292
rect -28577 -7372 -28530 -7308
rect -28466 -7372 -28450 -7308
rect -28577 -7388 -28450 -7372
rect -28577 -7452 -28530 -7388
rect -28466 -7452 -28450 -7388
rect -28577 -7468 -28450 -7452
rect -28577 -7532 -28530 -7468
rect -28466 -7532 -28450 -7468
rect -28577 -7548 -28450 -7532
rect -28577 -7612 -28530 -7548
rect -28466 -7612 -28450 -7548
rect -28577 -7628 -28450 -7612
rect -28577 -7692 -28530 -7628
rect -28466 -7692 -28450 -7628
rect -28577 -7708 -28450 -7692
rect -28577 -7772 -28530 -7708
rect -28466 -7772 -28450 -7708
rect -28577 -7788 -28450 -7772
rect -28577 -7852 -28530 -7788
rect -28466 -7852 -28450 -7788
rect -28577 -7868 -28450 -7852
rect -28577 -7932 -28530 -7868
rect -28466 -7932 -28450 -7868
rect -28577 -7948 -28450 -7932
rect -28577 -8012 -28530 -7948
rect -28466 -8012 -28450 -7948
rect -28577 -8028 -28450 -8012
rect -28577 -8092 -28530 -8028
rect -28466 -8092 -28450 -8028
rect -28577 -8108 -28450 -8092
rect -28577 -8172 -28530 -8108
rect -28466 -8172 -28450 -8108
rect -28577 -8188 -28450 -8172
rect -28577 -8252 -28530 -8188
rect -28466 -8252 -28450 -8188
rect -28577 -8268 -28450 -8252
rect -28577 -8332 -28530 -8268
rect -28466 -8332 -28450 -8268
rect -28577 -8348 -28450 -8332
rect -28577 -8412 -28530 -8348
rect -28466 -8412 -28450 -8348
rect -28577 -8428 -28450 -8412
rect -28577 -8492 -28530 -8428
rect -28466 -8492 -28450 -8428
rect -28577 -8508 -28450 -8492
rect -28577 -8572 -28530 -8508
rect -28466 -8572 -28450 -8508
rect -28577 -8588 -28450 -8572
rect -28577 -8652 -28530 -8588
rect -28466 -8652 -28450 -8588
rect -28577 -8668 -28450 -8652
rect -28577 -8732 -28530 -8668
rect -28466 -8732 -28450 -8668
rect -28577 -8748 -28450 -8732
rect -28577 -8812 -28530 -8748
rect -28466 -8812 -28450 -8748
rect -28577 -8828 -28450 -8812
rect -28577 -8892 -28530 -8828
rect -28466 -8892 -28450 -8828
rect -28577 -8908 -28450 -8892
rect -28577 -8972 -28530 -8908
rect -28466 -8972 -28450 -8908
rect -28577 -8988 -28450 -8972
rect -28577 -9052 -28530 -8988
rect -28466 -9052 -28450 -8988
rect -28577 -9068 -28450 -9052
rect -28577 -9132 -28530 -9068
rect -28466 -9132 -28450 -9068
rect -28577 -9148 -28450 -9132
rect -28577 -9212 -28530 -9148
rect -28466 -9212 -28450 -9148
rect -28577 -9228 -28450 -9212
rect -34896 -9308 -34769 -9292
rect -34896 -9372 -34849 -9308
rect -34785 -9372 -34769 -9308
rect -34896 -9388 -34769 -9372
rect -34896 -9512 -34792 -9388
rect -34896 -9528 -34769 -9512
rect -34896 -9592 -34849 -9528
rect -34785 -9592 -34769 -9528
rect -34896 -9608 -34769 -9592
rect -41215 -9688 -41088 -9672
rect -41215 -9752 -41168 -9688
rect -41104 -9752 -41088 -9688
rect -41215 -9768 -41088 -9752
rect -41215 -9832 -41168 -9768
rect -41104 -9832 -41088 -9768
rect -41215 -9848 -41088 -9832
rect -41215 -9912 -41168 -9848
rect -41104 -9912 -41088 -9848
rect -41215 -9928 -41088 -9912
rect -41215 -9992 -41168 -9928
rect -41104 -9992 -41088 -9928
rect -41215 -10008 -41088 -9992
rect -41215 -10072 -41168 -10008
rect -41104 -10072 -41088 -10008
rect -41215 -10088 -41088 -10072
rect -41215 -10152 -41168 -10088
rect -41104 -10152 -41088 -10088
rect -41215 -10168 -41088 -10152
rect -41215 -10232 -41168 -10168
rect -41104 -10232 -41088 -10168
rect -41215 -10248 -41088 -10232
rect -41215 -10312 -41168 -10248
rect -41104 -10312 -41088 -10248
rect -41215 -10328 -41088 -10312
rect -41215 -10392 -41168 -10328
rect -41104 -10392 -41088 -10328
rect -41215 -10408 -41088 -10392
rect -41215 -10472 -41168 -10408
rect -41104 -10472 -41088 -10408
rect -41215 -10488 -41088 -10472
rect -41215 -10552 -41168 -10488
rect -41104 -10552 -41088 -10488
rect -41215 -10568 -41088 -10552
rect -41215 -10632 -41168 -10568
rect -41104 -10632 -41088 -10568
rect -41215 -10648 -41088 -10632
rect -41215 -10712 -41168 -10648
rect -41104 -10712 -41088 -10648
rect -41215 -10728 -41088 -10712
rect -41215 -10792 -41168 -10728
rect -41104 -10792 -41088 -10728
rect -41215 -10808 -41088 -10792
rect -41215 -10872 -41168 -10808
rect -41104 -10872 -41088 -10808
rect -41215 -10888 -41088 -10872
rect -41215 -10952 -41168 -10888
rect -41104 -10952 -41088 -10888
rect -41215 -10968 -41088 -10952
rect -41215 -11032 -41168 -10968
rect -41104 -11032 -41088 -10968
rect -41215 -11048 -41088 -11032
rect -41215 -11112 -41168 -11048
rect -41104 -11112 -41088 -11048
rect -41215 -11128 -41088 -11112
rect -41215 -11192 -41168 -11128
rect -41104 -11192 -41088 -11128
rect -41215 -11208 -41088 -11192
rect -41215 -11272 -41168 -11208
rect -41104 -11272 -41088 -11208
rect -41215 -11288 -41088 -11272
rect -41215 -11352 -41168 -11288
rect -41104 -11352 -41088 -11288
rect -41215 -11368 -41088 -11352
rect -41215 -11432 -41168 -11368
rect -41104 -11432 -41088 -11368
rect -41215 -11448 -41088 -11432
rect -41215 -11512 -41168 -11448
rect -41104 -11512 -41088 -11448
rect -41215 -11528 -41088 -11512
rect -41215 -11592 -41168 -11528
rect -41104 -11592 -41088 -11528
rect -41215 -11608 -41088 -11592
rect -41215 -11672 -41168 -11608
rect -41104 -11672 -41088 -11608
rect -41215 -11688 -41088 -11672
rect -41215 -11752 -41168 -11688
rect -41104 -11752 -41088 -11688
rect -41215 -11768 -41088 -11752
rect -41215 -11832 -41168 -11768
rect -41104 -11832 -41088 -11768
rect -41215 -11848 -41088 -11832
rect -41215 -11912 -41168 -11848
rect -41104 -11912 -41088 -11848
rect -41215 -11928 -41088 -11912
rect -41215 -11992 -41168 -11928
rect -41104 -11992 -41088 -11928
rect -41215 -12008 -41088 -11992
rect -41215 -12072 -41168 -12008
rect -41104 -12072 -41088 -12008
rect -41215 -12088 -41088 -12072
rect -41215 -12152 -41168 -12088
rect -41104 -12152 -41088 -12088
rect -41215 -12168 -41088 -12152
rect -41215 -12232 -41168 -12168
rect -41104 -12232 -41088 -12168
rect -41215 -12248 -41088 -12232
rect -41215 -12312 -41168 -12248
rect -41104 -12312 -41088 -12248
rect -41215 -12328 -41088 -12312
rect -41215 -12392 -41168 -12328
rect -41104 -12392 -41088 -12328
rect -41215 -12408 -41088 -12392
rect -41215 -12472 -41168 -12408
rect -41104 -12472 -41088 -12408
rect -41215 -12488 -41088 -12472
rect -41215 -12552 -41168 -12488
rect -41104 -12552 -41088 -12488
rect -41215 -12568 -41088 -12552
rect -41215 -12632 -41168 -12568
rect -41104 -12632 -41088 -12568
rect -41215 -12648 -41088 -12632
rect -41215 -12712 -41168 -12648
rect -41104 -12712 -41088 -12648
rect -41215 -12728 -41088 -12712
rect -41215 -12792 -41168 -12728
rect -41104 -12792 -41088 -12728
rect -41215 -12808 -41088 -12792
rect -41215 -12872 -41168 -12808
rect -41104 -12872 -41088 -12808
rect -41215 -12888 -41088 -12872
rect -41215 -12952 -41168 -12888
rect -41104 -12952 -41088 -12888
rect -41215 -12968 -41088 -12952
rect -41215 -13032 -41168 -12968
rect -41104 -13032 -41088 -12968
rect -41215 -13048 -41088 -13032
rect -41215 -13112 -41168 -13048
rect -41104 -13112 -41088 -13048
rect -41215 -13128 -41088 -13112
rect -41215 -13192 -41168 -13128
rect -41104 -13192 -41088 -13128
rect -41215 -13208 -41088 -13192
rect -41215 -13272 -41168 -13208
rect -41104 -13272 -41088 -13208
rect -41215 -13288 -41088 -13272
rect -41215 -13352 -41168 -13288
rect -41104 -13352 -41088 -13288
rect -41215 -13368 -41088 -13352
rect -41215 -13432 -41168 -13368
rect -41104 -13432 -41088 -13368
rect -41215 -13448 -41088 -13432
rect -41215 -13512 -41168 -13448
rect -41104 -13512 -41088 -13448
rect -41215 -13528 -41088 -13512
rect -41215 -13592 -41168 -13528
rect -41104 -13592 -41088 -13528
rect -41215 -13608 -41088 -13592
rect -41215 -13672 -41168 -13608
rect -41104 -13672 -41088 -13608
rect -41215 -13688 -41088 -13672
rect -41215 -13752 -41168 -13688
rect -41104 -13752 -41088 -13688
rect -41215 -13768 -41088 -13752
rect -41215 -13832 -41168 -13768
rect -41104 -13832 -41088 -13768
rect -41215 -13848 -41088 -13832
rect -41215 -13912 -41168 -13848
rect -41104 -13912 -41088 -13848
rect -41215 -13928 -41088 -13912
rect -41215 -13992 -41168 -13928
rect -41104 -13992 -41088 -13928
rect -41215 -14008 -41088 -13992
rect -41215 -14072 -41168 -14008
rect -41104 -14072 -41088 -14008
rect -41215 -14088 -41088 -14072
rect -41215 -14152 -41168 -14088
rect -41104 -14152 -41088 -14088
rect -41215 -14168 -41088 -14152
rect -41215 -14232 -41168 -14168
rect -41104 -14232 -41088 -14168
rect -41215 -14248 -41088 -14232
rect -41215 -14312 -41168 -14248
rect -41104 -14312 -41088 -14248
rect -41215 -14328 -41088 -14312
rect -41215 -14392 -41168 -14328
rect -41104 -14392 -41088 -14328
rect -41215 -14408 -41088 -14392
rect -41215 -14472 -41168 -14408
rect -41104 -14472 -41088 -14408
rect -41215 -14488 -41088 -14472
rect -41215 -14552 -41168 -14488
rect -41104 -14552 -41088 -14488
rect -41215 -14568 -41088 -14552
rect -41215 -14632 -41168 -14568
rect -41104 -14632 -41088 -14568
rect -41215 -14648 -41088 -14632
rect -41215 -14712 -41168 -14648
rect -41104 -14712 -41088 -14648
rect -41215 -14728 -41088 -14712
rect -41215 -14792 -41168 -14728
rect -41104 -14792 -41088 -14728
rect -41215 -14808 -41088 -14792
rect -41215 -14872 -41168 -14808
rect -41104 -14872 -41088 -14808
rect -41215 -14888 -41088 -14872
rect -41215 -14952 -41168 -14888
rect -41104 -14952 -41088 -14888
rect -41215 -14968 -41088 -14952
rect -41215 -15032 -41168 -14968
rect -41104 -15032 -41088 -14968
rect -41215 -15048 -41088 -15032
rect -41215 -15112 -41168 -15048
rect -41104 -15112 -41088 -15048
rect -41215 -15128 -41088 -15112
rect -41215 -15192 -41168 -15128
rect -41104 -15192 -41088 -15128
rect -41215 -15208 -41088 -15192
rect -41215 -15272 -41168 -15208
rect -41104 -15272 -41088 -15208
rect -41215 -15288 -41088 -15272
rect -41215 -15352 -41168 -15288
rect -41104 -15352 -41088 -15288
rect -41215 -15368 -41088 -15352
rect -41215 -15432 -41168 -15368
rect -41104 -15432 -41088 -15368
rect -41215 -15448 -41088 -15432
rect -41215 -15512 -41168 -15448
rect -41104 -15512 -41088 -15448
rect -41215 -15528 -41088 -15512
rect -44335 -15939 -44231 -15561
rect -41215 -15592 -41168 -15528
rect -41104 -15592 -41088 -15528
rect -40925 -9648 -35003 -9639
rect -40925 -15552 -40916 -9648
rect -35012 -15552 -35003 -9648
rect -40925 -15561 -35003 -15552
rect -34896 -9672 -34849 -9608
rect -34785 -9672 -34769 -9608
rect -31697 -9639 -31593 -9261
rect -28577 -9292 -28530 -9228
rect -28466 -9292 -28450 -9228
rect -28287 -3348 -22365 -3339
rect -28287 -9252 -28278 -3348
rect -22374 -9252 -22365 -3348
rect -28287 -9261 -22365 -9252
rect -22258 -3372 -22211 -3308
rect -22147 -3372 -22131 -3308
rect -19059 -3339 -18955 -2961
rect -15939 -2992 -15892 -2928
rect -15828 -2992 -15812 -2928
rect -15649 2952 -9727 2961
rect -15649 -2952 -15640 2952
rect -9736 -2952 -9727 2952
rect -15649 -2961 -9727 -2952
rect -9620 2928 -9573 2992
rect -9509 2928 -9493 2992
rect -6421 2961 -6317 3339
rect -3301 3308 -3254 3372
rect -3190 3308 -3174 3372
rect -3011 9252 2911 9261
rect -3011 3348 -3002 9252
rect 2902 3348 2911 9252
rect -3011 3339 2911 3348
rect 3018 9228 3065 9292
rect 3129 9228 3145 9292
rect 6217 9261 6321 9639
rect 9337 9608 9384 9672
rect 9448 9608 9464 9672
rect 9627 15552 15549 15561
rect 9627 9648 9636 15552
rect 15540 9648 15549 15552
rect 9627 9639 15549 9648
rect 15656 15528 15703 15592
rect 15767 15528 15783 15592
rect 18855 15561 18959 15939
rect 21975 15908 22022 15972
rect 22086 15908 22102 15972
rect 22265 21852 28187 21861
rect 22265 15948 22274 21852
rect 28178 15948 28187 21852
rect 22265 15939 28187 15948
rect 28294 21828 28341 21892
rect 28405 21828 28421 21892
rect 31493 21861 31597 22239
rect 34613 22208 34660 22272
rect 34724 22208 34740 22272
rect 34903 28152 40825 28161
rect 34903 22248 34912 28152
rect 40816 22248 40825 28152
rect 34903 22239 40825 22248
rect 40932 28128 40979 28192
rect 41043 28128 41059 28192
rect 44131 28161 44235 28539
rect 47251 28508 47298 28572
rect 47362 28508 47378 28572
rect 47251 28492 47378 28508
rect 47251 28428 47298 28492
rect 47362 28428 47378 28492
rect 47251 28412 47378 28428
rect 47251 28288 47355 28412
rect 47251 28272 47378 28288
rect 47251 28208 47298 28272
rect 47362 28208 47378 28272
rect 47251 28192 47378 28208
rect 40932 28112 41059 28128
rect 40932 28048 40979 28112
rect 41043 28048 41059 28112
rect 40932 28032 41059 28048
rect 40932 27968 40979 28032
rect 41043 27968 41059 28032
rect 40932 27952 41059 27968
rect 40932 27888 40979 27952
rect 41043 27888 41059 27952
rect 40932 27872 41059 27888
rect 40932 27808 40979 27872
rect 41043 27808 41059 27872
rect 40932 27792 41059 27808
rect 40932 27728 40979 27792
rect 41043 27728 41059 27792
rect 40932 27712 41059 27728
rect 40932 27648 40979 27712
rect 41043 27648 41059 27712
rect 40932 27632 41059 27648
rect 40932 27568 40979 27632
rect 41043 27568 41059 27632
rect 40932 27552 41059 27568
rect 40932 27488 40979 27552
rect 41043 27488 41059 27552
rect 40932 27472 41059 27488
rect 40932 27408 40979 27472
rect 41043 27408 41059 27472
rect 40932 27392 41059 27408
rect 40932 27328 40979 27392
rect 41043 27328 41059 27392
rect 40932 27312 41059 27328
rect 40932 27248 40979 27312
rect 41043 27248 41059 27312
rect 40932 27232 41059 27248
rect 40932 27168 40979 27232
rect 41043 27168 41059 27232
rect 40932 27152 41059 27168
rect 40932 27088 40979 27152
rect 41043 27088 41059 27152
rect 40932 27072 41059 27088
rect 40932 27008 40979 27072
rect 41043 27008 41059 27072
rect 40932 26992 41059 27008
rect 40932 26928 40979 26992
rect 41043 26928 41059 26992
rect 40932 26912 41059 26928
rect 40932 26848 40979 26912
rect 41043 26848 41059 26912
rect 40932 26832 41059 26848
rect 40932 26768 40979 26832
rect 41043 26768 41059 26832
rect 40932 26752 41059 26768
rect 40932 26688 40979 26752
rect 41043 26688 41059 26752
rect 40932 26672 41059 26688
rect 40932 26608 40979 26672
rect 41043 26608 41059 26672
rect 40932 26592 41059 26608
rect 40932 26528 40979 26592
rect 41043 26528 41059 26592
rect 40932 26512 41059 26528
rect 40932 26448 40979 26512
rect 41043 26448 41059 26512
rect 40932 26432 41059 26448
rect 40932 26368 40979 26432
rect 41043 26368 41059 26432
rect 40932 26352 41059 26368
rect 40932 26288 40979 26352
rect 41043 26288 41059 26352
rect 40932 26272 41059 26288
rect 40932 26208 40979 26272
rect 41043 26208 41059 26272
rect 40932 26192 41059 26208
rect 40932 26128 40979 26192
rect 41043 26128 41059 26192
rect 40932 26112 41059 26128
rect 40932 26048 40979 26112
rect 41043 26048 41059 26112
rect 40932 26032 41059 26048
rect 40932 25968 40979 26032
rect 41043 25968 41059 26032
rect 40932 25952 41059 25968
rect 40932 25888 40979 25952
rect 41043 25888 41059 25952
rect 40932 25872 41059 25888
rect 40932 25808 40979 25872
rect 41043 25808 41059 25872
rect 40932 25792 41059 25808
rect 40932 25728 40979 25792
rect 41043 25728 41059 25792
rect 40932 25712 41059 25728
rect 40932 25648 40979 25712
rect 41043 25648 41059 25712
rect 40932 25632 41059 25648
rect 40932 25568 40979 25632
rect 41043 25568 41059 25632
rect 40932 25552 41059 25568
rect 40932 25488 40979 25552
rect 41043 25488 41059 25552
rect 40932 25472 41059 25488
rect 40932 25408 40979 25472
rect 41043 25408 41059 25472
rect 40932 25392 41059 25408
rect 40932 25328 40979 25392
rect 41043 25328 41059 25392
rect 40932 25312 41059 25328
rect 40932 25248 40979 25312
rect 41043 25248 41059 25312
rect 40932 25232 41059 25248
rect 40932 25168 40979 25232
rect 41043 25168 41059 25232
rect 40932 25152 41059 25168
rect 40932 25088 40979 25152
rect 41043 25088 41059 25152
rect 40932 25072 41059 25088
rect 40932 25008 40979 25072
rect 41043 25008 41059 25072
rect 40932 24992 41059 25008
rect 40932 24928 40979 24992
rect 41043 24928 41059 24992
rect 40932 24912 41059 24928
rect 40932 24848 40979 24912
rect 41043 24848 41059 24912
rect 40932 24832 41059 24848
rect 40932 24768 40979 24832
rect 41043 24768 41059 24832
rect 40932 24752 41059 24768
rect 40932 24688 40979 24752
rect 41043 24688 41059 24752
rect 40932 24672 41059 24688
rect 40932 24608 40979 24672
rect 41043 24608 41059 24672
rect 40932 24592 41059 24608
rect 40932 24528 40979 24592
rect 41043 24528 41059 24592
rect 40932 24512 41059 24528
rect 40932 24448 40979 24512
rect 41043 24448 41059 24512
rect 40932 24432 41059 24448
rect 40932 24368 40979 24432
rect 41043 24368 41059 24432
rect 40932 24352 41059 24368
rect 40932 24288 40979 24352
rect 41043 24288 41059 24352
rect 40932 24272 41059 24288
rect 40932 24208 40979 24272
rect 41043 24208 41059 24272
rect 40932 24192 41059 24208
rect 40932 24128 40979 24192
rect 41043 24128 41059 24192
rect 40932 24112 41059 24128
rect 40932 24048 40979 24112
rect 41043 24048 41059 24112
rect 40932 24032 41059 24048
rect 40932 23968 40979 24032
rect 41043 23968 41059 24032
rect 40932 23952 41059 23968
rect 40932 23888 40979 23952
rect 41043 23888 41059 23952
rect 40932 23872 41059 23888
rect 40932 23808 40979 23872
rect 41043 23808 41059 23872
rect 40932 23792 41059 23808
rect 40932 23728 40979 23792
rect 41043 23728 41059 23792
rect 40932 23712 41059 23728
rect 40932 23648 40979 23712
rect 41043 23648 41059 23712
rect 40932 23632 41059 23648
rect 40932 23568 40979 23632
rect 41043 23568 41059 23632
rect 40932 23552 41059 23568
rect 40932 23488 40979 23552
rect 41043 23488 41059 23552
rect 40932 23472 41059 23488
rect 40932 23408 40979 23472
rect 41043 23408 41059 23472
rect 40932 23392 41059 23408
rect 40932 23328 40979 23392
rect 41043 23328 41059 23392
rect 40932 23312 41059 23328
rect 40932 23248 40979 23312
rect 41043 23248 41059 23312
rect 40932 23232 41059 23248
rect 40932 23168 40979 23232
rect 41043 23168 41059 23232
rect 40932 23152 41059 23168
rect 40932 23088 40979 23152
rect 41043 23088 41059 23152
rect 40932 23072 41059 23088
rect 40932 23008 40979 23072
rect 41043 23008 41059 23072
rect 40932 22992 41059 23008
rect 40932 22928 40979 22992
rect 41043 22928 41059 22992
rect 40932 22912 41059 22928
rect 40932 22848 40979 22912
rect 41043 22848 41059 22912
rect 40932 22832 41059 22848
rect 40932 22768 40979 22832
rect 41043 22768 41059 22832
rect 40932 22752 41059 22768
rect 40932 22688 40979 22752
rect 41043 22688 41059 22752
rect 40932 22672 41059 22688
rect 40932 22608 40979 22672
rect 41043 22608 41059 22672
rect 40932 22592 41059 22608
rect 40932 22528 40979 22592
rect 41043 22528 41059 22592
rect 40932 22512 41059 22528
rect 40932 22448 40979 22512
rect 41043 22448 41059 22512
rect 40932 22432 41059 22448
rect 40932 22368 40979 22432
rect 41043 22368 41059 22432
rect 40932 22352 41059 22368
rect 40932 22288 40979 22352
rect 41043 22288 41059 22352
rect 40932 22272 41059 22288
rect 34613 22192 34740 22208
rect 34613 22128 34660 22192
rect 34724 22128 34740 22192
rect 34613 22112 34740 22128
rect 34613 21988 34717 22112
rect 34613 21972 34740 21988
rect 34613 21908 34660 21972
rect 34724 21908 34740 21972
rect 34613 21892 34740 21908
rect 28294 21812 28421 21828
rect 28294 21748 28341 21812
rect 28405 21748 28421 21812
rect 28294 21732 28421 21748
rect 28294 21668 28341 21732
rect 28405 21668 28421 21732
rect 28294 21652 28421 21668
rect 28294 21588 28341 21652
rect 28405 21588 28421 21652
rect 28294 21572 28421 21588
rect 28294 21508 28341 21572
rect 28405 21508 28421 21572
rect 28294 21492 28421 21508
rect 28294 21428 28341 21492
rect 28405 21428 28421 21492
rect 28294 21412 28421 21428
rect 28294 21348 28341 21412
rect 28405 21348 28421 21412
rect 28294 21332 28421 21348
rect 28294 21268 28341 21332
rect 28405 21268 28421 21332
rect 28294 21252 28421 21268
rect 28294 21188 28341 21252
rect 28405 21188 28421 21252
rect 28294 21172 28421 21188
rect 28294 21108 28341 21172
rect 28405 21108 28421 21172
rect 28294 21092 28421 21108
rect 28294 21028 28341 21092
rect 28405 21028 28421 21092
rect 28294 21012 28421 21028
rect 28294 20948 28341 21012
rect 28405 20948 28421 21012
rect 28294 20932 28421 20948
rect 28294 20868 28341 20932
rect 28405 20868 28421 20932
rect 28294 20852 28421 20868
rect 28294 20788 28341 20852
rect 28405 20788 28421 20852
rect 28294 20772 28421 20788
rect 28294 20708 28341 20772
rect 28405 20708 28421 20772
rect 28294 20692 28421 20708
rect 28294 20628 28341 20692
rect 28405 20628 28421 20692
rect 28294 20612 28421 20628
rect 28294 20548 28341 20612
rect 28405 20548 28421 20612
rect 28294 20532 28421 20548
rect 28294 20468 28341 20532
rect 28405 20468 28421 20532
rect 28294 20452 28421 20468
rect 28294 20388 28341 20452
rect 28405 20388 28421 20452
rect 28294 20372 28421 20388
rect 28294 20308 28341 20372
rect 28405 20308 28421 20372
rect 28294 20292 28421 20308
rect 28294 20228 28341 20292
rect 28405 20228 28421 20292
rect 28294 20212 28421 20228
rect 28294 20148 28341 20212
rect 28405 20148 28421 20212
rect 28294 20132 28421 20148
rect 28294 20068 28341 20132
rect 28405 20068 28421 20132
rect 28294 20052 28421 20068
rect 28294 19988 28341 20052
rect 28405 19988 28421 20052
rect 28294 19972 28421 19988
rect 28294 19908 28341 19972
rect 28405 19908 28421 19972
rect 28294 19892 28421 19908
rect 28294 19828 28341 19892
rect 28405 19828 28421 19892
rect 28294 19812 28421 19828
rect 28294 19748 28341 19812
rect 28405 19748 28421 19812
rect 28294 19732 28421 19748
rect 28294 19668 28341 19732
rect 28405 19668 28421 19732
rect 28294 19652 28421 19668
rect 28294 19588 28341 19652
rect 28405 19588 28421 19652
rect 28294 19572 28421 19588
rect 28294 19508 28341 19572
rect 28405 19508 28421 19572
rect 28294 19492 28421 19508
rect 28294 19428 28341 19492
rect 28405 19428 28421 19492
rect 28294 19412 28421 19428
rect 28294 19348 28341 19412
rect 28405 19348 28421 19412
rect 28294 19332 28421 19348
rect 28294 19268 28341 19332
rect 28405 19268 28421 19332
rect 28294 19252 28421 19268
rect 28294 19188 28341 19252
rect 28405 19188 28421 19252
rect 28294 19172 28421 19188
rect 28294 19108 28341 19172
rect 28405 19108 28421 19172
rect 28294 19092 28421 19108
rect 28294 19028 28341 19092
rect 28405 19028 28421 19092
rect 28294 19012 28421 19028
rect 28294 18948 28341 19012
rect 28405 18948 28421 19012
rect 28294 18932 28421 18948
rect 28294 18868 28341 18932
rect 28405 18868 28421 18932
rect 28294 18852 28421 18868
rect 28294 18788 28341 18852
rect 28405 18788 28421 18852
rect 28294 18772 28421 18788
rect 28294 18708 28341 18772
rect 28405 18708 28421 18772
rect 28294 18692 28421 18708
rect 28294 18628 28341 18692
rect 28405 18628 28421 18692
rect 28294 18612 28421 18628
rect 28294 18548 28341 18612
rect 28405 18548 28421 18612
rect 28294 18532 28421 18548
rect 28294 18468 28341 18532
rect 28405 18468 28421 18532
rect 28294 18452 28421 18468
rect 28294 18388 28341 18452
rect 28405 18388 28421 18452
rect 28294 18372 28421 18388
rect 28294 18308 28341 18372
rect 28405 18308 28421 18372
rect 28294 18292 28421 18308
rect 28294 18228 28341 18292
rect 28405 18228 28421 18292
rect 28294 18212 28421 18228
rect 28294 18148 28341 18212
rect 28405 18148 28421 18212
rect 28294 18132 28421 18148
rect 28294 18068 28341 18132
rect 28405 18068 28421 18132
rect 28294 18052 28421 18068
rect 28294 17988 28341 18052
rect 28405 17988 28421 18052
rect 28294 17972 28421 17988
rect 28294 17908 28341 17972
rect 28405 17908 28421 17972
rect 28294 17892 28421 17908
rect 28294 17828 28341 17892
rect 28405 17828 28421 17892
rect 28294 17812 28421 17828
rect 28294 17748 28341 17812
rect 28405 17748 28421 17812
rect 28294 17732 28421 17748
rect 28294 17668 28341 17732
rect 28405 17668 28421 17732
rect 28294 17652 28421 17668
rect 28294 17588 28341 17652
rect 28405 17588 28421 17652
rect 28294 17572 28421 17588
rect 28294 17508 28341 17572
rect 28405 17508 28421 17572
rect 28294 17492 28421 17508
rect 28294 17428 28341 17492
rect 28405 17428 28421 17492
rect 28294 17412 28421 17428
rect 28294 17348 28341 17412
rect 28405 17348 28421 17412
rect 28294 17332 28421 17348
rect 28294 17268 28341 17332
rect 28405 17268 28421 17332
rect 28294 17252 28421 17268
rect 28294 17188 28341 17252
rect 28405 17188 28421 17252
rect 28294 17172 28421 17188
rect 28294 17108 28341 17172
rect 28405 17108 28421 17172
rect 28294 17092 28421 17108
rect 28294 17028 28341 17092
rect 28405 17028 28421 17092
rect 28294 17012 28421 17028
rect 28294 16948 28341 17012
rect 28405 16948 28421 17012
rect 28294 16932 28421 16948
rect 28294 16868 28341 16932
rect 28405 16868 28421 16932
rect 28294 16852 28421 16868
rect 28294 16788 28341 16852
rect 28405 16788 28421 16852
rect 28294 16772 28421 16788
rect 28294 16708 28341 16772
rect 28405 16708 28421 16772
rect 28294 16692 28421 16708
rect 28294 16628 28341 16692
rect 28405 16628 28421 16692
rect 28294 16612 28421 16628
rect 28294 16548 28341 16612
rect 28405 16548 28421 16612
rect 28294 16532 28421 16548
rect 28294 16468 28341 16532
rect 28405 16468 28421 16532
rect 28294 16452 28421 16468
rect 28294 16388 28341 16452
rect 28405 16388 28421 16452
rect 28294 16372 28421 16388
rect 28294 16308 28341 16372
rect 28405 16308 28421 16372
rect 28294 16292 28421 16308
rect 28294 16228 28341 16292
rect 28405 16228 28421 16292
rect 28294 16212 28421 16228
rect 28294 16148 28341 16212
rect 28405 16148 28421 16212
rect 28294 16132 28421 16148
rect 28294 16068 28341 16132
rect 28405 16068 28421 16132
rect 28294 16052 28421 16068
rect 28294 15988 28341 16052
rect 28405 15988 28421 16052
rect 28294 15972 28421 15988
rect 21975 15892 22102 15908
rect 21975 15828 22022 15892
rect 22086 15828 22102 15892
rect 21975 15812 22102 15828
rect 21975 15688 22079 15812
rect 21975 15672 22102 15688
rect 21975 15608 22022 15672
rect 22086 15608 22102 15672
rect 21975 15592 22102 15608
rect 15656 15512 15783 15528
rect 15656 15448 15703 15512
rect 15767 15448 15783 15512
rect 15656 15432 15783 15448
rect 15656 15368 15703 15432
rect 15767 15368 15783 15432
rect 15656 15352 15783 15368
rect 15656 15288 15703 15352
rect 15767 15288 15783 15352
rect 15656 15272 15783 15288
rect 15656 15208 15703 15272
rect 15767 15208 15783 15272
rect 15656 15192 15783 15208
rect 15656 15128 15703 15192
rect 15767 15128 15783 15192
rect 15656 15112 15783 15128
rect 15656 15048 15703 15112
rect 15767 15048 15783 15112
rect 15656 15032 15783 15048
rect 15656 14968 15703 15032
rect 15767 14968 15783 15032
rect 15656 14952 15783 14968
rect 15656 14888 15703 14952
rect 15767 14888 15783 14952
rect 15656 14872 15783 14888
rect 15656 14808 15703 14872
rect 15767 14808 15783 14872
rect 15656 14792 15783 14808
rect 15656 14728 15703 14792
rect 15767 14728 15783 14792
rect 15656 14712 15783 14728
rect 15656 14648 15703 14712
rect 15767 14648 15783 14712
rect 15656 14632 15783 14648
rect 15656 14568 15703 14632
rect 15767 14568 15783 14632
rect 15656 14552 15783 14568
rect 15656 14488 15703 14552
rect 15767 14488 15783 14552
rect 15656 14472 15783 14488
rect 15656 14408 15703 14472
rect 15767 14408 15783 14472
rect 15656 14392 15783 14408
rect 15656 14328 15703 14392
rect 15767 14328 15783 14392
rect 15656 14312 15783 14328
rect 15656 14248 15703 14312
rect 15767 14248 15783 14312
rect 15656 14232 15783 14248
rect 15656 14168 15703 14232
rect 15767 14168 15783 14232
rect 15656 14152 15783 14168
rect 15656 14088 15703 14152
rect 15767 14088 15783 14152
rect 15656 14072 15783 14088
rect 15656 14008 15703 14072
rect 15767 14008 15783 14072
rect 15656 13992 15783 14008
rect 15656 13928 15703 13992
rect 15767 13928 15783 13992
rect 15656 13912 15783 13928
rect 15656 13848 15703 13912
rect 15767 13848 15783 13912
rect 15656 13832 15783 13848
rect 15656 13768 15703 13832
rect 15767 13768 15783 13832
rect 15656 13752 15783 13768
rect 15656 13688 15703 13752
rect 15767 13688 15783 13752
rect 15656 13672 15783 13688
rect 15656 13608 15703 13672
rect 15767 13608 15783 13672
rect 15656 13592 15783 13608
rect 15656 13528 15703 13592
rect 15767 13528 15783 13592
rect 15656 13512 15783 13528
rect 15656 13448 15703 13512
rect 15767 13448 15783 13512
rect 15656 13432 15783 13448
rect 15656 13368 15703 13432
rect 15767 13368 15783 13432
rect 15656 13352 15783 13368
rect 15656 13288 15703 13352
rect 15767 13288 15783 13352
rect 15656 13272 15783 13288
rect 15656 13208 15703 13272
rect 15767 13208 15783 13272
rect 15656 13192 15783 13208
rect 15656 13128 15703 13192
rect 15767 13128 15783 13192
rect 15656 13112 15783 13128
rect 15656 13048 15703 13112
rect 15767 13048 15783 13112
rect 15656 13032 15783 13048
rect 15656 12968 15703 13032
rect 15767 12968 15783 13032
rect 15656 12952 15783 12968
rect 15656 12888 15703 12952
rect 15767 12888 15783 12952
rect 15656 12872 15783 12888
rect 15656 12808 15703 12872
rect 15767 12808 15783 12872
rect 15656 12792 15783 12808
rect 15656 12728 15703 12792
rect 15767 12728 15783 12792
rect 15656 12712 15783 12728
rect 15656 12648 15703 12712
rect 15767 12648 15783 12712
rect 15656 12632 15783 12648
rect 15656 12568 15703 12632
rect 15767 12568 15783 12632
rect 15656 12552 15783 12568
rect 15656 12488 15703 12552
rect 15767 12488 15783 12552
rect 15656 12472 15783 12488
rect 15656 12408 15703 12472
rect 15767 12408 15783 12472
rect 15656 12392 15783 12408
rect 15656 12328 15703 12392
rect 15767 12328 15783 12392
rect 15656 12312 15783 12328
rect 15656 12248 15703 12312
rect 15767 12248 15783 12312
rect 15656 12232 15783 12248
rect 15656 12168 15703 12232
rect 15767 12168 15783 12232
rect 15656 12152 15783 12168
rect 15656 12088 15703 12152
rect 15767 12088 15783 12152
rect 15656 12072 15783 12088
rect 15656 12008 15703 12072
rect 15767 12008 15783 12072
rect 15656 11992 15783 12008
rect 15656 11928 15703 11992
rect 15767 11928 15783 11992
rect 15656 11912 15783 11928
rect 15656 11848 15703 11912
rect 15767 11848 15783 11912
rect 15656 11832 15783 11848
rect 15656 11768 15703 11832
rect 15767 11768 15783 11832
rect 15656 11752 15783 11768
rect 15656 11688 15703 11752
rect 15767 11688 15783 11752
rect 15656 11672 15783 11688
rect 15656 11608 15703 11672
rect 15767 11608 15783 11672
rect 15656 11592 15783 11608
rect 15656 11528 15703 11592
rect 15767 11528 15783 11592
rect 15656 11512 15783 11528
rect 15656 11448 15703 11512
rect 15767 11448 15783 11512
rect 15656 11432 15783 11448
rect 15656 11368 15703 11432
rect 15767 11368 15783 11432
rect 15656 11352 15783 11368
rect 15656 11288 15703 11352
rect 15767 11288 15783 11352
rect 15656 11272 15783 11288
rect 15656 11208 15703 11272
rect 15767 11208 15783 11272
rect 15656 11192 15783 11208
rect 15656 11128 15703 11192
rect 15767 11128 15783 11192
rect 15656 11112 15783 11128
rect 15656 11048 15703 11112
rect 15767 11048 15783 11112
rect 15656 11032 15783 11048
rect 15656 10968 15703 11032
rect 15767 10968 15783 11032
rect 15656 10952 15783 10968
rect 15656 10888 15703 10952
rect 15767 10888 15783 10952
rect 15656 10872 15783 10888
rect 15656 10808 15703 10872
rect 15767 10808 15783 10872
rect 15656 10792 15783 10808
rect 15656 10728 15703 10792
rect 15767 10728 15783 10792
rect 15656 10712 15783 10728
rect 15656 10648 15703 10712
rect 15767 10648 15783 10712
rect 15656 10632 15783 10648
rect 15656 10568 15703 10632
rect 15767 10568 15783 10632
rect 15656 10552 15783 10568
rect 15656 10488 15703 10552
rect 15767 10488 15783 10552
rect 15656 10472 15783 10488
rect 15656 10408 15703 10472
rect 15767 10408 15783 10472
rect 15656 10392 15783 10408
rect 15656 10328 15703 10392
rect 15767 10328 15783 10392
rect 15656 10312 15783 10328
rect 15656 10248 15703 10312
rect 15767 10248 15783 10312
rect 15656 10232 15783 10248
rect 15656 10168 15703 10232
rect 15767 10168 15783 10232
rect 15656 10152 15783 10168
rect 15656 10088 15703 10152
rect 15767 10088 15783 10152
rect 15656 10072 15783 10088
rect 15656 10008 15703 10072
rect 15767 10008 15783 10072
rect 15656 9992 15783 10008
rect 15656 9928 15703 9992
rect 15767 9928 15783 9992
rect 15656 9912 15783 9928
rect 15656 9848 15703 9912
rect 15767 9848 15783 9912
rect 15656 9832 15783 9848
rect 15656 9768 15703 9832
rect 15767 9768 15783 9832
rect 15656 9752 15783 9768
rect 15656 9688 15703 9752
rect 15767 9688 15783 9752
rect 15656 9672 15783 9688
rect 9337 9592 9464 9608
rect 9337 9528 9384 9592
rect 9448 9528 9464 9592
rect 9337 9512 9464 9528
rect 9337 9388 9441 9512
rect 9337 9372 9464 9388
rect 9337 9308 9384 9372
rect 9448 9308 9464 9372
rect 9337 9292 9464 9308
rect 3018 9212 3145 9228
rect 3018 9148 3065 9212
rect 3129 9148 3145 9212
rect 3018 9132 3145 9148
rect 3018 9068 3065 9132
rect 3129 9068 3145 9132
rect 3018 9052 3145 9068
rect 3018 8988 3065 9052
rect 3129 8988 3145 9052
rect 3018 8972 3145 8988
rect 3018 8908 3065 8972
rect 3129 8908 3145 8972
rect 3018 8892 3145 8908
rect 3018 8828 3065 8892
rect 3129 8828 3145 8892
rect 3018 8812 3145 8828
rect 3018 8748 3065 8812
rect 3129 8748 3145 8812
rect 3018 8732 3145 8748
rect 3018 8668 3065 8732
rect 3129 8668 3145 8732
rect 3018 8652 3145 8668
rect 3018 8588 3065 8652
rect 3129 8588 3145 8652
rect 3018 8572 3145 8588
rect 3018 8508 3065 8572
rect 3129 8508 3145 8572
rect 3018 8492 3145 8508
rect 3018 8428 3065 8492
rect 3129 8428 3145 8492
rect 3018 8412 3145 8428
rect 3018 8348 3065 8412
rect 3129 8348 3145 8412
rect 3018 8332 3145 8348
rect 3018 8268 3065 8332
rect 3129 8268 3145 8332
rect 3018 8252 3145 8268
rect 3018 8188 3065 8252
rect 3129 8188 3145 8252
rect 3018 8172 3145 8188
rect 3018 8108 3065 8172
rect 3129 8108 3145 8172
rect 3018 8092 3145 8108
rect 3018 8028 3065 8092
rect 3129 8028 3145 8092
rect 3018 8012 3145 8028
rect 3018 7948 3065 8012
rect 3129 7948 3145 8012
rect 3018 7932 3145 7948
rect 3018 7868 3065 7932
rect 3129 7868 3145 7932
rect 3018 7852 3145 7868
rect 3018 7788 3065 7852
rect 3129 7788 3145 7852
rect 3018 7772 3145 7788
rect 3018 7708 3065 7772
rect 3129 7708 3145 7772
rect 3018 7692 3145 7708
rect 3018 7628 3065 7692
rect 3129 7628 3145 7692
rect 3018 7612 3145 7628
rect 3018 7548 3065 7612
rect 3129 7548 3145 7612
rect 3018 7532 3145 7548
rect 3018 7468 3065 7532
rect 3129 7468 3145 7532
rect 3018 7452 3145 7468
rect 3018 7388 3065 7452
rect 3129 7388 3145 7452
rect 3018 7372 3145 7388
rect 3018 7308 3065 7372
rect 3129 7308 3145 7372
rect 3018 7292 3145 7308
rect 3018 7228 3065 7292
rect 3129 7228 3145 7292
rect 3018 7212 3145 7228
rect 3018 7148 3065 7212
rect 3129 7148 3145 7212
rect 3018 7132 3145 7148
rect 3018 7068 3065 7132
rect 3129 7068 3145 7132
rect 3018 7052 3145 7068
rect 3018 6988 3065 7052
rect 3129 6988 3145 7052
rect 3018 6972 3145 6988
rect 3018 6908 3065 6972
rect 3129 6908 3145 6972
rect 3018 6892 3145 6908
rect 3018 6828 3065 6892
rect 3129 6828 3145 6892
rect 3018 6812 3145 6828
rect 3018 6748 3065 6812
rect 3129 6748 3145 6812
rect 3018 6732 3145 6748
rect 3018 6668 3065 6732
rect 3129 6668 3145 6732
rect 3018 6652 3145 6668
rect 3018 6588 3065 6652
rect 3129 6588 3145 6652
rect 3018 6572 3145 6588
rect 3018 6508 3065 6572
rect 3129 6508 3145 6572
rect 3018 6492 3145 6508
rect 3018 6428 3065 6492
rect 3129 6428 3145 6492
rect 3018 6412 3145 6428
rect 3018 6348 3065 6412
rect 3129 6348 3145 6412
rect 3018 6332 3145 6348
rect 3018 6268 3065 6332
rect 3129 6268 3145 6332
rect 3018 6252 3145 6268
rect 3018 6188 3065 6252
rect 3129 6188 3145 6252
rect 3018 6172 3145 6188
rect 3018 6108 3065 6172
rect 3129 6108 3145 6172
rect 3018 6092 3145 6108
rect 3018 6028 3065 6092
rect 3129 6028 3145 6092
rect 3018 6012 3145 6028
rect 3018 5948 3065 6012
rect 3129 5948 3145 6012
rect 3018 5932 3145 5948
rect 3018 5868 3065 5932
rect 3129 5868 3145 5932
rect 3018 5852 3145 5868
rect 3018 5788 3065 5852
rect 3129 5788 3145 5852
rect 3018 5772 3145 5788
rect 3018 5708 3065 5772
rect 3129 5708 3145 5772
rect 3018 5692 3145 5708
rect 3018 5628 3065 5692
rect 3129 5628 3145 5692
rect 3018 5612 3145 5628
rect 3018 5548 3065 5612
rect 3129 5548 3145 5612
rect 3018 5532 3145 5548
rect 3018 5468 3065 5532
rect 3129 5468 3145 5532
rect 3018 5452 3145 5468
rect 3018 5388 3065 5452
rect 3129 5388 3145 5452
rect 3018 5372 3145 5388
rect 3018 5308 3065 5372
rect 3129 5308 3145 5372
rect 3018 5292 3145 5308
rect 3018 5228 3065 5292
rect 3129 5228 3145 5292
rect 3018 5212 3145 5228
rect 3018 5148 3065 5212
rect 3129 5148 3145 5212
rect 3018 5132 3145 5148
rect 3018 5068 3065 5132
rect 3129 5068 3145 5132
rect 3018 5052 3145 5068
rect 3018 4988 3065 5052
rect 3129 4988 3145 5052
rect 3018 4972 3145 4988
rect 3018 4908 3065 4972
rect 3129 4908 3145 4972
rect 3018 4892 3145 4908
rect 3018 4828 3065 4892
rect 3129 4828 3145 4892
rect 3018 4812 3145 4828
rect 3018 4748 3065 4812
rect 3129 4748 3145 4812
rect 3018 4732 3145 4748
rect 3018 4668 3065 4732
rect 3129 4668 3145 4732
rect 3018 4652 3145 4668
rect 3018 4588 3065 4652
rect 3129 4588 3145 4652
rect 3018 4572 3145 4588
rect 3018 4508 3065 4572
rect 3129 4508 3145 4572
rect 3018 4492 3145 4508
rect 3018 4428 3065 4492
rect 3129 4428 3145 4492
rect 3018 4412 3145 4428
rect 3018 4348 3065 4412
rect 3129 4348 3145 4412
rect 3018 4332 3145 4348
rect 3018 4268 3065 4332
rect 3129 4268 3145 4332
rect 3018 4252 3145 4268
rect 3018 4188 3065 4252
rect 3129 4188 3145 4252
rect 3018 4172 3145 4188
rect 3018 4108 3065 4172
rect 3129 4108 3145 4172
rect 3018 4092 3145 4108
rect 3018 4028 3065 4092
rect 3129 4028 3145 4092
rect 3018 4012 3145 4028
rect 3018 3948 3065 4012
rect 3129 3948 3145 4012
rect 3018 3932 3145 3948
rect 3018 3868 3065 3932
rect 3129 3868 3145 3932
rect 3018 3852 3145 3868
rect 3018 3788 3065 3852
rect 3129 3788 3145 3852
rect 3018 3772 3145 3788
rect 3018 3708 3065 3772
rect 3129 3708 3145 3772
rect 3018 3692 3145 3708
rect 3018 3628 3065 3692
rect 3129 3628 3145 3692
rect 3018 3612 3145 3628
rect 3018 3548 3065 3612
rect 3129 3548 3145 3612
rect 3018 3532 3145 3548
rect 3018 3468 3065 3532
rect 3129 3468 3145 3532
rect 3018 3452 3145 3468
rect 3018 3388 3065 3452
rect 3129 3388 3145 3452
rect 3018 3372 3145 3388
rect -3301 3292 -3174 3308
rect -3301 3228 -3254 3292
rect -3190 3228 -3174 3292
rect -3301 3212 -3174 3228
rect -3301 3088 -3197 3212
rect -3301 3072 -3174 3088
rect -3301 3008 -3254 3072
rect -3190 3008 -3174 3072
rect -3301 2992 -3174 3008
rect -9620 2912 -9493 2928
rect -9620 2848 -9573 2912
rect -9509 2848 -9493 2912
rect -9620 2832 -9493 2848
rect -9620 2768 -9573 2832
rect -9509 2768 -9493 2832
rect -9620 2752 -9493 2768
rect -9620 2688 -9573 2752
rect -9509 2688 -9493 2752
rect -9620 2672 -9493 2688
rect -9620 2608 -9573 2672
rect -9509 2608 -9493 2672
rect -9620 2592 -9493 2608
rect -9620 2528 -9573 2592
rect -9509 2528 -9493 2592
rect -9620 2512 -9493 2528
rect -9620 2448 -9573 2512
rect -9509 2448 -9493 2512
rect -9620 2432 -9493 2448
rect -9620 2368 -9573 2432
rect -9509 2368 -9493 2432
rect -9620 2352 -9493 2368
rect -9620 2288 -9573 2352
rect -9509 2288 -9493 2352
rect -9620 2272 -9493 2288
rect -9620 2208 -9573 2272
rect -9509 2208 -9493 2272
rect -9620 2192 -9493 2208
rect -9620 2128 -9573 2192
rect -9509 2128 -9493 2192
rect -9620 2112 -9493 2128
rect -9620 2048 -9573 2112
rect -9509 2048 -9493 2112
rect -9620 2032 -9493 2048
rect -9620 1968 -9573 2032
rect -9509 1968 -9493 2032
rect -9620 1952 -9493 1968
rect -9620 1888 -9573 1952
rect -9509 1888 -9493 1952
rect -9620 1872 -9493 1888
rect -9620 1808 -9573 1872
rect -9509 1808 -9493 1872
rect -9620 1792 -9493 1808
rect -9620 1728 -9573 1792
rect -9509 1728 -9493 1792
rect -9620 1712 -9493 1728
rect -9620 1648 -9573 1712
rect -9509 1648 -9493 1712
rect -9620 1632 -9493 1648
rect -9620 1568 -9573 1632
rect -9509 1568 -9493 1632
rect -9620 1552 -9493 1568
rect -9620 1488 -9573 1552
rect -9509 1488 -9493 1552
rect -9620 1472 -9493 1488
rect -9620 1408 -9573 1472
rect -9509 1408 -9493 1472
rect -9620 1392 -9493 1408
rect -9620 1328 -9573 1392
rect -9509 1328 -9493 1392
rect -9620 1312 -9493 1328
rect -9620 1248 -9573 1312
rect -9509 1248 -9493 1312
rect -9620 1232 -9493 1248
rect -9620 1168 -9573 1232
rect -9509 1168 -9493 1232
rect -9620 1152 -9493 1168
rect -9620 1088 -9573 1152
rect -9509 1088 -9493 1152
rect -9620 1072 -9493 1088
rect -9620 1008 -9573 1072
rect -9509 1008 -9493 1072
rect -9620 992 -9493 1008
rect -9620 928 -9573 992
rect -9509 928 -9493 992
rect -9620 912 -9493 928
rect -9620 848 -9573 912
rect -9509 848 -9493 912
rect -9620 832 -9493 848
rect -9620 768 -9573 832
rect -9509 768 -9493 832
rect -9620 752 -9493 768
rect -9620 688 -9573 752
rect -9509 688 -9493 752
rect -9620 672 -9493 688
rect -9620 608 -9573 672
rect -9509 608 -9493 672
rect -9620 592 -9493 608
rect -9620 528 -9573 592
rect -9509 528 -9493 592
rect -9620 512 -9493 528
rect -9620 448 -9573 512
rect -9509 448 -9493 512
rect -9620 432 -9493 448
rect -9620 368 -9573 432
rect -9509 368 -9493 432
rect -9620 352 -9493 368
rect -9620 288 -9573 352
rect -9509 288 -9493 352
rect -9620 272 -9493 288
rect -9620 208 -9573 272
rect -9509 208 -9493 272
rect -9620 192 -9493 208
rect -9620 128 -9573 192
rect -9509 128 -9493 192
rect -9620 112 -9493 128
rect -9620 48 -9573 112
rect -9509 48 -9493 112
rect -9620 32 -9493 48
rect -9620 -32 -9573 32
rect -9509 -32 -9493 32
rect -9620 -48 -9493 -32
rect -9620 -112 -9573 -48
rect -9509 -112 -9493 -48
rect -9620 -128 -9493 -112
rect -9620 -192 -9573 -128
rect -9509 -192 -9493 -128
rect -9620 -208 -9493 -192
rect -9620 -272 -9573 -208
rect -9509 -272 -9493 -208
rect -9620 -288 -9493 -272
rect -9620 -352 -9573 -288
rect -9509 -352 -9493 -288
rect -9620 -368 -9493 -352
rect -9620 -432 -9573 -368
rect -9509 -432 -9493 -368
rect -9620 -448 -9493 -432
rect -9620 -512 -9573 -448
rect -9509 -512 -9493 -448
rect -9620 -528 -9493 -512
rect -9620 -592 -9573 -528
rect -9509 -592 -9493 -528
rect -9620 -608 -9493 -592
rect -9620 -672 -9573 -608
rect -9509 -672 -9493 -608
rect -9620 -688 -9493 -672
rect -9620 -752 -9573 -688
rect -9509 -752 -9493 -688
rect -9620 -768 -9493 -752
rect -9620 -832 -9573 -768
rect -9509 -832 -9493 -768
rect -9620 -848 -9493 -832
rect -9620 -912 -9573 -848
rect -9509 -912 -9493 -848
rect -9620 -928 -9493 -912
rect -9620 -992 -9573 -928
rect -9509 -992 -9493 -928
rect -9620 -1008 -9493 -992
rect -9620 -1072 -9573 -1008
rect -9509 -1072 -9493 -1008
rect -9620 -1088 -9493 -1072
rect -9620 -1152 -9573 -1088
rect -9509 -1152 -9493 -1088
rect -9620 -1168 -9493 -1152
rect -9620 -1232 -9573 -1168
rect -9509 -1232 -9493 -1168
rect -9620 -1248 -9493 -1232
rect -9620 -1312 -9573 -1248
rect -9509 -1312 -9493 -1248
rect -9620 -1328 -9493 -1312
rect -9620 -1392 -9573 -1328
rect -9509 -1392 -9493 -1328
rect -9620 -1408 -9493 -1392
rect -9620 -1472 -9573 -1408
rect -9509 -1472 -9493 -1408
rect -9620 -1488 -9493 -1472
rect -9620 -1552 -9573 -1488
rect -9509 -1552 -9493 -1488
rect -9620 -1568 -9493 -1552
rect -9620 -1632 -9573 -1568
rect -9509 -1632 -9493 -1568
rect -9620 -1648 -9493 -1632
rect -9620 -1712 -9573 -1648
rect -9509 -1712 -9493 -1648
rect -9620 -1728 -9493 -1712
rect -9620 -1792 -9573 -1728
rect -9509 -1792 -9493 -1728
rect -9620 -1808 -9493 -1792
rect -9620 -1872 -9573 -1808
rect -9509 -1872 -9493 -1808
rect -9620 -1888 -9493 -1872
rect -9620 -1952 -9573 -1888
rect -9509 -1952 -9493 -1888
rect -9620 -1968 -9493 -1952
rect -9620 -2032 -9573 -1968
rect -9509 -2032 -9493 -1968
rect -9620 -2048 -9493 -2032
rect -9620 -2112 -9573 -2048
rect -9509 -2112 -9493 -2048
rect -9620 -2128 -9493 -2112
rect -9620 -2192 -9573 -2128
rect -9509 -2192 -9493 -2128
rect -9620 -2208 -9493 -2192
rect -9620 -2272 -9573 -2208
rect -9509 -2272 -9493 -2208
rect -9620 -2288 -9493 -2272
rect -9620 -2352 -9573 -2288
rect -9509 -2352 -9493 -2288
rect -9620 -2368 -9493 -2352
rect -9620 -2432 -9573 -2368
rect -9509 -2432 -9493 -2368
rect -9620 -2448 -9493 -2432
rect -9620 -2512 -9573 -2448
rect -9509 -2512 -9493 -2448
rect -9620 -2528 -9493 -2512
rect -9620 -2592 -9573 -2528
rect -9509 -2592 -9493 -2528
rect -9620 -2608 -9493 -2592
rect -9620 -2672 -9573 -2608
rect -9509 -2672 -9493 -2608
rect -9620 -2688 -9493 -2672
rect -9620 -2752 -9573 -2688
rect -9509 -2752 -9493 -2688
rect -9620 -2768 -9493 -2752
rect -9620 -2832 -9573 -2768
rect -9509 -2832 -9493 -2768
rect -9620 -2848 -9493 -2832
rect -9620 -2912 -9573 -2848
rect -9509 -2912 -9493 -2848
rect -9620 -2928 -9493 -2912
rect -15939 -3008 -15812 -2992
rect -15939 -3072 -15892 -3008
rect -15828 -3072 -15812 -3008
rect -15939 -3088 -15812 -3072
rect -15939 -3212 -15835 -3088
rect -15939 -3228 -15812 -3212
rect -15939 -3292 -15892 -3228
rect -15828 -3292 -15812 -3228
rect -15939 -3308 -15812 -3292
rect -22258 -3388 -22131 -3372
rect -22258 -3452 -22211 -3388
rect -22147 -3452 -22131 -3388
rect -22258 -3468 -22131 -3452
rect -22258 -3532 -22211 -3468
rect -22147 -3532 -22131 -3468
rect -22258 -3548 -22131 -3532
rect -22258 -3612 -22211 -3548
rect -22147 -3612 -22131 -3548
rect -22258 -3628 -22131 -3612
rect -22258 -3692 -22211 -3628
rect -22147 -3692 -22131 -3628
rect -22258 -3708 -22131 -3692
rect -22258 -3772 -22211 -3708
rect -22147 -3772 -22131 -3708
rect -22258 -3788 -22131 -3772
rect -22258 -3852 -22211 -3788
rect -22147 -3852 -22131 -3788
rect -22258 -3868 -22131 -3852
rect -22258 -3932 -22211 -3868
rect -22147 -3932 -22131 -3868
rect -22258 -3948 -22131 -3932
rect -22258 -4012 -22211 -3948
rect -22147 -4012 -22131 -3948
rect -22258 -4028 -22131 -4012
rect -22258 -4092 -22211 -4028
rect -22147 -4092 -22131 -4028
rect -22258 -4108 -22131 -4092
rect -22258 -4172 -22211 -4108
rect -22147 -4172 -22131 -4108
rect -22258 -4188 -22131 -4172
rect -22258 -4252 -22211 -4188
rect -22147 -4252 -22131 -4188
rect -22258 -4268 -22131 -4252
rect -22258 -4332 -22211 -4268
rect -22147 -4332 -22131 -4268
rect -22258 -4348 -22131 -4332
rect -22258 -4412 -22211 -4348
rect -22147 -4412 -22131 -4348
rect -22258 -4428 -22131 -4412
rect -22258 -4492 -22211 -4428
rect -22147 -4492 -22131 -4428
rect -22258 -4508 -22131 -4492
rect -22258 -4572 -22211 -4508
rect -22147 -4572 -22131 -4508
rect -22258 -4588 -22131 -4572
rect -22258 -4652 -22211 -4588
rect -22147 -4652 -22131 -4588
rect -22258 -4668 -22131 -4652
rect -22258 -4732 -22211 -4668
rect -22147 -4732 -22131 -4668
rect -22258 -4748 -22131 -4732
rect -22258 -4812 -22211 -4748
rect -22147 -4812 -22131 -4748
rect -22258 -4828 -22131 -4812
rect -22258 -4892 -22211 -4828
rect -22147 -4892 -22131 -4828
rect -22258 -4908 -22131 -4892
rect -22258 -4972 -22211 -4908
rect -22147 -4972 -22131 -4908
rect -22258 -4988 -22131 -4972
rect -22258 -5052 -22211 -4988
rect -22147 -5052 -22131 -4988
rect -22258 -5068 -22131 -5052
rect -22258 -5132 -22211 -5068
rect -22147 -5132 -22131 -5068
rect -22258 -5148 -22131 -5132
rect -22258 -5212 -22211 -5148
rect -22147 -5212 -22131 -5148
rect -22258 -5228 -22131 -5212
rect -22258 -5292 -22211 -5228
rect -22147 -5292 -22131 -5228
rect -22258 -5308 -22131 -5292
rect -22258 -5372 -22211 -5308
rect -22147 -5372 -22131 -5308
rect -22258 -5388 -22131 -5372
rect -22258 -5452 -22211 -5388
rect -22147 -5452 -22131 -5388
rect -22258 -5468 -22131 -5452
rect -22258 -5532 -22211 -5468
rect -22147 -5532 -22131 -5468
rect -22258 -5548 -22131 -5532
rect -22258 -5612 -22211 -5548
rect -22147 -5612 -22131 -5548
rect -22258 -5628 -22131 -5612
rect -22258 -5692 -22211 -5628
rect -22147 -5692 -22131 -5628
rect -22258 -5708 -22131 -5692
rect -22258 -5772 -22211 -5708
rect -22147 -5772 -22131 -5708
rect -22258 -5788 -22131 -5772
rect -22258 -5852 -22211 -5788
rect -22147 -5852 -22131 -5788
rect -22258 -5868 -22131 -5852
rect -22258 -5932 -22211 -5868
rect -22147 -5932 -22131 -5868
rect -22258 -5948 -22131 -5932
rect -22258 -6012 -22211 -5948
rect -22147 -6012 -22131 -5948
rect -22258 -6028 -22131 -6012
rect -22258 -6092 -22211 -6028
rect -22147 -6092 -22131 -6028
rect -22258 -6108 -22131 -6092
rect -22258 -6172 -22211 -6108
rect -22147 -6172 -22131 -6108
rect -22258 -6188 -22131 -6172
rect -22258 -6252 -22211 -6188
rect -22147 -6252 -22131 -6188
rect -22258 -6268 -22131 -6252
rect -22258 -6332 -22211 -6268
rect -22147 -6332 -22131 -6268
rect -22258 -6348 -22131 -6332
rect -22258 -6412 -22211 -6348
rect -22147 -6412 -22131 -6348
rect -22258 -6428 -22131 -6412
rect -22258 -6492 -22211 -6428
rect -22147 -6492 -22131 -6428
rect -22258 -6508 -22131 -6492
rect -22258 -6572 -22211 -6508
rect -22147 -6572 -22131 -6508
rect -22258 -6588 -22131 -6572
rect -22258 -6652 -22211 -6588
rect -22147 -6652 -22131 -6588
rect -22258 -6668 -22131 -6652
rect -22258 -6732 -22211 -6668
rect -22147 -6732 -22131 -6668
rect -22258 -6748 -22131 -6732
rect -22258 -6812 -22211 -6748
rect -22147 -6812 -22131 -6748
rect -22258 -6828 -22131 -6812
rect -22258 -6892 -22211 -6828
rect -22147 -6892 -22131 -6828
rect -22258 -6908 -22131 -6892
rect -22258 -6972 -22211 -6908
rect -22147 -6972 -22131 -6908
rect -22258 -6988 -22131 -6972
rect -22258 -7052 -22211 -6988
rect -22147 -7052 -22131 -6988
rect -22258 -7068 -22131 -7052
rect -22258 -7132 -22211 -7068
rect -22147 -7132 -22131 -7068
rect -22258 -7148 -22131 -7132
rect -22258 -7212 -22211 -7148
rect -22147 -7212 -22131 -7148
rect -22258 -7228 -22131 -7212
rect -22258 -7292 -22211 -7228
rect -22147 -7292 -22131 -7228
rect -22258 -7308 -22131 -7292
rect -22258 -7372 -22211 -7308
rect -22147 -7372 -22131 -7308
rect -22258 -7388 -22131 -7372
rect -22258 -7452 -22211 -7388
rect -22147 -7452 -22131 -7388
rect -22258 -7468 -22131 -7452
rect -22258 -7532 -22211 -7468
rect -22147 -7532 -22131 -7468
rect -22258 -7548 -22131 -7532
rect -22258 -7612 -22211 -7548
rect -22147 -7612 -22131 -7548
rect -22258 -7628 -22131 -7612
rect -22258 -7692 -22211 -7628
rect -22147 -7692 -22131 -7628
rect -22258 -7708 -22131 -7692
rect -22258 -7772 -22211 -7708
rect -22147 -7772 -22131 -7708
rect -22258 -7788 -22131 -7772
rect -22258 -7852 -22211 -7788
rect -22147 -7852 -22131 -7788
rect -22258 -7868 -22131 -7852
rect -22258 -7932 -22211 -7868
rect -22147 -7932 -22131 -7868
rect -22258 -7948 -22131 -7932
rect -22258 -8012 -22211 -7948
rect -22147 -8012 -22131 -7948
rect -22258 -8028 -22131 -8012
rect -22258 -8092 -22211 -8028
rect -22147 -8092 -22131 -8028
rect -22258 -8108 -22131 -8092
rect -22258 -8172 -22211 -8108
rect -22147 -8172 -22131 -8108
rect -22258 -8188 -22131 -8172
rect -22258 -8252 -22211 -8188
rect -22147 -8252 -22131 -8188
rect -22258 -8268 -22131 -8252
rect -22258 -8332 -22211 -8268
rect -22147 -8332 -22131 -8268
rect -22258 -8348 -22131 -8332
rect -22258 -8412 -22211 -8348
rect -22147 -8412 -22131 -8348
rect -22258 -8428 -22131 -8412
rect -22258 -8492 -22211 -8428
rect -22147 -8492 -22131 -8428
rect -22258 -8508 -22131 -8492
rect -22258 -8572 -22211 -8508
rect -22147 -8572 -22131 -8508
rect -22258 -8588 -22131 -8572
rect -22258 -8652 -22211 -8588
rect -22147 -8652 -22131 -8588
rect -22258 -8668 -22131 -8652
rect -22258 -8732 -22211 -8668
rect -22147 -8732 -22131 -8668
rect -22258 -8748 -22131 -8732
rect -22258 -8812 -22211 -8748
rect -22147 -8812 -22131 -8748
rect -22258 -8828 -22131 -8812
rect -22258 -8892 -22211 -8828
rect -22147 -8892 -22131 -8828
rect -22258 -8908 -22131 -8892
rect -22258 -8972 -22211 -8908
rect -22147 -8972 -22131 -8908
rect -22258 -8988 -22131 -8972
rect -22258 -9052 -22211 -8988
rect -22147 -9052 -22131 -8988
rect -22258 -9068 -22131 -9052
rect -22258 -9132 -22211 -9068
rect -22147 -9132 -22131 -9068
rect -22258 -9148 -22131 -9132
rect -22258 -9212 -22211 -9148
rect -22147 -9212 -22131 -9148
rect -22258 -9228 -22131 -9212
rect -28577 -9308 -28450 -9292
rect -28577 -9372 -28530 -9308
rect -28466 -9372 -28450 -9308
rect -28577 -9388 -28450 -9372
rect -28577 -9512 -28473 -9388
rect -28577 -9528 -28450 -9512
rect -28577 -9592 -28530 -9528
rect -28466 -9592 -28450 -9528
rect -28577 -9608 -28450 -9592
rect -34896 -9688 -34769 -9672
rect -34896 -9752 -34849 -9688
rect -34785 -9752 -34769 -9688
rect -34896 -9768 -34769 -9752
rect -34896 -9832 -34849 -9768
rect -34785 -9832 -34769 -9768
rect -34896 -9848 -34769 -9832
rect -34896 -9912 -34849 -9848
rect -34785 -9912 -34769 -9848
rect -34896 -9928 -34769 -9912
rect -34896 -9992 -34849 -9928
rect -34785 -9992 -34769 -9928
rect -34896 -10008 -34769 -9992
rect -34896 -10072 -34849 -10008
rect -34785 -10072 -34769 -10008
rect -34896 -10088 -34769 -10072
rect -34896 -10152 -34849 -10088
rect -34785 -10152 -34769 -10088
rect -34896 -10168 -34769 -10152
rect -34896 -10232 -34849 -10168
rect -34785 -10232 -34769 -10168
rect -34896 -10248 -34769 -10232
rect -34896 -10312 -34849 -10248
rect -34785 -10312 -34769 -10248
rect -34896 -10328 -34769 -10312
rect -34896 -10392 -34849 -10328
rect -34785 -10392 -34769 -10328
rect -34896 -10408 -34769 -10392
rect -34896 -10472 -34849 -10408
rect -34785 -10472 -34769 -10408
rect -34896 -10488 -34769 -10472
rect -34896 -10552 -34849 -10488
rect -34785 -10552 -34769 -10488
rect -34896 -10568 -34769 -10552
rect -34896 -10632 -34849 -10568
rect -34785 -10632 -34769 -10568
rect -34896 -10648 -34769 -10632
rect -34896 -10712 -34849 -10648
rect -34785 -10712 -34769 -10648
rect -34896 -10728 -34769 -10712
rect -34896 -10792 -34849 -10728
rect -34785 -10792 -34769 -10728
rect -34896 -10808 -34769 -10792
rect -34896 -10872 -34849 -10808
rect -34785 -10872 -34769 -10808
rect -34896 -10888 -34769 -10872
rect -34896 -10952 -34849 -10888
rect -34785 -10952 -34769 -10888
rect -34896 -10968 -34769 -10952
rect -34896 -11032 -34849 -10968
rect -34785 -11032 -34769 -10968
rect -34896 -11048 -34769 -11032
rect -34896 -11112 -34849 -11048
rect -34785 -11112 -34769 -11048
rect -34896 -11128 -34769 -11112
rect -34896 -11192 -34849 -11128
rect -34785 -11192 -34769 -11128
rect -34896 -11208 -34769 -11192
rect -34896 -11272 -34849 -11208
rect -34785 -11272 -34769 -11208
rect -34896 -11288 -34769 -11272
rect -34896 -11352 -34849 -11288
rect -34785 -11352 -34769 -11288
rect -34896 -11368 -34769 -11352
rect -34896 -11432 -34849 -11368
rect -34785 -11432 -34769 -11368
rect -34896 -11448 -34769 -11432
rect -34896 -11512 -34849 -11448
rect -34785 -11512 -34769 -11448
rect -34896 -11528 -34769 -11512
rect -34896 -11592 -34849 -11528
rect -34785 -11592 -34769 -11528
rect -34896 -11608 -34769 -11592
rect -34896 -11672 -34849 -11608
rect -34785 -11672 -34769 -11608
rect -34896 -11688 -34769 -11672
rect -34896 -11752 -34849 -11688
rect -34785 -11752 -34769 -11688
rect -34896 -11768 -34769 -11752
rect -34896 -11832 -34849 -11768
rect -34785 -11832 -34769 -11768
rect -34896 -11848 -34769 -11832
rect -34896 -11912 -34849 -11848
rect -34785 -11912 -34769 -11848
rect -34896 -11928 -34769 -11912
rect -34896 -11992 -34849 -11928
rect -34785 -11992 -34769 -11928
rect -34896 -12008 -34769 -11992
rect -34896 -12072 -34849 -12008
rect -34785 -12072 -34769 -12008
rect -34896 -12088 -34769 -12072
rect -34896 -12152 -34849 -12088
rect -34785 -12152 -34769 -12088
rect -34896 -12168 -34769 -12152
rect -34896 -12232 -34849 -12168
rect -34785 -12232 -34769 -12168
rect -34896 -12248 -34769 -12232
rect -34896 -12312 -34849 -12248
rect -34785 -12312 -34769 -12248
rect -34896 -12328 -34769 -12312
rect -34896 -12392 -34849 -12328
rect -34785 -12392 -34769 -12328
rect -34896 -12408 -34769 -12392
rect -34896 -12472 -34849 -12408
rect -34785 -12472 -34769 -12408
rect -34896 -12488 -34769 -12472
rect -34896 -12552 -34849 -12488
rect -34785 -12552 -34769 -12488
rect -34896 -12568 -34769 -12552
rect -34896 -12632 -34849 -12568
rect -34785 -12632 -34769 -12568
rect -34896 -12648 -34769 -12632
rect -34896 -12712 -34849 -12648
rect -34785 -12712 -34769 -12648
rect -34896 -12728 -34769 -12712
rect -34896 -12792 -34849 -12728
rect -34785 -12792 -34769 -12728
rect -34896 -12808 -34769 -12792
rect -34896 -12872 -34849 -12808
rect -34785 -12872 -34769 -12808
rect -34896 -12888 -34769 -12872
rect -34896 -12952 -34849 -12888
rect -34785 -12952 -34769 -12888
rect -34896 -12968 -34769 -12952
rect -34896 -13032 -34849 -12968
rect -34785 -13032 -34769 -12968
rect -34896 -13048 -34769 -13032
rect -34896 -13112 -34849 -13048
rect -34785 -13112 -34769 -13048
rect -34896 -13128 -34769 -13112
rect -34896 -13192 -34849 -13128
rect -34785 -13192 -34769 -13128
rect -34896 -13208 -34769 -13192
rect -34896 -13272 -34849 -13208
rect -34785 -13272 -34769 -13208
rect -34896 -13288 -34769 -13272
rect -34896 -13352 -34849 -13288
rect -34785 -13352 -34769 -13288
rect -34896 -13368 -34769 -13352
rect -34896 -13432 -34849 -13368
rect -34785 -13432 -34769 -13368
rect -34896 -13448 -34769 -13432
rect -34896 -13512 -34849 -13448
rect -34785 -13512 -34769 -13448
rect -34896 -13528 -34769 -13512
rect -34896 -13592 -34849 -13528
rect -34785 -13592 -34769 -13528
rect -34896 -13608 -34769 -13592
rect -34896 -13672 -34849 -13608
rect -34785 -13672 -34769 -13608
rect -34896 -13688 -34769 -13672
rect -34896 -13752 -34849 -13688
rect -34785 -13752 -34769 -13688
rect -34896 -13768 -34769 -13752
rect -34896 -13832 -34849 -13768
rect -34785 -13832 -34769 -13768
rect -34896 -13848 -34769 -13832
rect -34896 -13912 -34849 -13848
rect -34785 -13912 -34769 -13848
rect -34896 -13928 -34769 -13912
rect -34896 -13992 -34849 -13928
rect -34785 -13992 -34769 -13928
rect -34896 -14008 -34769 -13992
rect -34896 -14072 -34849 -14008
rect -34785 -14072 -34769 -14008
rect -34896 -14088 -34769 -14072
rect -34896 -14152 -34849 -14088
rect -34785 -14152 -34769 -14088
rect -34896 -14168 -34769 -14152
rect -34896 -14232 -34849 -14168
rect -34785 -14232 -34769 -14168
rect -34896 -14248 -34769 -14232
rect -34896 -14312 -34849 -14248
rect -34785 -14312 -34769 -14248
rect -34896 -14328 -34769 -14312
rect -34896 -14392 -34849 -14328
rect -34785 -14392 -34769 -14328
rect -34896 -14408 -34769 -14392
rect -34896 -14472 -34849 -14408
rect -34785 -14472 -34769 -14408
rect -34896 -14488 -34769 -14472
rect -34896 -14552 -34849 -14488
rect -34785 -14552 -34769 -14488
rect -34896 -14568 -34769 -14552
rect -34896 -14632 -34849 -14568
rect -34785 -14632 -34769 -14568
rect -34896 -14648 -34769 -14632
rect -34896 -14712 -34849 -14648
rect -34785 -14712 -34769 -14648
rect -34896 -14728 -34769 -14712
rect -34896 -14792 -34849 -14728
rect -34785 -14792 -34769 -14728
rect -34896 -14808 -34769 -14792
rect -34896 -14872 -34849 -14808
rect -34785 -14872 -34769 -14808
rect -34896 -14888 -34769 -14872
rect -34896 -14952 -34849 -14888
rect -34785 -14952 -34769 -14888
rect -34896 -14968 -34769 -14952
rect -34896 -15032 -34849 -14968
rect -34785 -15032 -34769 -14968
rect -34896 -15048 -34769 -15032
rect -34896 -15112 -34849 -15048
rect -34785 -15112 -34769 -15048
rect -34896 -15128 -34769 -15112
rect -34896 -15192 -34849 -15128
rect -34785 -15192 -34769 -15128
rect -34896 -15208 -34769 -15192
rect -34896 -15272 -34849 -15208
rect -34785 -15272 -34769 -15208
rect -34896 -15288 -34769 -15272
rect -34896 -15352 -34849 -15288
rect -34785 -15352 -34769 -15288
rect -34896 -15368 -34769 -15352
rect -34896 -15432 -34849 -15368
rect -34785 -15432 -34769 -15368
rect -34896 -15448 -34769 -15432
rect -34896 -15512 -34849 -15448
rect -34785 -15512 -34769 -15448
rect -34896 -15528 -34769 -15512
rect -41215 -15608 -41088 -15592
rect -41215 -15672 -41168 -15608
rect -41104 -15672 -41088 -15608
rect -41215 -15688 -41088 -15672
rect -41215 -15812 -41111 -15688
rect -41215 -15828 -41088 -15812
rect -41215 -15892 -41168 -15828
rect -41104 -15892 -41088 -15828
rect -41215 -15908 -41088 -15892
rect -47244 -15948 -41322 -15939
rect -47244 -21852 -47235 -15948
rect -41331 -21852 -41322 -15948
rect -47244 -21861 -41322 -21852
rect -41215 -15972 -41168 -15908
rect -41104 -15972 -41088 -15908
rect -38016 -15939 -37912 -15561
rect -34896 -15592 -34849 -15528
rect -34785 -15592 -34769 -15528
rect -34606 -9648 -28684 -9639
rect -34606 -15552 -34597 -9648
rect -28693 -15552 -28684 -9648
rect -34606 -15561 -28684 -15552
rect -28577 -9672 -28530 -9608
rect -28466 -9672 -28450 -9608
rect -25378 -9639 -25274 -9261
rect -22258 -9292 -22211 -9228
rect -22147 -9292 -22131 -9228
rect -21968 -3348 -16046 -3339
rect -21968 -9252 -21959 -3348
rect -16055 -9252 -16046 -3348
rect -21968 -9261 -16046 -9252
rect -15939 -3372 -15892 -3308
rect -15828 -3372 -15812 -3308
rect -12740 -3339 -12636 -2961
rect -9620 -2992 -9573 -2928
rect -9509 -2992 -9493 -2928
rect -9330 2952 -3408 2961
rect -9330 -2952 -9321 2952
rect -3417 -2952 -3408 2952
rect -9330 -2961 -3408 -2952
rect -3301 2928 -3254 2992
rect -3190 2928 -3174 2992
rect -102 2961 2 3339
rect 3018 3308 3065 3372
rect 3129 3308 3145 3372
rect 3308 9252 9230 9261
rect 3308 3348 3317 9252
rect 9221 3348 9230 9252
rect 3308 3339 9230 3348
rect 9337 9228 9384 9292
rect 9448 9228 9464 9292
rect 12536 9261 12640 9639
rect 15656 9608 15703 9672
rect 15767 9608 15783 9672
rect 15946 15552 21868 15561
rect 15946 9648 15955 15552
rect 21859 9648 21868 15552
rect 15946 9639 21868 9648
rect 21975 15528 22022 15592
rect 22086 15528 22102 15592
rect 25174 15561 25278 15939
rect 28294 15908 28341 15972
rect 28405 15908 28421 15972
rect 28584 21852 34506 21861
rect 28584 15948 28593 21852
rect 34497 15948 34506 21852
rect 28584 15939 34506 15948
rect 34613 21828 34660 21892
rect 34724 21828 34740 21892
rect 37812 21861 37916 22239
rect 40932 22208 40979 22272
rect 41043 22208 41059 22272
rect 41222 28152 47144 28161
rect 41222 22248 41231 28152
rect 47135 22248 47144 28152
rect 41222 22239 47144 22248
rect 47251 28128 47298 28192
rect 47362 28128 47378 28192
rect 47251 28112 47378 28128
rect 47251 28048 47298 28112
rect 47362 28048 47378 28112
rect 47251 28032 47378 28048
rect 47251 27968 47298 28032
rect 47362 27968 47378 28032
rect 47251 27952 47378 27968
rect 47251 27888 47298 27952
rect 47362 27888 47378 27952
rect 47251 27872 47378 27888
rect 47251 27808 47298 27872
rect 47362 27808 47378 27872
rect 47251 27792 47378 27808
rect 47251 27728 47298 27792
rect 47362 27728 47378 27792
rect 47251 27712 47378 27728
rect 47251 27648 47298 27712
rect 47362 27648 47378 27712
rect 47251 27632 47378 27648
rect 47251 27568 47298 27632
rect 47362 27568 47378 27632
rect 47251 27552 47378 27568
rect 47251 27488 47298 27552
rect 47362 27488 47378 27552
rect 47251 27472 47378 27488
rect 47251 27408 47298 27472
rect 47362 27408 47378 27472
rect 47251 27392 47378 27408
rect 47251 27328 47298 27392
rect 47362 27328 47378 27392
rect 47251 27312 47378 27328
rect 47251 27248 47298 27312
rect 47362 27248 47378 27312
rect 47251 27232 47378 27248
rect 47251 27168 47298 27232
rect 47362 27168 47378 27232
rect 47251 27152 47378 27168
rect 47251 27088 47298 27152
rect 47362 27088 47378 27152
rect 47251 27072 47378 27088
rect 47251 27008 47298 27072
rect 47362 27008 47378 27072
rect 47251 26992 47378 27008
rect 47251 26928 47298 26992
rect 47362 26928 47378 26992
rect 47251 26912 47378 26928
rect 47251 26848 47298 26912
rect 47362 26848 47378 26912
rect 47251 26832 47378 26848
rect 47251 26768 47298 26832
rect 47362 26768 47378 26832
rect 47251 26752 47378 26768
rect 47251 26688 47298 26752
rect 47362 26688 47378 26752
rect 47251 26672 47378 26688
rect 47251 26608 47298 26672
rect 47362 26608 47378 26672
rect 47251 26592 47378 26608
rect 47251 26528 47298 26592
rect 47362 26528 47378 26592
rect 47251 26512 47378 26528
rect 47251 26448 47298 26512
rect 47362 26448 47378 26512
rect 47251 26432 47378 26448
rect 47251 26368 47298 26432
rect 47362 26368 47378 26432
rect 47251 26352 47378 26368
rect 47251 26288 47298 26352
rect 47362 26288 47378 26352
rect 47251 26272 47378 26288
rect 47251 26208 47298 26272
rect 47362 26208 47378 26272
rect 47251 26192 47378 26208
rect 47251 26128 47298 26192
rect 47362 26128 47378 26192
rect 47251 26112 47378 26128
rect 47251 26048 47298 26112
rect 47362 26048 47378 26112
rect 47251 26032 47378 26048
rect 47251 25968 47298 26032
rect 47362 25968 47378 26032
rect 47251 25952 47378 25968
rect 47251 25888 47298 25952
rect 47362 25888 47378 25952
rect 47251 25872 47378 25888
rect 47251 25808 47298 25872
rect 47362 25808 47378 25872
rect 47251 25792 47378 25808
rect 47251 25728 47298 25792
rect 47362 25728 47378 25792
rect 47251 25712 47378 25728
rect 47251 25648 47298 25712
rect 47362 25648 47378 25712
rect 47251 25632 47378 25648
rect 47251 25568 47298 25632
rect 47362 25568 47378 25632
rect 47251 25552 47378 25568
rect 47251 25488 47298 25552
rect 47362 25488 47378 25552
rect 47251 25472 47378 25488
rect 47251 25408 47298 25472
rect 47362 25408 47378 25472
rect 47251 25392 47378 25408
rect 47251 25328 47298 25392
rect 47362 25328 47378 25392
rect 47251 25312 47378 25328
rect 47251 25248 47298 25312
rect 47362 25248 47378 25312
rect 47251 25232 47378 25248
rect 47251 25168 47298 25232
rect 47362 25168 47378 25232
rect 47251 25152 47378 25168
rect 47251 25088 47298 25152
rect 47362 25088 47378 25152
rect 47251 25072 47378 25088
rect 47251 25008 47298 25072
rect 47362 25008 47378 25072
rect 47251 24992 47378 25008
rect 47251 24928 47298 24992
rect 47362 24928 47378 24992
rect 47251 24912 47378 24928
rect 47251 24848 47298 24912
rect 47362 24848 47378 24912
rect 47251 24832 47378 24848
rect 47251 24768 47298 24832
rect 47362 24768 47378 24832
rect 47251 24752 47378 24768
rect 47251 24688 47298 24752
rect 47362 24688 47378 24752
rect 47251 24672 47378 24688
rect 47251 24608 47298 24672
rect 47362 24608 47378 24672
rect 47251 24592 47378 24608
rect 47251 24528 47298 24592
rect 47362 24528 47378 24592
rect 47251 24512 47378 24528
rect 47251 24448 47298 24512
rect 47362 24448 47378 24512
rect 47251 24432 47378 24448
rect 47251 24368 47298 24432
rect 47362 24368 47378 24432
rect 47251 24352 47378 24368
rect 47251 24288 47298 24352
rect 47362 24288 47378 24352
rect 47251 24272 47378 24288
rect 47251 24208 47298 24272
rect 47362 24208 47378 24272
rect 47251 24192 47378 24208
rect 47251 24128 47298 24192
rect 47362 24128 47378 24192
rect 47251 24112 47378 24128
rect 47251 24048 47298 24112
rect 47362 24048 47378 24112
rect 47251 24032 47378 24048
rect 47251 23968 47298 24032
rect 47362 23968 47378 24032
rect 47251 23952 47378 23968
rect 47251 23888 47298 23952
rect 47362 23888 47378 23952
rect 47251 23872 47378 23888
rect 47251 23808 47298 23872
rect 47362 23808 47378 23872
rect 47251 23792 47378 23808
rect 47251 23728 47298 23792
rect 47362 23728 47378 23792
rect 47251 23712 47378 23728
rect 47251 23648 47298 23712
rect 47362 23648 47378 23712
rect 47251 23632 47378 23648
rect 47251 23568 47298 23632
rect 47362 23568 47378 23632
rect 47251 23552 47378 23568
rect 47251 23488 47298 23552
rect 47362 23488 47378 23552
rect 47251 23472 47378 23488
rect 47251 23408 47298 23472
rect 47362 23408 47378 23472
rect 47251 23392 47378 23408
rect 47251 23328 47298 23392
rect 47362 23328 47378 23392
rect 47251 23312 47378 23328
rect 47251 23248 47298 23312
rect 47362 23248 47378 23312
rect 47251 23232 47378 23248
rect 47251 23168 47298 23232
rect 47362 23168 47378 23232
rect 47251 23152 47378 23168
rect 47251 23088 47298 23152
rect 47362 23088 47378 23152
rect 47251 23072 47378 23088
rect 47251 23008 47298 23072
rect 47362 23008 47378 23072
rect 47251 22992 47378 23008
rect 47251 22928 47298 22992
rect 47362 22928 47378 22992
rect 47251 22912 47378 22928
rect 47251 22848 47298 22912
rect 47362 22848 47378 22912
rect 47251 22832 47378 22848
rect 47251 22768 47298 22832
rect 47362 22768 47378 22832
rect 47251 22752 47378 22768
rect 47251 22688 47298 22752
rect 47362 22688 47378 22752
rect 47251 22672 47378 22688
rect 47251 22608 47298 22672
rect 47362 22608 47378 22672
rect 47251 22592 47378 22608
rect 47251 22528 47298 22592
rect 47362 22528 47378 22592
rect 47251 22512 47378 22528
rect 47251 22448 47298 22512
rect 47362 22448 47378 22512
rect 47251 22432 47378 22448
rect 47251 22368 47298 22432
rect 47362 22368 47378 22432
rect 47251 22352 47378 22368
rect 47251 22288 47298 22352
rect 47362 22288 47378 22352
rect 47251 22272 47378 22288
rect 40932 22192 41059 22208
rect 40932 22128 40979 22192
rect 41043 22128 41059 22192
rect 40932 22112 41059 22128
rect 40932 21988 41036 22112
rect 40932 21972 41059 21988
rect 40932 21908 40979 21972
rect 41043 21908 41059 21972
rect 40932 21892 41059 21908
rect 34613 21812 34740 21828
rect 34613 21748 34660 21812
rect 34724 21748 34740 21812
rect 34613 21732 34740 21748
rect 34613 21668 34660 21732
rect 34724 21668 34740 21732
rect 34613 21652 34740 21668
rect 34613 21588 34660 21652
rect 34724 21588 34740 21652
rect 34613 21572 34740 21588
rect 34613 21508 34660 21572
rect 34724 21508 34740 21572
rect 34613 21492 34740 21508
rect 34613 21428 34660 21492
rect 34724 21428 34740 21492
rect 34613 21412 34740 21428
rect 34613 21348 34660 21412
rect 34724 21348 34740 21412
rect 34613 21332 34740 21348
rect 34613 21268 34660 21332
rect 34724 21268 34740 21332
rect 34613 21252 34740 21268
rect 34613 21188 34660 21252
rect 34724 21188 34740 21252
rect 34613 21172 34740 21188
rect 34613 21108 34660 21172
rect 34724 21108 34740 21172
rect 34613 21092 34740 21108
rect 34613 21028 34660 21092
rect 34724 21028 34740 21092
rect 34613 21012 34740 21028
rect 34613 20948 34660 21012
rect 34724 20948 34740 21012
rect 34613 20932 34740 20948
rect 34613 20868 34660 20932
rect 34724 20868 34740 20932
rect 34613 20852 34740 20868
rect 34613 20788 34660 20852
rect 34724 20788 34740 20852
rect 34613 20772 34740 20788
rect 34613 20708 34660 20772
rect 34724 20708 34740 20772
rect 34613 20692 34740 20708
rect 34613 20628 34660 20692
rect 34724 20628 34740 20692
rect 34613 20612 34740 20628
rect 34613 20548 34660 20612
rect 34724 20548 34740 20612
rect 34613 20532 34740 20548
rect 34613 20468 34660 20532
rect 34724 20468 34740 20532
rect 34613 20452 34740 20468
rect 34613 20388 34660 20452
rect 34724 20388 34740 20452
rect 34613 20372 34740 20388
rect 34613 20308 34660 20372
rect 34724 20308 34740 20372
rect 34613 20292 34740 20308
rect 34613 20228 34660 20292
rect 34724 20228 34740 20292
rect 34613 20212 34740 20228
rect 34613 20148 34660 20212
rect 34724 20148 34740 20212
rect 34613 20132 34740 20148
rect 34613 20068 34660 20132
rect 34724 20068 34740 20132
rect 34613 20052 34740 20068
rect 34613 19988 34660 20052
rect 34724 19988 34740 20052
rect 34613 19972 34740 19988
rect 34613 19908 34660 19972
rect 34724 19908 34740 19972
rect 34613 19892 34740 19908
rect 34613 19828 34660 19892
rect 34724 19828 34740 19892
rect 34613 19812 34740 19828
rect 34613 19748 34660 19812
rect 34724 19748 34740 19812
rect 34613 19732 34740 19748
rect 34613 19668 34660 19732
rect 34724 19668 34740 19732
rect 34613 19652 34740 19668
rect 34613 19588 34660 19652
rect 34724 19588 34740 19652
rect 34613 19572 34740 19588
rect 34613 19508 34660 19572
rect 34724 19508 34740 19572
rect 34613 19492 34740 19508
rect 34613 19428 34660 19492
rect 34724 19428 34740 19492
rect 34613 19412 34740 19428
rect 34613 19348 34660 19412
rect 34724 19348 34740 19412
rect 34613 19332 34740 19348
rect 34613 19268 34660 19332
rect 34724 19268 34740 19332
rect 34613 19252 34740 19268
rect 34613 19188 34660 19252
rect 34724 19188 34740 19252
rect 34613 19172 34740 19188
rect 34613 19108 34660 19172
rect 34724 19108 34740 19172
rect 34613 19092 34740 19108
rect 34613 19028 34660 19092
rect 34724 19028 34740 19092
rect 34613 19012 34740 19028
rect 34613 18948 34660 19012
rect 34724 18948 34740 19012
rect 34613 18932 34740 18948
rect 34613 18868 34660 18932
rect 34724 18868 34740 18932
rect 34613 18852 34740 18868
rect 34613 18788 34660 18852
rect 34724 18788 34740 18852
rect 34613 18772 34740 18788
rect 34613 18708 34660 18772
rect 34724 18708 34740 18772
rect 34613 18692 34740 18708
rect 34613 18628 34660 18692
rect 34724 18628 34740 18692
rect 34613 18612 34740 18628
rect 34613 18548 34660 18612
rect 34724 18548 34740 18612
rect 34613 18532 34740 18548
rect 34613 18468 34660 18532
rect 34724 18468 34740 18532
rect 34613 18452 34740 18468
rect 34613 18388 34660 18452
rect 34724 18388 34740 18452
rect 34613 18372 34740 18388
rect 34613 18308 34660 18372
rect 34724 18308 34740 18372
rect 34613 18292 34740 18308
rect 34613 18228 34660 18292
rect 34724 18228 34740 18292
rect 34613 18212 34740 18228
rect 34613 18148 34660 18212
rect 34724 18148 34740 18212
rect 34613 18132 34740 18148
rect 34613 18068 34660 18132
rect 34724 18068 34740 18132
rect 34613 18052 34740 18068
rect 34613 17988 34660 18052
rect 34724 17988 34740 18052
rect 34613 17972 34740 17988
rect 34613 17908 34660 17972
rect 34724 17908 34740 17972
rect 34613 17892 34740 17908
rect 34613 17828 34660 17892
rect 34724 17828 34740 17892
rect 34613 17812 34740 17828
rect 34613 17748 34660 17812
rect 34724 17748 34740 17812
rect 34613 17732 34740 17748
rect 34613 17668 34660 17732
rect 34724 17668 34740 17732
rect 34613 17652 34740 17668
rect 34613 17588 34660 17652
rect 34724 17588 34740 17652
rect 34613 17572 34740 17588
rect 34613 17508 34660 17572
rect 34724 17508 34740 17572
rect 34613 17492 34740 17508
rect 34613 17428 34660 17492
rect 34724 17428 34740 17492
rect 34613 17412 34740 17428
rect 34613 17348 34660 17412
rect 34724 17348 34740 17412
rect 34613 17332 34740 17348
rect 34613 17268 34660 17332
rect 34724 17268 34740 17332
rect 34613 17252 34740 17268
rect 34613 17188 34660 17252
rect 34724 17188 34740 17252
rect 34613 17172 34740 17188
rect 34613 17108 34660 17172
rect 34724 17108 34740 17172
rect 34613 17092 34740 17108
rect 34613 17028 34660 17092
rect 34724 17028 34740 17092
rect 34613 17012 34740 17028
rect 34613 16948 34660 17012
rect 34724 16948 34740 17012
rect 34613 16932 34740 16948
rect 34613 16868 34660 16932
rect 34724 16868 34740 16932
rect 34613 16852 34740 16868
rect 34613 16788 34660 16852
rect 34724 16788 34740 16852
rect 34613 16772 34740 16788
rect 34613 16708 34660 16772
rect 34724 16708 34740 16772
rect 34613 16692 34740 16708
rect 34613 16628 34660 16692
rect 34724 16628 34740 16692
rect 34613 16612 34740 16628
rect 34613 16548 34660 16612
rect 34724 16548 34740 16612
rect 34613 16532 34740 16548
rect 34613 16468 34660 16532
rect 34724 16468 34740 16532
rect 34613 16452 34740 16468
rect 34613 16388 34660 16452
rect 34724 16388 34740 16452
rect 34613 16372 34740 16388
rect 34613 16308 34660 16372
rect 34724 16308 34740 16372
rect 34613 16292 34740 16308
rect 34613 16228 34660 16292
rect 34724 16228 34740 16292
rect 34613 16212 34740 16228
rect 34613 16148 34660 16212
rect 34724 16148 34740 16212
rect 34613 16132 34740 16148
rect 34613 16068 34660 16132
rect 34724 16068 34740 16132
rect 34613 16052 34740 16068
rect 34613 15988 34660 16052
rect 34724 15988 34740 16052
rect 34613 15972 34740 15988
rect 28294 15892 28421 15908
rect 28294 15828 28341 15892
rect 28405 15828 28421 15892
rect 28294 15812 28421 15828
rect 28294 15688 28398 15812
rect 28294 15672 28421 15688
rect 28294 15608 28341 15672
rect 28405 15608 28421 15672
rect 28294 15592 28421 15608
rect 21975 15512 22102 15528
rect 21975 15448 22022 15512
rect 22086 15448 22102 15512
rect 21975 15432 22102 15448
rect 21975 15368 22022 15432
rect 22086 15368 22102 15432
rect 21975 15352 22102 15368
rect 21975 15288 22022 15352
rect 22086 15288 22102 15352
rect 21975 15272 22102 15288
rect 21975 15208 22022 15272
rect 22086 15208 22102 15272
rect 21975 15192 22102 15208
rect 21975 15128 22022 15192
rect 22086 15128 22102 15192
rect 21975 15112 22102 15128
rect 21975 15048 22022 15112
rect 22086 15048 22102 15112
rect 21975 15032 22102 15048
rect 21975 14968 22022 15032
rect 22086 14968 22102 15032
rect 21975 14952 22102 14968
rect 21975 14888 22022 14952
rect 22086 14888 22102 14952
rect 21975 14872 22102 14888
rect 21975 14808 22022 14872
rect 22086 14808 22102 14872
rect 21975 14792 22102 14808
rect 21975 14728 22022 14792
rect 22086 14728 22102 14792
rect 21975 14712 22102 14728
rect 21975 14648 22022 14712
rect 22086 14648 22102 14712
rect 21975 14632 22102 14648
rect 21975 14568 22022 14632
rect 22086 14568 22102 14632
rect 21975 14552 22102 14568
rect 21975 14488 22022 14552
rect 22086 14488 22102 14552
rect 21975 14472 22102 14488
rect 21975 14408 22022 14472
rect 22086 14408 22102 14472
rect 21975 14392 22102 14408
rect 21975 14328 22022 14392
rect 22086 14328 22102 14392
rect 21975 14312 22102 14328
rect 21975 14248 22022 14312
rect 22086 14248 22102 14312
rect 21975 14232 22102 14248
rect 21975 14168 22022 14232
rect 22086 14168 22102 14232
rect 21975 14152 22102 14168
rect 21975 14088 22022 14152
rect 22086 14088 22102 14152
rect 21975 14072 22102 14088
rect 21975 14008 22022 14072
rect 22086 14008 22102 14072
rect 21975 13992 22102 14008
rect 21975 13928 22022 13992
rect 22086 13928 22102 13992
rect 21975 13912 22102 13928
rect 21975 13848 22022 13912
rect 22086 13848 22102 13912
rect 21975 13832 22102 13848
rect 21975 13768 22022 13832
rect 22086 13768 22102 13832
rect 21975 13752 22102 13768
rect 21975 13688 22022 13752
rect 22086 13688 22102 13752
rect 21975 13672 22102 13688
rect 21975 13608 22022 13672
rect 22086 13608 22102 13672
rect 21975 13592 22102 13608
rect 21975 13528 22022 13592
rect 22086 13528 22102 13592
rect 21975 13512 22102 13528
rect 21975 13448 22022 13512
rect 22086 13448 22102 13512
rect 21975 13432 22102 13448
rect 21975 13368 22022 13432
rect 22086 13368 22102 13432
rect 21975 13352 22102 13368
rect 21975 13288 22022 13352
rect 22086 13288 22102 13352
rect 21975 13272 22102 13288
rect 21975 13208 22022 13272
rect 22086 13208 22102 13272
rect 21975 13192 22102 13208
rect 21975 13128 22022 13192
rect 22086 13128 22102 13192
rect 21975 13112 22102 13128
rect 21975 13048 22022 13112
rect 22086 13048 22102 13112
rect 21975 13032 22102 13048
rect 21975 12968 22022 13032
rect 22086 12968 22102 13032
rect 21975 12952 22102 12968
rect 21975 12888 22022 12952
rect 22086 12888 22102 12952
rect 21975 12872 22102 12888
rect 21975 12808 22022 12872
rect 22086 12808 22102 12872
rect 21975 12792 22102 12808
rect 21975 12728 22022 12792
rect 22086 12728 22102 12792
rect 21975 12712 22102 12728
rect 21975 12648 22022 12712
rect 22086 12648 22102 12712
rect 21975 12632 22102 12648
rect 21975 12568 22022 12632
rect 22086 12568 22102 12632
rect 21975 12552 22102 12568
rect 21975 12488 22022 12552
rect 22086 12488 22102 12552
rect 21975 12472 22102 12488
rect 21975 12408 22022 12472
rect 22086 12408 22102 12472
rect 21975 12392 22102 12408
rect 21975 12328 22022 12392
rect 22086 12328 22102 12392
rect 21975 12312 22102 12328
rect 21975 12248 22022 12312
rect 22086 12248 22102 12312
rect 21975 12232 22102 12248
rect 21975 12168 22022 12232
rect 22086 12168 22102 12232
rect 21975 12152 22102 12168
rect 21975 12088 22022 12152
rect 22086 12088 22102 12152
rect 21975 12072 22102 12088
rect 21975 12008 22022 12072
rect 22086 12008 22102 12072
rect 21975 11992 22102 12008
rect 21975 11928 22022 11992
rect 22086 11928 22102 11992
rect 21975 11912 22102 11928
rect 21975 11848 22022 11912
rect 22086 11848 22102 11912
rect 21975 11832 22102 11848
rect 21975 11768 22022 11832
rect 22086 11768 22102 11832
rect 21975 11752 22102 11768
rect 21975 11688 22022 11752
rect 22086 11688 22102 11752
rect 21975 11672 22102 11688
rect 21975 11608 22022 11672
rect 22086 11608 22102 11672
rect 21975 11592 22102 11608
rect 21975 11528 22022 11592
rect 22086 11528 22102 11592
rect 21975 11512 22102 11528
rect 21975 11448 22022 11512
rect 22086 11448 22102 11512
rect 21975 11432 22102 11448
rect 21975 11368 22022 11432
rect 22086 11368 22102 11432
rect 21975 11352 22102 11368
rect 21975 11288 22022 11352
rect 22086 11288 22102 11352
rect 21975 11272 22102 11288
rect 21975 11208 22022 11272
rect 22086 11208 22102 11272
rect 21975 11192 22102 11208
rect 21975 11128 22022 11192
rect 22086 11128 22102 11192
rect 21975 11112 22102 11128
rect 21975 11048 22022 11112
rect 22086 11048 22102 11112
rect 21975 11032 22102 11048
rect 21975 10968 22022 11032
rect 22086 10968 22102 11032
rect 21975 10952 22102 10968
rect 21975 10888 22022 10952
rect 22086 10888 22102 10952
rect 21975 10872 22102 10888
rect 21975 10808 22022 10872
rect 22086 10808 22102 10872
rect 21975 10792 22102 10808
rect 21975 10728 22022 10792
rect 22086 10728 22102 10792
rect 21975 10712 22102 10728
rect 21975 10648 22022 10712
rect 22086 10648 22102 10712
rect 21975 10632 22102 10648
rect 21975 10568 22022 10632
rect 22086 10568 22102 10632
rect 21975 10552 22102 10568
rect 21975 10488 22022 10552
rect 22086 10488 22102 10552
rect 21975 10472 22102 10488
rect 21975 10408 22022 10472
rect 22086 10408 22102 10472
rect 21975 10392 22102 10408
rect 21975 10328 22022 10392
rect 22086 10328 22102 10392
rect 21975 10312 22102 10328
rect 21975 10248 22022 10312
rect 22086 10248 22102 10312
rect 21975 10232 22102 10248
rect 21975 10168 22022 10232
rect 22086 10168 22102 10232
rect 21975 10152 22102 10168
rect 21975 10088 22022 10152
rect 22086 10088 22102 10152
rect 21975 10072 22102 10088
rect 21975 10008 22022 10072
rect 22086 10008 22102 10072
rect 21975 9992 22102 10008
rect 21975 9928 22022 9992
rect 22086 9928 22102 9992
rect 21975 9912 22102 9928
rect 21975 9848 22022 9912
rect 22086 9848 22102 9912
rect 21975 9832 22102 9848
rect 21975 9768 22022 9832
rect 22086 9768 22102 9832
rect 21975 9752 22102 9768
rect 21975 9688 22022 9752
rect 22086 9688 22102 9752
rect 21975 9672 22102 9688
rect 15656 9592 15783 9608
rect 15656 9528 15703 9592
rect 15767 9528 15783 9592
rect 15656 9512 15783 9528
rect 15656 9388 15760 9512
rect 15656 9372 15783 9388
rect 15656 9308 15703 9372
rect 15767 9308 15783 9372
rect 15656 9292 15783 9308
rect 9337 9212 9464 9228
rect 9337 9148 9384 9212
rect 9448 9148 9464 9212
rect 9337 9132 9464 9148
rect 9337 9068 9384 9132
rect 9448 9068 9464 9132
rect 9337 9052 9464 9068
rect 9337 8988 9384 9052
rect 9448 8988 9464 9052
rect 9337 8972 9464 8988
rect 9337 8908 9384 8972
rect 9448 8908 9464 8972
rect 9337 8892 9464 8908
rect 9337 8828 9384 8892
rect 9448 8828 9464 8892
rect 9337 8812 9464 8828
rect 9337 8748 9384 8812
rect 9448 8748 9464 8812
rect 9337 8732 9464 8748
rect 9337 8668 9384 8732
rect 9448 8668 9464 8732
rect 9337 8652 9464 8668
rect 9337 8588 9384 8652
rect 9448 8588 9464 8652
rect 9337 8572 9464 8588
rect 9337 8508 9384 8572
rect 9448 8508 9464 8572
rect 9337 8492 9464 8508
rect 9337 8428 9384 8492
rect 9448 8428 9464 8492
rect 9337 8412 9464 8428
rect 9337 8348 9384 8412
rect 9448 8348 9464 8412
rect 9337 8332 9464 8348
rect 9337 8268 9384 8332
rect 9448 8268 9464 8332
rect 9337 8252 9464 8268
rect 9337 8188 9384 8252
rect 9448 8188 9464 8252
rect 9337 8172 9464 8188
rect 9337 8108 9384 8172
rect 9448 8108 9464 8172
rect 9337 8092 9464 8108
rect 9337 8028 9384 8092
rect 9448 8028 9464 8092
rect 9337 8012 9464 8028
rect 9337 7948 9384 8012
rect 9448 7948 9464 8012
rect 9337 7932 9464 7948
rect 9337 7868 9384 7932
rect 9448 7868 9464 7932
rect 9337 7852 9464 7868
rect 9337 7788 9384 7852
rect 9448 7788 9464 7852
rect 9337 7772 9464 7788
rect 9337 7708 9384 7772
rect 9448 7708 9464 7772
rect 9337 7692 9464 7708
rect 9337 7628 9384 7692
rect 9448 7628 9464 7692
rect 9337 7612 9464 7628
rect 9337 7548 9384 7612
rect 9448 7548 9464 7612
rect 9337 7532 9464 7548
rect 9337 7468 9384 7532
rect 9448 7468 9464 7532
rect 9337 7452 9464 7468
rect 9337 7388 9384 7452
rect 9448 7388 9464 7452
rect 9337 7372 9464 7388
rect 9337 7308 9384 7372
rect 9448 7308 9464 7372
rect 9337 7292 9464 7308
rect 9337 7228 9384 7292
rect 9448 7228 9464 7292
rect 9337 7212 9464 7228
rect 9337 7148 9384 7212
rect 9448 7148 9464 7212
rect 9337 7132 9464 7148
rect 9337 7068 9384 7132
rect 9448 7068 9464 7132
rect 9337 7052 9464 7068
rect 9337 6988 9384 7052
rect 9448 6988 9464 7052
rect 9337 6972 9464 6988
rect 9337 6908 9384 6972
rect 9448 6908 9464 6972
rect 9337 6892 9464 6908
rect 9337 6828 9384 6892
rect 9448 6828 9464 6892
rect 9337 6812 9464 6828
rect 9337 6748 9384 6812
rect 9448 6748 9464 6812
rect 9337 6732 9464 6748
rect 9337 6668 9384 6732
rect 9448 6668 9464 6732
rect 9337 6652 9464 6668
rect 9337 6588 9384 6652
rect 9448 6588 9464 6652
rect 9337 6572 9464 6588
rect 9337 6508 9384 6572
rect 9448 6508 9464 6572
rect 9337 6492 9464 6508
rect 9337 6428 9384 6492
rect 9448 6428 9464 6492
rect 9337 6412 9464 6428
rect 9337 6348 9384 6412
rect 9448 6348 9464 6412
rect 9337 6332 9464 6348
rect 9337 6268 9384 6332
rect 9448 6268 9464 6332
rect 9337 6252 9464 6268
rect 9337 6188 9384 6252
rect 9448 6188 9464 6252
rect 9337 6172 9464 6188
rect 9337 6108 9384 6172
rect 9448 6108 9464 6172
rect 9337 6092 9464 6108
rect 9337 6028 9384 6092
rect 9448 6028 9464 6092
rect 9337 6012 9464 6028
rect 9337 5948 9384 6012
rect 9448 5948 9464 6012
rect 9337 5932 9464 5948
rect 9337 5868 9384 5932
rect 9448 5868 9464 5932
rect 9337 5852 9464 5868
rect 9337 5788 9384 5852
rect 9448 5788 9464 5852
rect 9337 5772 9464 5788
rect 9337 5708 9384 5772
rect 9448 5708 9464 5772
rect 9337 5692 9464 5708
rect 9337 5628 9384 5692
rect 9448 5628 9464 5692
rect 9337 5612 9464 5628
rect 9337 5548 9384 5612
rect 9448 5548 9464 5612
rect 9337 5532 9464 5548
rect 9337 5468 9384 5532
rect 9448 5468 9464 5532
rect 9337 5452 9464 5468
rect 9337 5388 9384 5452
rect 9448 5388 9464 5452
rect 9337 5372 9464 5388
rect 9337 5308 9384 5372
rect 9448 5308 9464 5372
rect 9337 5292 9464 5308
rect 9337 5228 9384 5292
rect 9448 5228 9464 5292
rect 9337 5212 9464 5228
rect 9337 5148 9384 5212
rect 9448 5148 9464 5212
rect 9337 5132 9464 5148
rect 9337 5068 9384 5132
rect 9448 5068 9464 5132
rect 9337 5052 9464 5068
rect 9337 4988 9384 5052
rect 9448 4988 9464 5052
rect 9337 4972 9464 4988
rect 9337 4908 9384 4972
rect 9448 4908 9464 4972
rect 9337 4892 9464 4908
rect 9337 4828 9384 4892
rect 9448 4828 9464 4892
rect 9337 4812 9464 4828
rect 9337 4748 9384 4812
rect 9448 4748 9464 4812
rect 9337 4732 9464 4748
rect 9337 4668 9384 4732
rect 9448 4668 9464 4732
rect 9337 4652 9464 4668
rect 9337 4588 9384 4652
rect 9448 4588 9464 4652
rect 9337 4572 9464 4588
rect 9337 4508 9384 4572
rect 9448 4508 9464 4572
rect 9337 4492 9464 4508
rect 9337 4428 9384 4492
rect 9448 4428 9464 4492
rect 9337 4412 9464 4428
rect 9337 4348 9384 4412
rect 9448 4348 9464 4412
rect 9337 4332 9464 4348
rect 9337 4268 9384 4332
rect 9448 4268 9464 4332
rect 9337 4252 9464 4268
rect 9337 4188 9384 4252
rect 9448 4188 9464 4252
rect 9337 4172 9464 4188
rect 9337 4108 9384 4172
rect 9448 4108 9464 4172
rect 9337 4092 9464 4108
rect 9337 4028 9384 4092
rect 9448 4028 9464 4092
rect 9337 4012 9464 4028
rect 9337 3948 9384 4012
rect 9448 3948 9464 4012
rect 9337 3932 9464 3948
rect 9337 3868 9384 3932
rect 9448 3868 9464 3932
rect 9337 3852 9464 3868
rect 9337 3788 9384 3852
rect 9448 3788 9464 3852
rect 9337 3772 9464 3788
rect 9337 3708 9384 3772
rect 9448 3708 9464 3772
rect 9337 3692 9464 3708
rect 9337 3628 9384 3692
rect 9448 3628 9464 3692
rect 9337 3612 9464 3628
rect 9337 3548 9384 3612
rect 9448 3548 9464 3612
rect 9337 3532 9464 3548
rect 9337 3468 9384 3532
rect 9448 3468 9464 3532
rect 9337 3452 9464 3468
rect 9337 3388 9384 3452
rect 9448 3388 9464 3452
rect 9337 3372 9464 3388
rect 3018 3292 3145 3308
rect 3018 3228 3065 3292
rect 3129 3228 3145 3292
rect 3018 3212 3145 3228
rect 3018 3088 3122 3212
rect 3018 3072 3145 3088
rect 3018 3008 3065 3072
rect 3129 3008 3145 3072
rect 3018 2992 3145 3008
rect -3301 2912 -3174 2928
rect -3301 2848 -3254 2912
rect -3190 2848 -3174 2912
rect -3301 2832 -3174 2848
rect -3301 2768 -3254 2832
rect -3190 2768 -3174 2832
rect -3301 2752 -3174 2768
rect -3301 2688 -3254 2752
rect -3190 2688 -3174 2752
rect -3301 2672 -3174 2688
rect -3301 2608 -3254 2672
rect -3190 2608 -3174 2672
rect -3301 2592 -3174 2608
rect -3301 2528 -3254 2592
rect -3190 2528 -3174 2592
rect -3301 2512 -3174 2528
rect -3301 2448 -3254 2512
rect -3190 2448 -3174 2512
rect -3301 2432 -3174 2448
rect -3301 2368 -3254 2432
rect -3190 2368 -3174 2432
rect -3301 2352 -3174 2368
rect -3301 2288 -3254 2352
rect -3190 2288 -3174 2352
rect -3301 2272 -3174 2288
rect -3301 2208 -3254 2272
rect -3190 2208 -3174 2272
rect -3301 2192 -3174 2208
rect -3301 2128 -3254 2192
rect -3190 2128 -3174 2192
rect -3301 2112 -3174 2128
rect -3301 2048 -3254 2112
rect -3190 2048 -3174 2112
rect -3301 2032 -3174 2048
rect -3301 1968 -3254 2032
rect -3190 1968 -3174 2032
rect -3301 1952 -3174 1968
rect -3301 1888 -3254 1952
rect -3190 1888 -3174 1952
rect -3301 1872 -3174 1888
rect -3301 1808 -3254 1872
rect -3190 1808 -3174 1872
rect -3301 1792 -3174 1808
rect -3301 1728 -3254 1792
rect -3190 1728 -3174 1792
rect -3301 1712 -3174 1728
rect -3301 1648 -3254 1712
rect -3190 1648 -3174 1712
rect -3301 1632 -3174 1648
rect -3301 1568 -3254 1632
rect -3190 1568 -3174 1632
rect -3301 1552 -3174 1568
rect -3301 1488 -3254 1552
rect -3190 1488 -3174 1552
rect -3301 1472 -3174 1488
rect -3301 1408 -3254 1472
rect -3190 1408 -3174 1472
rect -3301 1392 -3174 1408
rect -3301 1328 -3254 1392
rect -3190 1328 -3174 1392
rect -3301 1312 -3174 1328
rect -3301 1248 -3254 1312
rect -3190 1248 -3174 1312
rect -3301 1232 -3174 1248
rect -3301 1168 -3254 1232
rect -3190 1168 -3174 1232
rect -3301 1152 -3174 1168
rect -3301 1088 -3254 1152
rect -3190 1088 -3174 1152
rect -3301 1072 -3174 1088
rect -3301 1008 -3254 1072
rect -3190 1008 -3174 1072
rect -3301 992 -3174 1008
rect -3301 928 -3254 992
rect -3190 928 -3174 992
rect -3301 912 -3174 928
rect -3301 848 -3254 912
rect -3190 848 -3174 912
rect -3301 832 -3174 848
rect -3301 768 -3254 832
rect -3190 768 -3174 832
rect -3301 752 -3174 768
rect -3301 688 -3254 752
rect -3190 688 -3174 752
rect -3301 672 -3174 688
rect -3301 608 -3254 672
rect -3190 608 -3174 672
rect -3301 592 -3174 608
rect -3301 528 -3254 592
rect -3190 528 -3174 592
rect -3301 512 -3174 528
rect -3301 448 -3254 512
rect -3190 448 -3174 512
rect -3301 432 -3174 448
rect -3301 368 -3254 432
rect -3190 368 -3174 432
rect -3301 352 -3174 368
rect -3301 288 -3254 352
rect -3190 288 -3174 352
rect -3301 272 -3174 288
rect -3301 208 -3254 272
rect -3190 208 -3174 272
rect -3301 192 -3174 208
rect -3301 128 -3254 192
rect -3190 128 -3174 192
rect -3301 112 -3174 128
rect -3301 48 -3254 112
rect -3190 48 -3174 112
rect -3301 32 -3174 48
rect -3301 -32 -3254 32
rect -3190 -32 -3174 32
rect -3301 -48 -3174 -32
rect -3301 -112 -3254 -48
rect -3190 -112 -3174 -48
rect -3301 -128 -3174 -112
rect -3301 -192 -3254 -128
rect -3190 -192 -3174 -128
rect -3301 -208 -3174 -192
rect -3301 -272 -3254 -208
rect -3190 -272 -3174 -208
rect -3301 -288 -3174 -272
rect -3301 -352 -3254 -288
rect -3190 -352 -3174 -288
rect -3301 -368 -3174 -352
rect -3301 -432 -3254 -368
rect -3190 -432 -3174 -368
rect -3301 -448 -3174 -432
rect -3301 -512 -3254 -448
rect -3190 -512 -3174 -448
rect -3301 -528 -3174 -512
rect -3301 -592 -3254 -528
rect -3190 -592 -3174 -528
rect -3301 -608 -3174 -592
rect -3301 -672 -3254 -608
rect -3190 -672 -3174 -608
rect -3301 -688 -3174 -672
rect -3301 -752 -3254 -688
rect -3190 -752 -3174 -688
rect -3301 -768 -3174 -752
rect -3301 -832 -3254 -768
rect -3190 -832 -3174 -768
rect -3301 -848 -3174 -832
rect -3301 -912 -3254 -848
rect -3190 -912 -3174 -848
rect -3301 -928 -3174 -912
rect -3301 -992 -3254 -928
rect -3190 -992 -3174 -928
rect -3301 -1008 -3174 -992
rect -3301 -1072 -3254 -1008
rect -3190 -1072 -3174 -1008
rect -3301 -1088 -3174 -1072
rect -3301 -1152 -3254 -1088
rect -3190 -1152 -3174 -1088
rect -3301 -1168 -3174 -1152
rect -3301 -1232 -3254 -1168
rect -3190 -1232 -3174 -1168
rect -3301 -1248 -3174 -1232
rect -3301 -1312 -3254 -1248
rect -3190 -1312 -3174 -1248
rect -3301 -1328 -3174 -1312
rect -3301 -1392 -3254 -1328
rect -3190 -1392 -3174 -1328
rect -3301 -1408 -3174 -1392
rect -3301 -1472 -3254 -1408
rect -3190 -1472 -3174 -1408
rect -3301 -1488 -3174 -1472
rect -3301 -1552 -3254 -1488
rect -3190 -1552 -3174 -1488
rect -3301 -1568 -3174 -1552
rect -3301 -1632 -3254 -1568
rect -3190 -1632 -3174 -1568
rect -3301 -1648 -3174 -1632
rect -3301 -1712 -3254 -1648
rect -3190 -1712 -3174 -1648
rect -3301 -1728 -3174 -1712
rect -3301 -1792 -3254 -1728
rect -3190 -1792 -3174 -1728
rect -3301 -1808 -3174 -1792
rect -3301 -1872 -3254 -1808
rect -3190 -1872 -3174 -1808
rect -3301 -1888 -3174 -1872
rect -3301 -1952 -3254 -1888
rect -3190 -1952 -3174 -1888
rect -3301 -1968 -3174 -1952
rect -3301 -2032 -3254 -1968
rect -3190 -2032 -3174 -1968
rect -3301 -2048 -3174 -2032
rect -3301 -2112 -3254 -2048
rect -3190 -2112 -3174 -2048
rect -3301 -2128 -3174 -2112
rect -3301 -2192 -3254 -2128
rect -3190 -2192 -3174 -2128
rect -3301 -2208 -3174 -2192
rect -3301 -2272 -3254 -2208
rect -3190 -2272 -3174 -2208
rect -3301 -2288 -3174 -2272
rect -3301 -2352 -3254 -2288
rect -3190 -2352 -3174 -2288
rect -3301 -2368 -3174 -2352
rect -3301 -2432 -3254 -2368
rect -3190 -2432 -3174 -2368
rect -3301 -2448 -3174 -2432
rect -3301 -2512 -3254 -2448
rect -3190 -2512 -3174 -2448
rect -3301 -2528 -3174 -2512
rect -3301 -2592 -3254 -2528
rect -3190 -2592 -3174 -2528
rect -3301 -2608 -3174 -2592
rect -3301 -2672 -3254 -2608
rect -3190 -2672 -3174 -2608
rect -3301 -2688 -3174 -2672
rect -3301 -2752 -3254 -2688
rect -3190 -2752 -3174 -2688
rect -3301 -2768 -3174 -2752
rect -3301 -2832 -3254 -2768
rect -3190 -2832 -3174 -2768
rect -3301 -2848 -3174 -2832
rect -3301 -2912 -3254 -2848
rect -3190 -2912 -3174 -2848
rect -3301 -2928 -3174 -2912
rect -9620 -3008 -9493 -2992
rect -9620 -3072 -9573 -3008
rect -9509 -3072 -9493 -3008
rect -9620 -3088 -9493 -3072
rect -9620 -3212 -9516 -3088
rect -9620 -3228 -9493 -3212
rect -9620 -3292 -9573 -3228
rect -9509 -3292 -9493 -3228
rect -9620 -3308 -9493 -3292
rect -15939 -3388 -15812 -3372
rect -15939 -3452 -15892 -3388
rect -15828 -3452 -15812 -3388
rect -15939 -3468 -15812 -3452
rect -15939 -3532 -15892 -3468
rect -15828 -3532 -15812 -3468
rect -15939 -3548 -15812 -3532
rect -15939 -3612 -15892 -3548
rect -15828 -3612 -15812 -3548
rect -15939 -3628 -15812 -3612
rect -15939 -3692 -15892 -3628
rect -15828 -3692 -15812 -3628
rect -15939 -3708 -15812 -3692
rect -15939 -3772 -15892 -3708
rect -15828 -3772 -15812 -3708
rect -15939 -3788 -15812 -3772
rect -15939 -3852 -15892 -3788
rect -15828 -3852 -15812 -3788
rect -15939 -3868 -15812 -3852
rect -15939 -3932 -15892 -3868
rect -15828 -3932 -15812 -3868
rect -15939 -3948 -15812 -3932
rect -15939 -4012 -15892 -3948
rect -15828 -4012 -15812 -3948
rect -15939 -4028 -15812 -4012
rect -15939 -4092 -15892 -4028
rect -15828 -4092 -15812 -4028
rect -15939 -4108 -15812 -4092
rect -15939 -4172 -15892 -4108
rect -15828 -4172 -15812 -4108
rect -15939 -4188 -15812 -4172
rect -15939 -4252 -15892 -4188
rect -15828 -4252 -15812 -4188
rect -15939 -4268 -15812 -4252
rect -15939 -4332 -15892 -4268
rect -15828 -4332 -15812 -4268
rect -15939 -4348 -15812 -4332
rect -15939 -4412 -15892 -4348
rect -15828 -4412 -15812 -4348
rect -15939 -4428 -15812 -4412
rect -15939 -4492 -15892 -4428
rect -15828 -4492 -15812 -4428
rect -15939 -4508 -15812 -4492
rect -15939 -4572 -15892 -4508
rect -15828 -4572 -15812 -4508
rect -15939 -4588 -15812 -4572
rect -15939 -4652 -15892 -4588
rect -15828 -4652 -15812 -4588
rect -15939 -4668 -15812 -4652
rect -15939 -4732 -15892 -4668
rect -15828 -4732 -15812 -4668
rect -15939 -4748 -15812 -4732
rect -15939 -4812 -15892 -4748
rect -15828 -4812 -15812 -4748
rect -15939 -4828 -15812 -4812
rect -15939 -4892 -15892 -4828
rect -15828 -4892 -15812 -4828
rect -15939 -4908 -15812 -4892
rect -15939 -4972 -15892 -4908
rect -15828 -4972 -15812 -4908
rect -15939 -4988 -15812 -4972
rect -15939 -5052 -15892 -4988
rect -15828 -5052 -15812 -4988
rect -15939 -5068 -15812 -5052
rect -15939 -5132 -15892 -5068
rect -15828 -5132 -15812 -5068
rect -15939 -5148 -15812 -5132
rect -15939 -5212 -15892 -5148
rect -15828 -5212 -15812 -5148
rect -15939 -5228 -15812 -5212
rect -15939 -5292 -15892 -5228
rect -15828 -5292 -15812 -5228
rect -15939 -5308 -15812 -5292
rect -15939 -5372 -15892 -5308
rect -15828 -5372 -15812 -5308
rect -15939 -5388 -15812 -5372
rect -15939 -5452 -15892 -5388
rect -15828 -5452 -15812 -5388
rect -15939 -5468 -15812 -5452
rect -15939 -5532 -15892 -5468
rect -15828 -5532 -15812 -5468
rect -15939 -5548 -15812 -5532
rect -15939 -5612 -15892 -5548
rect -15828 -5612 -15812 -5548
rect -15939 -5628 -15812 -5612
rect -15939 -5692 -15892 -5628
rect -15828 -5692 -15812 -5628
rect -15939 -5708 -15812 -5692
rect -15939 -5772 -15892 -5708
rect -15828 -5772 -15812 -5708
rect -15939 -5788 -15812 -5772
rect -15939 -5852 -15892 -5788
rect -15828 -5852 -15812 -5788
rect -15939 -5868 -15812 -5852
rect -15939 -5932 -15892 -5868
rect -15828 -5932 -15812 -5868
rect -15939 -5948 -15812 -5932
rect -15939 -6012 -15892 -5948
rect -15828 -6012 -15812 -5948
rect -15939 -6028 -15812 -6012
rect -15939 -6092 -15892 -6028
rect -15828 -6092 -15812 -6028
rect -15939 -6108 -15812 -6092
rect -15939 -6172 -15892 -6108
rect -15828 -6172 -15812 -6108
rect -15939 -6188 -15812 -6172
rect -15939 -6252 -15892 -6188
rect -15828 -6252 -15812 -6188
rect -15939 -6268 -15812 -6252
rect -15939 -6332 -15892 -6268
rect -15828 -6332 -15812 -6268
rect -15939 -6348 -15812 -6332
rect -15939 -6412 -15892 -6348
rect -15828 -6412 -15812 -6348
rect -15939 -6428 -15812 -6412
rect -15939 -6492 -15892 -6428
rect -15828 -6492 -15812 -6428
rect -15939 -6508 -15812 -6492
rect -15939 -6572 -15892 -6508
rect -15828 -6572 -15812 -6508
rect -15939 -6588 -15812 -6572
rect -15939 -6652 -15892 -6588
rect -15828 -6652 -15812 -6588
rect -15939 -6668 -15812 -6652
rect -15939 -6732 -15892 -6668
rect -15828 -6732 -15812 -6668
rect -15939 -6748 -15812 -6732
rect -15939 -6812 -15892 -6748
rect -15828 -6812 -15812 -6748
rect -15939 -6828 -15812 -6812
rect -15939 -6892 -15892 -6828
rect -15828 -6892 -15812 -6828
rect -15939 -6908 -15812 -6892
rect -15939 -6972 -15892 -6908
rect -15828 -6972 -15812 -6908
rect -15939 -6988 -15812 -6972
rect -15939 -7052 -15892 -6988
rect -15828 -7052 -15812 -6988
rect -15939 -7068 -15812 -7052
rect -15939 -7132 -15892 -7068
rect -15828 -7132 -15812 -7068
rect -15939 -7148 -15812 -7132
rect -15939 -7212 -15892 -7148
rect -15828 -7212 -15812 -7148
rect -15939 -7228 -15812 -7212
rect -15939 -7292 -15892 -7228
rect -15828 -7292 -15812 -7228
rect -15939 -7308 -15812 -7292
rect -15939 -7372 -15892 -7308
rect -15828 -7372 -15812 -7308
rect -15939 -7388 -15812 -7372
rect -15939 -7452 -15892 -7388
rect -15828 -7452 -15812 -7388
rect -15939 -7468 -15812 -7452
rect -15939 -7532 -15892 -7468
rect -15828 -7532 -15812 -7468
rect -15939 -7548 -15812 -7532
rect -15939 -7612 -15892 -7548
rect -15828 -7612 -15812 -7548
rect -15939 -7628 -15812 -7612
rect -15939 -7692 -15892 -7628
rect -15828 -7692 -15812 -7628
rect -15939 -7708 -15812 -7692
rect -15939 -7772 -15892 -7708
rect -15828 -7772 -15812 -7708
rect -15939 -7788 -15812 -7772
rect -15939 -7852 -15892 -7788
rect -15828 -7852 -15812 -7788
rect -15939 -7868 -15812 -7852
rect -15939 -7932 -15892 -7868
rect -15828 -7932 -15812 -7868
rect -15939 -7948 -15812 -7932
rect -15939 -8012 -15892 -7948
rect -15828 -8012 -15812 -7948
rect -15939 -8028 -15812 -8012
rect -15939 -8092 -15892 -8028
rect -15828 -8092 -15812 -8028
rect -15939 -8108 -15812 -8092
rect -15939 -8172 -15892 -8108
rect -15828 -8172 -15812 -8108
rect -15939 -8188 -15812 -8172
rect -15939 -8252 -15892 -8188
rect -15828 -8252 -15812 -8188
rect -15939 -8268 -15812 -8252
rect -15939 -8332 -15892 -8268
rect -15828 -8332 -15812 -8268
rect -15939 -8348 -15812 -8332
rect -15939 -8412 -15892 -8348
rect -15828 -8412 -15812 -8348
rect -15939 -8428 -15812 -8412
rect -15939 -8492 -15892 -8428
rect -15828 -8492 -15812 -8428
rect -15939 -8508 -15812 -8492
rect -15939 -8572 -15892 -8508
rect -15828 -8572 -15812 -8508
rect -15939 -8588 -15812 -8572
rect -15939 -8652 -15892 -8588
rect -15828 -8652 -15812 -8588
rect -15939 -8668 -15812 -8652
rect -15939 -8732 -15892 -8668
rect -15828 -8732 -15812 -8668
rect -15939 -8748 -15812 -8732
rect -15939 -8812 -15892 -8748
rect -15828 -8812 -15812 -8748
rect -15939 -8828 -15812 -8812
rect -15939 -8892 -15892 -8828
rect -15828 -8892 -15812 -8828
rect -15939 -8908 -15812 -8892
rect -15939 -8972 -15892 -8908
rect -15828 -8972 -15812 -8908
rect -15939 -8988 -15812 -8972
rect -15939 -9052 -15892 -8988
rect -15828 -9052 -15812 -8988
rect -15939 -9068 -15812 -9052
rect -15939 -9132 -15892 -9068
rect -15828 -9132 -15812 -9068
rect -15939 -9148 -15812 -9132
rect -15939 -9212 -15892 -9148
rect -15828 -9212 -15812 -9148
rect -15939 -9228 -15812 -9212
rect -22258 -9308 -22131 -9292
rect -22258 -9372 -22211 -9308
rect -22147 -9372 -22131 -9308
rect -22258 -9388 -22131 -9372
rect -22258 -9512 -22154 -9388
rect -22258 -9528 -22131 -9512
rect -22258 -9592 -22211 -9528
rect -22147 -9592 -22131 -9528
rect -22258 -9608 -22131 -9592
rect -28577 -9688 -28450 -9672
rect -28577 -9752 -28530 -9688
rect -28466 -9752 -28450 -9688
rect -28577 -9768 -28450 -9752
rect -28577 -9832 -28530 -9768
rect -28466 -9832 -28450 -9768
rect -28577 -9848 -28450 -9832
rect -28577 -9912 -28530 -9848
rect -28466 -9912 -28450 -9848
rect -28577 -9928 -28450 -9912
rect -28577 -9992 -28530 -9928
rect -28466 -9992 -28450 -9928
rect -28577 -10008 -28450 -9992
rect -28577 -10072 -28530 -10008
rect -28466 -10072 -28450 -10008
rect -28577 -10088 -28450 -10072
rect -28577 -10152 -28530 -10088
rect -28466 -10152 -28450 -10088
rect -28577 -10168 -28450 -10152
rect -28577 -10232 -28530 -10168
rect -28466 -10232 -28450 -10168
rect -28577 -10248 -28450 -10232
rect -28577 -10312 -28530 -10248
rect -28466 -10312 -28450 -10248
rect -28577 -10328 -28450 -10312
rect -28577 -10392 -28530 -10328
rect -28466 -10392 -28450 -10328
rect -28577 -10408 -28450 -10392
rect -28577 -10472 -28530 -10408
rect -28466 -10472 -28450 -10408
rect -28577 -10488 -28450 -10472
rect -28577 -10552 -28530 -10488
rect -28466 -10552 -28450 -10488
rect -28577 -10568 -28450 -10552
rect -28577 -10632 -28530 -10568
rect -28466 -10632 -28450 -10568
rect -28577 -10648 -28450 -10632
rect -28577 -10712 -28530 -10648
rect -28466 -10712 -28450 -10648
rect -28577 -10728 -28450 -10712
rect -28577 -10792 -28530 -10728
rect -28466 -10792 -28450 -10728
rect -28577 -10808 -28450 -10792
rect -28577 -10872 -28530 -10808
rect -28466 -10872 -28450 -10808
rect -28577 -10888 -28450 -10872
rect -28577 -10952 -28530 -10888
rect -28466 -10952 -28450 -10888
rect -28577 -10968 -28450 -10952
rect -28577 -11032 -28530 -10968
rect -28466 -11032 -28450 -10968
rect -28577 -11048 -28450 -11032
rect -28577 -11112 -28530 -11048
rect -28466 -11112 -28450 -11048
rect -28577 -11128 -28450 -11112
rect -28577 -11192 -28530 -11128
rect -28466 -11192 -28450 -11128
rect -28577 -11208 -28450 -11192
rect -28577 -11272 -28530 -11208
rect -28466 -11272 -28450 -11208
rect -28577 -11288 -28450 -11272
rect -28577 -11352 -28530 -11288
rect -28466 -11352 -28450 -11288
rect -28577 -11368 -28450 -11352
rect -28577 -11432 -28530 -11368
rect -28466 -11432 -28450 -11368
rect -28577 -11448 -28450 -11432
rect -28577 -11512 -28530 -11448
rect -28466 -11512 -28450 -11448
rect -28577 -11528 -28450 -11512
rect -28577 -11592 -28530 -11528
rect -28466 -11592 -28450 -11528
rect -28577 -11608 -28450 -11592
rect -28577 -11672 -28530 -11608
rect -28466 -11672 -28450 -11608
rect -28577 -11688 -28450 -11672
rect -28577 -11752 -28530 -11688
rect -28466 -11752 -28450 -11688
rect -28577 -11768 -28450 -11752
rect -28577 -11832 -28530 -11768
rect -28466 -11832 -28450 -11768
rect -28577 -11848 -28450 -11832
rect -28577 -11912 -28530 -11848
rect -28466 -11912 -28450 -11848
rect -28577 -11928 -28450 -11912
rect -28577 -11992 -28530 -11928
rect -28466 -11992 -28450 -11928
rect -28577 -12008 -28450 -11992
rect -28577 -12072 -28530 -12008
rect -28466 -12072 -28450 -12008
rect -28577 -12088 -28450 -12072
rect -28577 -12152 -28530 -12088
rect -28466 -12152 -28450 -12088
rect -28577 -12168 -28450 -12152
rect -28577 -12232 -28530 -12168
rect -28466 -12232 -28450 -12168
rect -28577 -12248 -28450 -12232
rect -28577 -12312 -28530 -12248
rect -28466 -12312 -28450 -12248
rect -28577 -12328 -28450 -12312
rect -28577 -12392 -28530 -12328
rect -28466 -12392 -28450 -12328
rect -28577 -12408 -28450 -12392
rect -28577 -12472 -28530 -12408
rect -28466 -12472 -28450 -12408
rect -28577 -12488 -28450 -12472
rect -28577 -12552 -28530 -12488
rect -28466 -12552 -28450 -12488
rect -28577 -12568 -28450 -12552
rect -28577 -12632 -28530 -12568
rect -28466 -12632 -28450 -12568
rect -28577 -12648 -28450 -12632
rect -28577 -12712 -28530 -12648
rect -28466 -12712 -28450 -12648
rect -28577 -12728 -28450 -12712
rect -28577 -12792 -28530 -12728
rect -28466 -12792 -28450 -12728
rect -28577 -12808 -28450 -12792
rect -28577 -12872 -28530 -12808
rect -28466 -12872 -28450 -12808
rect -28577 -12888 -28450 -12872
rect -28577 -12952 -28530 -12888
rect -28466 -12952 -28450 -12888
rect -28577 -12968 -28450 -12952
rect -28577 -13032 -28530 -12968
rect -28466 -13032 -28450 -12968
rect -28577 -13048 -28450 -13032
rect -28577 -13112 -28530 -13048
rect -28466 -13112 -28450 -13048
rect -28577 -13128 -28450 -13112
rect -28577 -13192 -28530 -13128
rect -28466 -13192 -28450 -13128
rect -28577 -13208 -28450 -13192
rect -28577 -13272 -28530 -13208
rect -28466 -13272 -28450 -13208
rect -28577 -13288 -28450 -13272
rect -28577 -13352 -28530 -13288
rect -28466 -13352 -28450 -13288
rect -28577 -13368 -28450 -13352
rect -28577 -13432 -28530 -13368
rect -28466 -13432 -28450 -13368
rect -28577 -13448 -28450 -13432
rect -28577 -13512 -28530 -13448
rect -28466 -13512 -28450 -13448
rect -28577 -13528 -28450 -13512
rect -28577 -13592 -28530 -13528
rect -28466 -13592 -28450 -13528
rect -28577 -13608 -28450 -13592
rect -28577 -13672 -28530 -13608
rect -28466 -13672 -28450 -13608
rect -28577 -13688 -28450 -13672
rect -28577 -13752 -28530 -13688
rect -28466 -13752 -28450 -13688
rect -28577 -13768 -28450 -13752
rect -28577 -13832 -28530 -13768
rect -28466 -13832 -28450 -13768
rect -28577 -13848 -28450 -13832
rect -28577 -13912 -28530 -13848
rect -28466 -13912 -28450 -13848
rect -28577 -13928 -28450 -13912
rect -28577 -13992 -28530 -13928
rect -28466 -13992 -28450 -13928
rect -28577 -14008 -28450 -13992
rect -28577 -14072 -28530 -14008
rect -28466 -14072 -28450 -14008
rect -28577 -14088 -28450 -14072
rect -28577 -14152 -28530 -14088
rect -28466 -14152 -28450 -14088
rect -28577 -14168 -28450 -14152
rect -28577 -14232 -28530 -14168
rect -28466 -14232 -28450 -14168
rect -28577 -14248 -28450 -14232
rect -28577 -14312 -28530 -14248
rect -28466 -14312 -28450 -14248
rect -28577 -14328 -28450 -14312
rect -28577 -14392 -28530 -14328
rect -28466 -14392 -28450 -14328
rect -28577 -14408 -28450 -14392
rect -28577 -14472 -28530 -14408
rect -28466 -14472 -28450 -14408
rect -28577 -14488 -28450 -14472
rect -28577 -14552 -28530 -14488
rect -28466 -14552 -28450 -14488
rect -28577 -14568 -28450 -14552
rect -28577 -14632 -28530 -14568
rect -28466 -14632 -28450 -14568
rect -28577 -14648 -28450 -14632
rect -28577 -14712 -28530 -14648
rect -28466 -14712 -28450 -14648
rect -28577 -14728 -28450 -14712
rect -28577 -14792 -28530 -14728
rect -28466 -14792 -28450 -14728
rect -28577 -14808 -28450 -14792
rect -28577 -14872 -28530 -14808
rect -28466 -14872 -28450 -14808
rect -28577 -14888 -28450 -14872
rect -28577 -14952 -28530 -14888
rect -28466 -14952 -28450 -14888
rect -28577 -14968 -28450 -14952
rect -28577 -15032 -28530 -14968
rect -28466 -15032 -28450 -14968
rect -28577 -15048 -28450 -15032
rect -28577 -15112 -28530 -15048
rect -28466 -15112 -28450 -15048
rect -28577 -15128 -28450 -15112
rect -28577 -15192 -28530 -15128
rect -28466 -15192 -28450 -15128
rect -28577 -15208 -28450 -15192
rect -28577 -15272 -28530 -15208
rect -28466 -15272 -28450 -15208
rect -28577 -15288 -28450 -15272
rect -28577 -15352 -28530 -15288
rect -28466 -15352 -28450 -15288
rect -28577 -15368 -28450 -15352
rect -28577 -15432 -28530 -15368
rect -28466 -15432 -28450 -15368
rect -28577 -15448 -28450 -15432
rect -28577 -15512 -28530 -15448
rect -28466 -15512 -28450 -15448
rect -28577 -15528 -28450 -15512
rect -34896 -15608 -34769 -15592
rect -34896 -15672 -34849 -15608
rect -34785 -15672 -34769 -15608
rect -34896 -15688 -34769 -15672
rect -34896 -15812 -34792 -15688
rect -34896 -15828 -34769 -15812
rect -34896 -15892 -34849 -15828
rect -34785 -15892 -34769 -15828
rect -34896 -15908 -34769 -15892
rect -41215 -15988 -41088 -15972
rect -41215 -16052 -41168 -15988
rect -41104 -16052 -41088 -15988
rect -41215 -16068 -41088 -16052
rect -41215 -16132 -41168 -16068
rect -41104 -16132 -41088 -16068
rect -41215 -16148 -41088 -16132
rect -41215 -16212 -41168 -16148
rect -41104 -16212 -41088 -16148
rect -41215 -16228 -41088 -16212
rect -41215 -16292 -41168 -16228
rect -41104 -16292 -41088 -16228
rect -41215 -16308 -41088 -16292
rect -41215 -16372 -41168 -16308
rect -41104 -16372 -41088 -16308
rect -41215 -16388 -41088 -16372
rect -41215 -16452 -41168 -16388
rect -41104 -16452 -41088 -16388
rect -41215 -16468 -41088 -16452
rect -41215 -16532 -41168 -16468
rect -41104 -16532 -41088 -16468
rect -41215 -16548 -41088 -16532
rect -41215 -16612 -41168 -16548
rect -41104 -16612 -41088 -16548
rect -41215 -16628 -41088 -16612
rect -41215 -16692 -41168 -16628
rect -41104 -16692 -41088 -16628
rect -41215 -16708 -41088 -16692
rect -41215 -16772 -41168 -16708
rect -41104 -16772 -41088 -16708
rect -41215 -16788 -41088 -16772
rect -41215 -16852 -41168 -16788
rect -41104 -16852 -41088 -16788
rect -41215 -16868 -41088 -16852
rect -41215 -16932 -41168 -16868
rect -41104 -16932 -41088 -16868
rect -41215 -16948 -41088 -16932
rect -41215 -17012 -41168 -16948
rect -41104 -17012 -41088 -16948
rect -41215 -17028 -41088 -17012
rect -41215 -17092 -41168 -17028
rect -41104 -17092 -41088 -17028
rect -41215 -17108 -41088 -17092
rect -41215 -17172 -41168 -17108
rect -41104 -17172 -41088 -17108
rect -41215 -17188 -41088 -17172
rect -41215 -17252 -41168 -17188
rect -41104 -17252 -41088 -17188
rect -41215 -17268 -41088 -17252
rect -41215 -17332 -41168 -17268
rect -41104 -17332 -41088 -17268
rect -41215 -17348 -41088 -17332
rect -41215 -17412 -41168 -17348
rect -41104 -17412 -41088 -17348
rect -41215 -17428 -41088 -17412
rect -41215 -17492 -41168 -17428
rect -41104 -17492 -41088 -17428
rect -41215 -17508 -41088 -17492
rect -41215 -17572 -41168 -17508
rect -41104 -17572 -41088 -17508
rect -41215 -17588 -41088 -17572
rect -41215 -17652 -41168 -17588
rect -41104 -17652 -41088 -17588
rect -41215 -17668 -41088 -17652
rect -41215 -17732 -41168 -17668
rect -41104 -17732 -41088 -17668
rect -41215 -17748 -41088 -17732
rect -41215 -17812 -41168 -17748
rect -41104 -17812 -41088 -17748
rect -41215 -17828 -41088 -17812
rect -41215 -17892 -41168 -17828
rect -41104 -17892 -41088 -17828
rect -41215 -17908 -41088 -17892
rect -41215 -17972 -41168 -17908
rect -41104 -17972 -41088 -17908
rect -41215 -17988 -41088 -17972
rect -41215 -18052 -41168 -17988
rect -41104 -18052 -41088 -17988
rect -41215 -18068 -41088 -18052
rect -41215 -18132 -41168 -18068
rect -41104 -18132 -41088 -18068
rect -41215 -18148 -41088 -18132
rect -41215 -18212 -41168 -18148
rect -41104 -18212 -41088 -18148
rect -41215 -18228 -41088 -18212
rect -41215 -18292 -41168 -18228
rect -41104 -18292 -41088 -18228
rect -41215 -18308 -41088 -18292
rect -41215 -18372 -41168 -18308
rect -41104 -18372 -41088 -18308
rect -41215 -18388 -41088 -18372
rect -41215 -18452 -41168 -18388
rect -41104 -18452 -41088 -18388
rect -41215 -18468 -41088 -18452
rect -41215 -18532 -41168 -18468
rect -41104 -18532 -41088 -18468
rect -41215 -18548 -41088 -18532
rect -41215 -18612 -41168 -18548
rect -41104 -18612 -41088 -18548
rect -41215 -18628 -41088 -18612
rect -41215 -18692 -41168 -18628
rect -41104 -18692 -41088 -18628
rect -41215 -18708 -41088 -18692
rect -41215 -18772 -41168 -18708
rect -41104 -18772 -41088 -18708
rect -41215 -18788 -41088 -18772
rect -41215 -18852 -41168 -18788
rect -41104 -18852 -41088 -18788
rect -41215 -18868 -41088 -18852
rect -41215 -18932 -41168 -18868
rect -41104 -18932 -41088 -18868
rect -41215 -18948 -41088 -18932
rect -41215 -19012 -41168 -18948
rect -41104 -19012 -41088 -18948
rect -41215 -19028 -41088 -19012
rect -41215 -19092 -41168 -19028
rect -41104 -19092 -41088 -19028
rect -41215 -19108 -41088 -19092
rect -41215 -19172 -41168 -19108
rect -41104 -19172 -41088 -19108
rect -41215 -19188 -41088 -19172
rect -41215 -19252 -41168 -19188
rect -41104 -19252 -41088 -19188
rect -41215 -19268 -41088 -19252
rect -41215 -19332 -41168 -19268
rect -41104 -19332 -41088 -19268
rect -41215 -19348 -41088 -19332
rect -41215 -19412 -41168 -19348
rect -41104 -19412 -41088 -19348
rect -41215 -19428 -41088 -19412
rect -41215 -19492 -41168 -19428
rect -41104 -19492 -41088 -19428
rect -41215 -19508 -41088 -19492
rect -41215 -19572 -41168 -19508
rect -41104 -19572 -41088 -19508
rect -41215 -19588 -41088 -19572
rect -41215 -19652 -41168 -19588
rect -41104 -19652 -41088 -19588
rect -41215 -19668 -41088 -19652
rect -41215 -19732 -41168 -19668
rect -41104 -19732 -41088 -19668
rect -41215 -19748 -41088 -19732
rect -41215 -19812 -41168 -19748
rect -41104 -19812 -41088 -19748
rect -41215 -19828 -41088 -19812
rect -41215 -19892 -41168 -19828
rect -41104 -19892 -41088 -19828
rect -41215 -19908 -41088 -19892
rect -41215 -19972 -41168 -19908
rect -41104 -19972 -41088 -19908
rect -41215 -19988 -41088 -19972
rect -41215 -20052 -41168 -19988
rect -41104 -20052 -41088 -19988
rect -41215 -20068 -41088 -20052
rect -41215 -20132 -41168 -20068
rect -41104 -20132 -41088 -20068
rect -41215 -20148 -41088 -20132
rect -41215 -20212 -41168 -20148
rect -41104 -20212 -41088 -20148
rect -41215 -20228 -41088 -20212
rect -41215 -20292 -41168 -20228
rect -41104 -20292 -41088 -20228
rect -41215 -20308 -41088 -20292
rect -41215 -20372 -41168 -20308
rect -41104 -20372 -41088 -20308
rect -41215 -20388 -41088 -20372
rect -41215 -20452 -41168 -20388
rect -41104 -20452 -41088 -20388
rect -41215 -20468 -41088 -20452
rect -41215 -20532 -41168 -20468
rect -41104 -20532 -41088 -20468
rect -41215 -20548 -41088 -20532
rect -41215 -20612 -41168 -20548
rect -41104 -20612 -41088 -20548
rect -41215 -20628 -41088 -20612
rect -41215 -20692 -41168 -20628
rect -41104 -20692 -41088 -20628
rect -41215 -20708 -41088 -20692
rect -41215 -20772 -41168 -20708
rect -41104 -20772 -41088 -20708
rect -41215 -20788 -41088 -20772
rect -41215 -20852 -41168 -20788
rect -41104 -20852 -41088 -20788
rect -41215 -20868 -41088 -20852
rect -41215 -20932 -41168 -20868
rect -41104 -20932 -41088 -20868
rect -41215 -20948 -41088 -20932
rect -41215 -21012 -41168 -20948
rect -41104 -21012 -41088 -20948
rect -41215 -21028 -41088 -21012
rect -41215 -21092 -41168 -21028
rect -41104 -21092 -41088 -21028
rect -41215 -21108 -41088 -21092
rect -41215 -21172 -41168 -21108
rect -41104 -21172 -41088 -21108
rect -41215 -21188 -41088 -21172
rect -41215 -21252 -41168 -21188
rect -41104 -21252 -41088 -21188
rect -41215 -21268 -41088 -21252
rect -41215 -21332 -41168 -21268
rect -41104 -21332 -41088 -21268
rect -41215 -21348 -41088 -21332
rect -41215 -21412 -41168 -21348
rect -41104 -21412 -41088 -21348
rect -41215 -21428 -41088 -21412
rect -41215 -21492 -41168 -21428
rect -41104 -21492 -41088 -21428
rect -41215 -21508 -41088 -21492
rect -41215 -21572 -41168 -21508
rect -41104 -21572 -41088 -21508
rect -41215 -21588 -41088 -21572
rect -41215 -21652 -41168 -21588
rect -41104 -21652 -41088 -21588
rect -41215 -21668 -41088 -21652
rect -41215 -21732 -41168 -21668
rect -41104 -21732 -41088 -21668
rect -41215 -21748 -41088 -21732
rect -41215 -21812 -41168 -21748
rect -41104 -21812 -41088 -21748
rect -41215 -21828 -41088 -21812
rect -44335 -22239 -44231 -21861
rect -41215 -21892 -41168 -21828
rect -41104 -21892 -41088 -21828
rect -40925 -15948 -35003 -15939
rect -40925 -21852 -40916 -15948
rect -35012 -21852 -35003 -15948
rect -40925 -21861 -35003 -21852
rect -34896 -15972 -34849 -15908
rect -34785 -15972 -34769 -15908
rect -31697 -15939 -31593 -15561
rect -28577 -15592 -28530 -15528
rect -28466 -15592 -28450 -15528
rect -28287 -9648 -22365 -9639
rect -28287 -15552 -28278 -9648
rect -22374 -15552 -22365 -9648
rect -28287 -15561 -22365 -15552
rect -22258 -9672 -22211 -9608
rect -22147 -9672 -22131 -9608
rect -19059 -9639 -18955 -9261
rect -15939 -9292 -15892 -9228
rect -15828 -9292 -15812 -9228
rect -15649 -3348 -9727 -3339
rect -15649 -9252 -15640 -3348
rect -9736 -9252 -9727 -3348
rect -15649 -9261 -9727 -9252
rect -9620 -3372 -9573 -3308
rect -9509 -3372 -9493 -3308
rect -6421 -3339 -6317 -2961
rect -3301 -2992 -3254 -2928
rect -3190 -2992 -3174 -2928
rect -3011 2952 2911 2961
rect -3011 -2952 -3002 2952
rect 2902 -2952 2911 2952
rect -3011 -2961 2911 -2952
rect 3018 2928 3065 2992
rect 3129 2928 3145 2992
rect 6217 2961 6321 3339
rect 9337 3308 9384 3372
rect 9448 3308 9464 3372
rect 9627 9252 15549 9261
rect 9627 3348 9636 9252
rect 15540 3348 15549 9252
rect 9627 3339 15549 3348
rect 15656 9228 15703 9292
rect 15767 9228 15783 9292
rect 18855 9261 18959 9639
rect 21975 9608 22022 9672
rect 22086 9608 22102 9672
rect 22265 15552 28187 15561
rect 22265 9648 22274 15552
rect 28178 9648 28187 15552
rect 22265 9639 28187 9648
rect 28294 15528 28341 15592
rect 28405 15528 28421 15592
rect 31493 15561 31597 15939
rect 34613 15908 34660 15972
rect 34724 15908 34740 15972
rect 34903 21852 40825 21861
rect 34903 15948 34912 21852
rect 40816 15948 40825 21852
rect 34903 15939 40825 15948
rect 40932 21828 40979 21892
rect 41043 21828 41059 21892
rect 44131 21861 44235 22239
rect 47251 22208 47298 22272
rect 47362 22208 47378 22272
rect 47251 22192 47378 22208
rect 47251 22128 47298 22192
rect 47362 22128 47378 22192
rect 47251 22112 47378 22128
rect 47251 21988 47355 22112
rect 47251 21972 47378 21988
rect 47251 21908 47298 21972
rect 47362 21908 47378 21972
rect 47251 21892 47378 21908
rect 40932 21812 41059 21828
rect 40932 21748 40979 21812
rect 41043 21748 41059 21812
rect 40932 21732 41059 21748
rect 40932 21668 40979 21732
rect 41043 21668 41059 21732
rect 40932 21652 41059 21668
rect 40932 21588 40979 21652
rect 41043 21588 41059 21652
rect 40932 21572 41059 21588
rect 40932 21508 40979 21572
rect 41043 21508 41059 21572
rect 40932 21492 41059 21508
rect 40932 21428 40979 21492
rect 41043 21428 41059 21492
rect 40932 21412 41059 21428
rect 40932 21348 40979 21412
rect 41043 21348 41059 21412
rect 40932 21332 41059 21348
rect 40932 21268 40979 21332
rect 41043 21268 41059 21332
rect 40932 21252 41059 21268
rect 40932 21188 40979 21252
rect 41043 21188 41059 21252
rect 40932 21172 41059 21188
rect 40932 21108 40979 21172
rect 41043 21108 41059 21172
rect 40932 21092 41059 21108
rect 40932 21028 40979 21092
rect 41043 21028 41059 21092
rect 40932 21012 41059 21028
rect 40932 20948 40979 21012
rect 41043 20948 41059 21012
rect 40932 20932 41059 20948
rect 40932 20868 40979 20932
rect 41043 20868 41059 20932
rect 40932 20852 41059 20868
rect 40932 20788 40979 20852
rect 41043 20788 41059 20852
rect 40932 20772 41059 20788
rect 40932 20708 40979 20772
rect 41043 20708 41059 20772
rect 40932 20692 41059 20708
rect 40932 20628 40979 20692
rect 41043 20628 41059 20692
rect 40932 20612 41059 20628
rect 40932 20548 40979 20612
rect 41043 20548 41059 20612
rect 40932 20532 41059 20548
rect 40932 20468 40979 20532
rect 41043 20468 41059 20532
rect 40932 20452 41059 20468
rect 40932 20388 40979 20452
rect 41043 20388 41059 20452
rect 40932 20372 41059 20388
rect 40932 20308 40979 20372
rect 41043 20308 41059 20372
rect 40932 20292 41059 20308
rect 40932 20228 40979 20292
rect 41043 20228 41059 20292
rect 40932 20212 41059 20228
rect 40932 20148 40979 20212
rect 41043 20148 41059 20212
rect 40932 20132 41059 20148
rect 40932 20068 40979 20132
rect 41043 20068 41059 20132
rect 40932 20052 41059 20068
rect 40932 19988 40979 20052
rect 41043 19988 41059 20052
rect 40932 19972 41059 19988
rect 40932 19908 40979 19972
rect 41043 19908 41059 19972
rect 40932 19892 41059 19908
rect 40932 19828 40979 19892
rect 41043 19828 41059 19892
rect 40932 19812 41059 19828
rect 40932 19748 40979 19812
rect 41043 19748 41059 19812
rect 40932 19732 41059 19748
rect 40932 19668 40979 19732
rect 41043 19668 41059 19732
rect 40932 19652 41059 19668
rect 40932 19588 40979 19652
rect 41043 19588 41059 19652
rect 40932 19572 41059 19588
rect 40932 19508 40979 19572
rect 41043 19508 41059 19572
rect 40932 19492 41059 19508
rect 40932 19428 40979 19492
rect 41043 19428 41059 19492
rect 40932 19412 41059 19428
rect 40932 19348 40979 19412
rect 41043 19348 41059 19412
rect 40932 19332 41059 19348
rect 40932 19268 40979 19332
rect 41043 19268 41059 19332
rect 40932 19252 41059 19268
rect 40932 19188 40979 19252
rect 41043 19188 41059 19252
rect 40932 19172 41059 19188
rect 40932 19108 40979 19172
rect 41043 19108 41059 19172
rect 40932 19092 41059 19108
rect 40932 19028 40979 19092
rect 41043 19028 41059 19092
rect 40932 19012 41059 19028
rect 40932 18948 40979 19012
rect 41043 18948 41059 19012
rect 40932 18932 41059 18948
rect 40932 18868 40979 18932
rect 41043 18868 41059 18932
rect 40932 18852 41059 18868
rect 40932 18788 40979 18852
rect 41043 18788 41059 18852
rect 40932 18772 41059 18788
rect 40932 18708 40979 18772
rect 41043 18708 41059 18772
rect 40932 18692 41059 18708
rect 40932 18628 40979 18692
rect 41043 18628 41059 18692
rect 40932 18612 41059 18628
rect 40932 18548 40979 18612
rect 41043 18548 41059 18612
rect 40932 18532 41059 18548
rect 40932 18468 40979 18532
rect 41043 18468 41059 18532
rect 40932 18452 41059 18468
rect 40932 18388 40979 18452
rect 41043 18388 41059 18452
rect 40932 18372 41059 18388
rect 40932 18308 40979 18372
rect 41043 18308 41059 18372
rect 40932 18292 41059 18308
rect 40932 18228 40979 18292
rect 41043 18228 41059 18292
rect 40932 18212 41059 18228
rect 40932 18148 40979 18212
rect 41043 18148 41059 18212
rect 40932 18132 41059 18148
rect 40932 18068 40979 18132
rect 41043 18068 41059 18132
rect 40932 18052 41059 18068
rect 40932 17988 40979 18052
rect 41043 17988 41059 18052
rect 40932 17972 41059 17988
rect 40932 17908 40979 17972
rect 41043 17908 41059 17972
rect 40932 17892 41059 17908
rect 40932 17828 40979 17892
rect 41043 17828 41059 17892
rect 40932 17812 41059 17828
rect 40932 17748 40979 17812
rect 41043 17748 41059 17812
rect 40932 17732 41059 17748
rect 40932 17668 40979 17732
rect 41043 17668 41059 17732
rect 40932 17652 41059 17668
rect 40932 17588 40979 17652
rect 41043 17588 41059 17652
rect 40932 17572 41059 17588
rect 40932 17508 40979 17572
rect 41043 17508 41059 17572
rect 40932 17492 41059 17508
rect 40932 17428 40979 17492
rect 41043 17428 41059 17492
rect 40932 17412 41059 17428
rect 40932 17348 40979 17412
rect 41043 17348 41059 17412
rect 40932 17332 41059 17348
rect 40932 17268 40979 17332
rect 41043 17268 41059 17332
rect 40932 17252 41059 17268
rect 40932 17188 40979 17252
rect 41043 17188 41059 17252
rect 40932 17172 41059 17188
rect 40932 17108 40979 17172
rect 41043 17108 41059 17172
rect 40932 17092 41059 17108
rect 40932 17028 40979 17092
rect 41043 17028 41059 17092
rect 40932 17012 41059 17028
rect 40932 16948 40979 17012
rect 41043 16948 41059 17012
rect 40932 16932 41059 16948
rect 40932 16868 40979 16932
rect 41043 16868 41059 16932
rect 40932 16852 41059 16868
rect 40932 16788 40979 16852
rect 41043 16788 41059 16852
rect 40932 16772 41059 16788
rect 40932 16708 40979 16772
rect 41043 16708 41059 16772
rect 40932 16692 41059 16708
rect 40932 16628 40979 16692
rect 41043 16628 41059 16692
rect 40932 16612 41059 16628
rect 40932 16548 40979 16612
rect 41043 16548 41059 16612
rect 40932 16532 41059 16548
rect 40932 16468 40979 16532
rect 41043 16468 41059 16532
rect 40932 16452 41059 16468
rect 40932 16388 40979 16452
rect 41043 16388 41059 16452
rect 40932 16372 41059 16388
rect 40932 16308 40979 16372
rect 41043 16308 41059 16372
rect 40932 16292 41059 16308
rect 40932 16228 40979 16292
rect 41043 16228 41059 16292
rect 40932 16212 41059 16228
rect 40932 16148 40979 16212
rect 41043 16148 41059 16212
rect 40932 16132 41059 16148
rect 40932 16068 40979 16132
rect 41043 16068 41059 16132
rect 40932 16052 41059 16068
rect 40932 15988 40979 16052
rect 41043 15988 41059 16052
rect 40932 15972 41059 15988
rect 34613 15892 34740 15908
rect 34613 15828 34660 15892
rect 34724 15828 34740 15892
rect 34613 15812 34740 15828
rect 34613 15688 34717 15812
rect 34613 15672 34740 15688
rect 34613 15608 34660 15672
rect 34724 15608 34740 15672
rect 34613 15592 34740 15608
rect 28294 15512 28421 15528
rect 28294 15448 28341 15512
rect 28405 15448 28421 15512
rect 28294 15432 28421 15448
rect 28294 15368 28341 15432
rect 28405 15368 28421 15432
rect 28294 15352 28421 15368
rect 28294 15288 28341 15352
rect 28405 15288 28421 15352
rect 28294 15272 28421 15288
rect 28294 15208 28341 15272
rect 28405 15208 28421 15272
rect 28294 15192 28421 15208
rect 28294 15128 28341 15192
rect 28405 15128 28421 15192
rect 28294 15112 28421 15128
rect 28294 15048 28341 15112
rect 28405 15048 28421 15112
rect 28294 15032 28421 15048
rect 28294 14968 28341 15032
rect 28405 14968 28421 15032
rect 28294 14952 28421 14968
rect 28294 14888 28341 14952
rect 28405 14888 28421 14952
rect 28294 14872 28421 14888
rect 28294 14808 28341 14872
rect 28405 14808 28421 14872
rect 28294 14792 28421 14808
rect 28294 14728 28341 14792
rect 28405 14728 28421 14792
rect 28294 14712 28421 14728
rect 28294 14648 28341 14712
rect 28405 14648 28421 14712
rect 28294 14632 28421 14648
rect 28294 14568 28341 14632
rect 28405 14568 28421 14632
rect 28294 14552 28421 14568
rect 28294 14488 28341 14552
rect 28405 14488 28421 14552
rect 28294 14472 28421 14488
rect 28294 14408 28341 14472
rect 28405 14408 28421 14472
rect 28294 14392 28421 14408
rect 28294 14328 28341 14392
rect 28405 14328 28421 14392
rect 28294 14312 28421 14328
rect 28294 14248 28341 14312
rect 28405 14248 28421 14312
rect 28294 14232 28421 14248
rect 28294 14168 28341 14232
rect 28405 14168 28421 14232
rect 28294 14152 28421 14168
rect 28294 14088 28341 14152
rect 28405 14088 28421 14152
rect 28294 14072 28421 14088
rect 28294 14008 28341 14072
rect 28405 14008 28421 14072
rect 28294 13992 28421 14008
rect 28294 13928 28341 13992
rect 28405 13928 28421 13992
rect 28294 13912 28421 13928
rect 28294 13848 28341 13912
rect 28405 13848 28421 13912
rect 28294 13832 28421 13848
rect 28294 13768 28341 13832
rect 28405 13768 28421 13832
rect 28294 13752 28421 13768
rect 28294 13688 28341 13752
rect 28405 13688 28421 13752
rect 28294 13672 28421 13688
rect 28294 13608 28341 13672
rect 28405 13608 28421 13672
rect 28294 13592 28421 13608
rect 28294 13528 28341 13592
rect 28405 13528 28421 13592
rect 28294 13512 28421 13528
rect 28294 13448 28341 13512
rect 28405 13448 28421 13512
rect 28294 13432 28421 13448
rect 28294 13368 28341 13432
rect 28405 13368 28421 13432
rect 28294 13352 28421 13368
rect 28294 13288 28341 13352
rect 28405 13288 28421 13352
rect 28294 13272 28421 13288
rect 28294 13208 28341 13272
rect 28405 13208 28421 13272
rect 28294 13192 28421 13208
rect 28294 13128 28341 13192
rect 28405 13128 28421 13192
rect 28294 13112 28421 13128
rect 28294 13048 28341 13112
rect 28405 13048 28421 13112
rect 28294 13032 28421 13048
rect 28294 12968 28341 13032
rect 28405 12968 28421 13032
rect 28294 12952 28421 12968
rect 28294 12888 28341 12952
rect 28405 12888 28421 12952
rect 28294 12872 28421 12888
rect 28294 12808 28341 12872
rect 28405 12808 28421 12872
rect 28294 12792 28421 12808
rect 28294 12728 28341 12792
rect 28405 12728 28421 12792
rect 28294 12712 28421 12728
rect 28294 12648 28341 12712
rect 28405 12648 28421 12712
rect 28294 12632 28421 12648
rect 28294 12568 28341 12632
rect 28405 12568 28421 12632
rect 28294 12552 28421 12568
rect 28294 12488 28341 12552
rect 28405 12488 28421 12552
rect 28294 12472 28421 12488
rect 28294 12408 28341 12472
rect 28405 12408 28421 12472
rect 28294 12392 28421 12408
rect 28294 12328 28341 12392
rect 28405 12328 28421 12392
rect 28294 12312 28421 12328
rect 28294 12248 28341 12312
rect 28405 12248 28421 12312
rect 28294 12232 28421 12248
rect 28294 12168 28341 12232
rect 28405 12168 28421 12232
rect 28294 12152 28421 12168
rect 28294 12088 28341 12152
rect 28405 12088 28421 12152
rect 28294 12072 28421 12088
rect 28294 12008 28341 12072
rect 28405 12008 28421 12072
rect 28294 11992 28421 12008
rect 28294 11928 28341 11992
rect 28405 11928 28421 11992
rect 28294 11912 28421 11928
rect 28294 11848 28341 11912
rect 28405 11848 28421 11912
rect 28294 11832 28421 11848
rect 28294 11768 28341 11832
rect 28405 11768 28421 11832
rect 28294 11752 28421 11768
rect 28294 11688 28341 11752
rect 28405 11688 28421 11752
rect 28294 11672 28421 11688
rect 28294 11608 28341 11672
rect 28405 11608 28421 11672
rect 28294 11592 28421 11608
rect 28294 11528 28341 11592
rect 28405 11528 28421 11592
rect 28294 11512 28421 11528
rect 28294 11448 28341 11512
rect 28405 11448 28421 11512
rect 28294 11432 28421 11448
rect 28294 11368 28341 11432
rect 28405 11368 28421 11432
rect 28294 11352 28421 11368
rect 28294 11288 28341 11352
rect 28405 11288 28421 11352
rect 28294 11272 28421 11288
rect 28294 11208 28341 11272
rect 28405 11208 28421 11272
rect 28294 11192 28421 11208
rect 28294 11128 28341 11192
rect 28405 11128 28421 11192
rect 28294 11112 28421 11128
rect 28294 11048 28341 11112
rect 28405 11048 28421 11112
rect 28294 11032 28421 11048
rect 28294 10968 28341 11032
rect 28405 10968 28421 11032
rect 28294 10952 28421 10968
rect 28294 10888 28341 10952
rect 28405 10888 28421 10952
rect 28294 10872 28421 10888
rect 28294 10808 28341 10872
rect 28405 10808 28421 10872
rect 28294 10792 28421 10808
rect 28294 10728 28341 10792
rect 28405 10728 28421 10792
rect 28294 10712 28421 10728
rect 28294 10648 28341 10712
rect 28405 10648 28421 10712
rect 28294 10632 28421 10648
rect 28294 10568 28341 10632
rect 28405 10568 28421 10632
rect 28294 10552 28421 10568
rect 28294 10488 28341 10552
rect 28405 10488 28421 10552
rect 28294 10472 28421 10488
rect 28294 10408 28341 10472
rect 28405 10408 28421 10472
rect 28294 10392 28421 10408
rect 28294 10328 28341 10392
rect 28405 10328 28421 10392
rect 28294 10312 28421 10328
rect 28294 10248 28341 10312
rect 28405 10248 28421 10312
rect 28294 10232 28421 10248
rect 28294 10168 28341 10232
rect 28405 10168 28421 10232
rect 28294 10152 28421 10168
rect 28294 10088 28341 10152
rect 28405 10088 28421 10152
rect 28294 10072 28421 10088
rect 28294 10008 28341 10072
rect 28405 10008 28421 10072
rect 28294 9992 28421 10008
rect 28294 9928 28341 9992
rect 28405 9928 28421 9992
rect 28294 9912 28421 9928
rect 28294 9848 28341 9912
rect 28405 9848 28421 9912
rect 28294 9832 28421 9848
rect 28294 9768 28341 9832
rect 28405 9768 28421 9832
rect 28294 9752 28421 9768
rect 28294 9688 28341 9752
rect 28405 9688 28421 9752
rect 28294 9672 28421 9688
rect 21975 9592 22102 9608
rect 21975 9528 22022 9592
rect 22086 9528 22102 9592
rect 21975 9512 22102 9528
rect 21975 9388 22079 9512
rect 21975 9372 22102 9388
rect 21975 9308 22022 9372
rect 22086 9308 22102 9372
rect 21975 9292 22102 9308
rect 15656 9212 15783 9228
rect 15656 9148 15703 9212
rect 15767 9148 15783 9212
rect 15656 9132 15783 9148
rect 15656 9068 15703 9132
rect 15767 9068 15783 9132
rect 15656 9052 15783 9068
rect 15656 8988 15703 9052
rect 15767 8988 15783 9052
rect 15656 8972 15783 8988
rect 15656 8908 15703 8972
rect 15767 8908 15783 8972
rect 15656 8892 15783 8908
rect 15656 8828 15703 8892
rect 15767 8828 15783 8892
rect 15656 8812 15783 8828
rect 15656 8748 15703 8812
rect 15767 8748 15783 8812
rect 15656 8732 15783 8748
rect 15656 8668 15703 8732
rect 15767 8668 15783 8732
rect 15656 8652 15783 8668
rect 15656 8588 15703 8652
rect 15767 8588 15783 8652
rect 15656 8572 15783 8588
rect 15656 8508 15703 8572
rect 15767 8508 15783 8572
rect 15656 8492 15783 8508
rect 15656 8428 15703 8492
rect 15767 8428 15783 8492
rect 15656 8412 15783 8428
rect 15656 8348 15703 8412
rect 15767 8348 15783 8412
rect 15656 8332 15783 8348
rect 15656 8268 15703 8332
rect 15767 8268 15783 8332
rect 15656 8252 15783 8268
rect 15656 8188 15703 8252
rect 15767 8188 15783 8252
rect 15656 8172 15783 8188
rect 15656 8108 15703 8172
rect 15767 8108 15783 8172
rect 15656 8092 15783 8108
rect 15656 8028 15703 8092
rect 15767 8028 15783 8092
rect 15656 8012 15783 8028
rect 15656 7948 15703 8012
rect 15767 7948 15783 8012
rect 15656 7932 15783 7948
rect 15656 7868 15703 7932
rect 15767 7868 15783 7932
rect 15656 7852 15783 7868
rect 15656 7788 15703 7852
rect 15767 7788 15783 7852
rect 15656 7772 15783 7788
rect 15656 7708 15703 7772
rect 15767 7708 15783 7772
rect 15656 7692 15783 7708
rect 15656 7628 15703 7692
rect 15767 7628 15783 7692
rect 15656 7612 15783 7628
rect 15656 7548 15703 7612
rect 15767 7548 15783 7612
rect 15656 7532 15783 7548
rect 15656 7468 15703 7532
rect 15767 7468 15783 7532
rect 15656 7452 15783 7468
rect 15656 7388 15703 7452
rect 15767 7388 15783 7452
rect 15656 7372 15783 7388
rect 15656 7308 15703 7372
rect 15767 7308 15783 7372
rect 15656 7292 15783 7308
rect 15656 7228 15703 7292
rect 15767 7228 15783 7292
rect 15656 7212 15783 7228
rect 15656 7148 15703 7212
rect 15767 7148 15783 7212
rect 15656 7132 15783 7148
rect 15656 7068 15703 7132
rect 15767 7068 15783 7132
rect 15656 7052 15783 7068
rect 15656 6988 15703 7052
rect 15767 6988 15783 7052
rect 15656 6972 15783 6988
rect 15656 6908 15703 6972
rect 15767 6908 15783 6972
rect 15656 6892 15783 6908
rect 15656 6828 15703 6892
rect 15767 6828 15783 6892
rect 15656 6812 15783 6828
rect 15656 6748 15703 6812
rect 15767 6748 15783 6812
rect 15656 6732 15783 6748
rect 15656 6668 15703 6732
rect 15767 6668 15783 6732
rect 15656 6652 15783 6668
rect 15656 6588 15703 6652
rect 15767 6588 15783 6652
rect 15656 6572 15783 6588
rect 15656 6508 15703 6572
rect 15767 6508 15783 6572
rect 15656 6492 15783 6508
rect 15656 6428 15703 6492
rect 15767 6428 15783 6492
rect 15656 6412 15783 6428
rect 15656 6348 15703 6412
rect 15767 6348 15783 6412
rect 15656 6332 15783 6348
rect 15656 6268 15703 6332
rect 15767 6268 15783 6332
rect 15656 6252 15783 6268
rect 15656 6188 15703 6252
rect 15767 6188 15783 6252
rect 15656 6172 15783 6188
rect 15656 6108 15703 6172
rect 15767 6108 15783 6172
rect 15656 6092 15783 6108
rect 15656 6028 15703 6092
rect 15767 6028 15783 6092
rect 15656 6012 15783 6028
rect 15656 5948 15703 6012
rect 15767 5948 15783 6012
rect 15656 5932 15783 5948
rect 15656 5868 15703 5932
rect 15767 5868 15783 5932
rect 15656 5852 15783 5868
rect 15656 5788 15703 5852
rect 15767 5788 15783 5852
rect 15656 5772 15783 5788
rect 15656 5708 15703 5772
rect 15767 5708 15783 5772
rect 15656 5692 15783 5708
rect 15656 5628 15703 5692
rect 15767 5628 15783 5692
rect 15656 5612 15783 5628
rect 15656 5548 15703 5612
rect 15767 5548 15783 5612
rect 15656 5532 15783 5548
rect 15656 5468 15703 5532
rect 15767 5468 15783 5532
rect 15656 5452 15783 5468
rect 15656 5388 15703 5452
rect 15767 5388 15783 5452
rect 15656 5372 15783 5388
rect 15656 5308 15703 5372
rect 15767 5308 15783 5372
rect 15656 5292 15783 5308
rect 15656 5228 15703 5292
rect 15767 5228 15783 5292
rect 15656 5212 15783 5228
rect 15656 5148 15703 5212
rect 15767 5148 15783 5212
rect 15656 5132 15783 5148
rect 15656 5068 15703 5132
rect 15767 5068 15783 5132
rect 15656 5052 15783 5068
rect 15656 4988 15703 5052
rect 15767 4988 15783 5052
rect 15656 4972 15783 4988
rect 15656 4908 15703 4972
rect 15767 4908 15783 4972
rect 15656 4892 15783 4908
rect 15656 4828 15703 4892
rect 15767 4828 15783 4892
rect 15656 4812 15783 4828
rect 15656 4748 15703 4812
rect 15767 4748 15783 4812
rect 15656 4732 15783 4748
rect 15656 4668 15703 4732
rect 15767 4668 15783 4732
rect 15656 4652 15783 4668
rect 15656 4588 15703 4652
rect 15767 4588 15783 4652
rect 15656 4572 15783 4588
rect 15656 4508 15703 4572
rect 15767 4508 15783 4572
rect 15656 4492 15783 4508
rect 15656 4428 15703 4492
rect 15767 4428 15783 4492
rect 15656 4412 15783 4428
rect 15656 4348 15703 4412
rect 15767 4348 15783 4412
rect 15656 4332 15783 4348
rect 15656 4268 15703 4332
rect 15767 4268 15783 4332
rect 15656 4252 15783 4268
rect 15656 4188 15703 4252
rect 15767 4188 15783 4252
rect 15656 4172 15783 4188
rect 15656 4108 15703 4172
rect 15767 4108 15783 4172
rect 15656 4092 15783 4108
rect 15656 4028 15703 4092
rect 15767 4028 15783 4092
rect 15656 4012 15783 4028
rect 15656 3948 15703 4012
rect 15767 3948 15783 4012
rect 15656 3932 15783 3948
rect 15656 3868 15703 3932
rect 15767 3868 15783 3932
rect 15656 3852 15783 3868
rect 15656 3788 15703 3852
rect 15767 3788 15783 3852
rect 15656 3772 15783 3788
rect 15656 3708 15703 3772
rect 15767 3708 15783 3772
rect 15656 3692 15783 3708
rect 15656 3628 15703 3692
rect 15767 3628 15783 3692
rect 15656 3612 15783 3628
rect 15656 3548 15703 3612
rect 15767 3548 15783 3612
rect 15656 3532 15783 3548
rect 15656 3468 15703 3532
rect 15767 3468 15783 3532
rect 15656 3452 15783 3468
rect 15656 3388 15703 3452
rect 15767 3388 15783 3452
rect 15656 3372 15783 3388
rect 9337 3292 9464 3308
rect 9337 3228 9384 3292
rect 9448 3228 9464 3292
rect 9337 3212 9464 3228
rect 9337 3088 9441 3212
rect 9337 3072 9464 3088
rect 9337 3008 9384 3072
rect 9448 3008 9464 3072
rect 9337 2992 9464 3008
rect 3018 2912 3145 2928
rect 3018 2848 3065 2912
rect 3129 2848 3145 2912
rect 3018 2832 3145 2848
rect 3018 2768 3065 2832
rect 3129 2768 3145 2832
rect 3018 2752 3145 2768
rect 3018 2688 3065 2752
rect 3129 2688 3145 2752
rect 3018 2672 3145 2688
rect 3018 2608 3065 2672
rect 3129 2608 3145 2672
rect 3018 2592 3145 2608
rect 3018 2528 3065 2592
rect 3129 2528 3145 2592
rect 3018 2512 3145 2528
rect 3018 2448 3065 2512
rect 3129 2448 3145 2512
rect 3018 2432 3145 2448
rect 3018 2368 3065 2432
rect 3129 2368 3145 2432
rect 3018 2352 3145 2368
rect 3018 2288 3065 2352
rect 3129 2288 3145 2352
rect 3018 2272 3145 2288
rect 3018 2208 3065 2272
rect 3129 2208 3145 2272
rect 3018 2192 3145 2208
rect 3018 2128 3065 2192
rect 3129 2128 3145 2192
rect 3018 2112 3145 2128
rect 3018 2048 3065 2112
rect 3129 2048 3145 2112
rect 3018 2032 3145 2048
rect 3018 1968 3065 2032
rect 3129 1968 3145 2032
rect 3018 1952 3145 1968
rect 3018 1888 3065 1952
rect 3129 1888 3145 1952
rect 3018 1872 3145 1888
rect 3018 1808 3065 1872
rect 3129 1808 3145 1872
rect 3018 1792 3145 1808
rect 3018 1728 3065 1792
rect 3129 1728 3145 1792
rect 3018 1712 3145 1728
rect 3018 1648 3065 1712
rect 3129 1648 3145 1712
rect 3018 1632 3145 1648
rect 3018 1568 3065 1632
rect 3129 1568 3145 1632
rect 3018 1552 3145 1568
rect 3018 1488 3065 1552
rect 3129 1488 3145 1552
rect 3018 1472 3145 1488
rect 3018 1408 3065 1472
rect 3129 1408 3145 1472
rect 3018 1392 3145 1408
rect 3018 1328 3065 1392
rect 3129 1328 3145 1392
rect 3018 1312 3145 1328
rect 3018 1248 3065 1312
rect 3129 1248 3145 1312
rect 3018 1232 3145 1248
rect 3018 1168 3065 1232
rect 3129 1168 3145 1232
rect 3018 1152 3145 1168
rect 3018 1088 3065 1152
rect 3129 1088 3145 1152
rect 3018 1072 3145 1088
rect 3018 1008 3065 1072
rect 3129 1008 3145 1072
rect 3018 992 3145 1008
rect 3018 928 3065 992
rect 3129 928 3145 992
rect 3018 912 3145 928
rect 3018 848 3065 912
rect 3129 848 3145 912
rect 3018 832 3145 848
rect 3018 768 3065 832
rect 3129 768 3145 832
rect 3018 752 3145 768
rect 3018 688 3065 752
rect 3129 688 3145 752
rect 3018 672 3145 688
rect 3018 608 3065 672
rect 3129 608 3145 672
rect 3018 592 3145 608
rect 3018 528 3065 592
rect 3129 528 3145 592
rect 3018 512 3145 528
rect 3018 448 3065 512
rect 3129 448 3145 512
rect 3018 432 3145 448
rect 3018 368 3065 432
rect 3129 368 3145 432
rect 3018 352 3145 368
rect 3018 288 3065 352
rect 3129 288 3145 352
rect 3018 272 3145 288
rect 3018 208 3065 272
rect 3129 208 3145 272
rect 3018 192 3145 208
rect 3018 128 3065 192
rect 3129 128 3145 192
rect 3018 112 3145 128
rect 3018 48 3065 112
rect 3129 48 3145 112
rect 3018 32 3145 48
rect 3018 -32 3065 32
rect 3129 -32 3145 32
rect 3018 -48 3145 -32
rect 3018 -112 3065 -48
rect 3129 -112 3145 -48
rect 3018 -128 3145 -112
rect 3018 -192 3065 -128
rect 3129 -192 3145 -128
rect 3018 -208 3145 -192
rect 3018 -272 3065 -208
rect 3129 -272 3145 -208
rect 3018 -288 3145 -272
rect 3018 -352 3065 -288
rect 3129 -352 3145 -288
rect 3018 -368 3145 -352
rect 3018 -432 3065 -368
rect 3129 -432 3145 -368
rect 3018 -448 3145 -432
rect 3018 -512 3065 -448
rect 3129 -512 3145 -448
rect 3018 -528 3145 -512
rect 3018 -592 3065 -528
rect 3129 -592 3145 -528
rect 3018 -608 3145 -592
rect 3018 -672 3065 -608
rect 3129 -672 3145 -608
rect 3018 -688 3145 -672
rect 3018 -752 3065 -688
rect 3129 -752 3145 -688
rect 3018 -768 3145 -752
rect 3018 -832 3065 -768
rect 3129 -832 3145 -768
rect 3018 -848 3145 -832
rect 3018 -912 3065 -848
rect 3129 -912 3145 -848
rect 3018 -928 3145 -912
rect 3018 -992 3065 -928
rect 3129 -992 3145 -928
rect 3018 -1008 3145 -992
rect 3018 -1072 3065 -1008
rect 3129 -1072 3145 -1008
rect 3018 -1088 3145 -1072
rect 3018 -1152 3065 -1088
rect 3129 -1152 3145 -1088
rect 3018 -1168 3145 -1152
rect 3018 -1232 3065 -1168
rect 3129 -1232 3145 -1168
rect 3018 -1248 3145 -1232
rect 3018 -1312 3065 -1248
rect 3129 -1312 3145 -1248
rect 3018 -1328 3145 -1312
rect 3018 -1392 3065 -1328
rect 3129 -1392 3145 -1328
rect 3018 -1408 3145 -1392
rect 3018 -1472 3065 -1408
rect 3129 -1472 3145 -1408
rect 3018 -1488 3145 -1472
rect 3018 -1552 3065 -1488
rect 3129 -1552 3145 -1488
rect 3018 -1568 3145 -1552
rect 3018 -1632 3065 -1568
rect 3129 -1632 3145 -1568
rect 3018 -1648 3145 -1632
rect 3018 -1712 3065 -1648
rect 3129 -1712 3145 -1648
rect 3018 -1728 3145 -1712
rect 3018 -1792 3065 -1728
rect 3129 -1792 3145 -1728
rect 3018 -1808 3145 -1792
rect 3018 -1872 3065 -1808
rect 3129 -1872 3145 -1808
rect 3018 -1888 3145 -1872
rect 3018 -1952 3065 -1888
rect 3129 -1952 3145 -1888
rect 3018 -1968 3145 -1952
rect 3018 -2032 3065 -1968
rect 3129 -2032 3145 -1968
rect 3018 -2048 3145 -2032
rect 3018 -2112 3065 -2048
rect 3129 -2112 3145 -2048
rect 3018 -2128 3145 -2112
rect 3018 -2192 3065 -2128
rect 3129 -2192 3145 -2128
rect 3018 -2208 3145 -2192
rect 3018 -2272 3065 -2208
rect 3129 -2272 3145 -2208
rect 3018 -2288 3145 -2272
rect 3018 -2352 3065 -2288
rect 3129 -2352 3145 -2288
rect 3018 -2368 3145 -2352
rect 3018 -2432 3065 -2368
rect 3129 -2432 3145 -2368
rect 3018 -2448 3145 -2432
rect 3018 -2512 3065 -2448
rect 3129 -2512 3145 -2448
rect 3018 -2528 3145 -2512
rect 3018 -2592 3065 -2528
rect 3129 -2592 3145 -2528
rect 3018 -2608 3145 -2592
rect 3018 -2672 3065 -2608
rect 3129 -2672 3145 -2608
rect 3018 -2688 3145 -2672
rect 3018 -2752 3065 -2688
rect 3129 -2752 3145 -2688
rect 3018 -2768 3145 -2752
rect 3018 -2832 3065 -2768
rect 3129 -2832 3145 -2768
rect 3018 -2848 3145 -2832
rect 3018 -2912 3065 -2848
rect 3129 -2912 3145 -2848
rect 3018 -2928 3145 -2912
rect -3301 -3008 -3174 -2992
rect -3301 -3072 -3254 -3008
rect -3190 -3072 -3174 -3008
rect -3301 -3088 -3174 -3072
rect -3301 -3212 -3197 -3088
rect -3301 -3228 -3174 -3212
rect -3301 -3292 -3254 -3228
rect -3190 -3292 -3174 -3228
rect -3301 -3308 -3174 -3292
rect -9620 -3388 -9493 -3372
rect -9620 -3452 -9573 -3388
rect -9509 -3452 -9493 -3388
rect -9620 -3468 -9493 -3452
rect -9620 -3532 -9573 -3468
rect -9509 -3532 -9493 -3468
rect -9620 -3548 -9493 -3532
rect -9620 -3612 -9573 -3548
rect -9509 -3612 -9493 -3548
rect -9620 -3628 -9493 -3612
rect -9620 -3692 -9573 -3628
rect -9509 -3692 -9493 -3628
rect -9620 -3708 -9493 -3692
rect -9620 -3772 -9573 -3708
rect -9509 -3772 -9493 -3708
rect -9620 -3788 -9493 -3772
rect -9620 -3852 -9573 -3788
rect -9509 -3852 -9493 -3788
rect -9620 -3868 -9493 -3852
rect -9620 -3932 -9573 -3868
rect -9509 -3932 -9493 -3868
rect -9620 -3948 -9493 -3932
rect -9620 -4012 -9573 -3948
rect -9509 -4012 -9493 -3948
rect -9620 -4028 -9493 -4012
rect -9620 -4092 -9573 -4028
rect -9509 -4092 -9493 -4028
rect -9620 -4108 -9493 -4092
rect -9620 -4172 -9573 -4108
rect -9509 -4172 -9493 -4108
rect -9620 -4188 -9493 -4172
rect -9620 -4252 -9573 -4188
rect -9509 -4252 -9493 -4188
rect -9620 -4268 -9493 -4252
rect -9620 -4332 -9573 -4268
rect -9509 -4332 -9493 -4268
rect -9620 -4348 -9493 -4332
rect -9620 -4412 -9573 -4348
rect -9509 -4412 -9493 -4348
rect -9620 -4428 -9493 -4412
rect -9620 -4492 -9573 -4428
rect -9509 -4492 -9493 -4428
rect -9620 -4508 -9493 -4492
rect -9620 -4572 -9573 -4508
rect -9509 -4572 -9493 -4508
rect -9620 -4588 -9493 -4572
rect -9620 -4652 -9573 -4588
rect -9509 -4652 -9493 -4588
rect -9620 -4668 -9493 -4652
rect -9620 -4732 -9573 -4668
rect -9509 -4732 -9493 -4668
rect -9620 -4748 -9493 -4732
rect -9620 -4812 -9573 -4748
rect -9509 -4812 -9493 -4748
rect -9620 -4828 -9493 -4812
rect -9620 -4892 -9573 -4828
rect -9509 -4892 -9493 -4828
rect -9620 -4908 -9493 -4892
rect -9620 -4972 -9573 -4908
rect -9509 -4972 -9493 -4908
rect -9620 -4988 -9493 -4972
rect -9620 -5052 -9573 -4988
rect -9509 -5052 -9493 -4988
rect -9620 -5068 -9493 -5052
rect -9620 -5132 -9573 -5068
rect -9509 -5132 -9493 -5068
rect -9620 -5148 -9493 -5132
rect -9620 -5212 -9573 -5148
rect -9509 -5212 -9493 -5148
rect -9620 -5228 -9493 -5212
rect -9620 -5292 -9573 -5228
rect -9509 -5292 -9493 -5228
rect -9620 -5308 -9493 -5292
rect -9620 -5372 -9573 -5308
rect -9509 -5372 -9493 -5308
rect -9620 -5388 -9493 -5372
rect -9620 -5452 -9573 -5388
rect -9509 -5452 -9493 -5388
rect -9620 -5468 -9493 -5452
rect -9620 -5532 -9573 -5468
rect -9509 -5532 -9493 -5468
rect -9620 -5548 -9493 -5532
rect -9620 -5612 -9573 -5548
rect -9509 -5612 -9493 -5548
rect -9620 -5628 -9493 -5612
rect -9620 -5692 -9573 -5628
rect -9509 -5692 -9493 -5628
rect -9620 -5708 -9493 -5692
rect -9620 -5772 -9573 -5708
rect -9509 -5772 -9493 -5708
rect -9620 -5788 -9493 -5772
rect -9620 -5852 -9573 -5788
rect -9509 -5852 -9493 -5788
rect -9620 -5868 -9493 -5852
rect -9620 -5932 -9573 -5868
rect -9509 -5932 -9493 -5868
rect -9620 -5948 -9493 -5932
rect -9620 -6012 -9573 -5948
rect -9509 -6012 -9493 -5948
rect -9620 -6028 -9493 -6012
rect -9620 -6092 -9573 -6028
rect -9509 -6092 -9493 -6028
rect -9620 -6108 -9493 -6092
rect -9620 -6172 -9573 -6108
rect -9509 -6172 -9493 -6108
rect -9620 -6188 -9493 -6172
rect -9620 -6252 -9573 -6188
rect -9509 -6252 -9493 -6188
rect -9620 -6268 -9493 -6252
rect -9620 -6332 -9573 -6268
rect -9509 -6332 -9493 -6268
rect -9620 -6348 -9493 -6332
rect -9620 -6412 -9573 -6348
rect -9509 -6412 -9493 -6348
rect -9620 -6428 -9493 -6412
rect -9620 -6492 -9573 -6428
rect -9509 -6492 -9493 -6428
rect -9620 -6508 -9493 -6492
rect -9620 -6572 -9573 -6508
rect -9509 -6572 -9493 -6508
rect -9620 -6588 -9493 -6572
rect -9620 -6652 -9573 -6588
rect -9509 -6652 -9493 -6588
rect -9620 -6668 -9493 -6652
rect -9620 -6732 -9573 -6668
rect -9509 -6732 -9493 -6668
rect -9620 -6748 -9493 -6732
rect -9620 -6812 -9573 -6748
rect -9509 -6812 -9493 -6748
rect -9620 -6828 -9493 -6812
rect -9620 -6892 -9573 -6828
rect -9509 -6892 -9493 -6828
rect -9620 -6908 -9493 -6892
rect -9620 -6972 -9573 -6908
rect -9509 -6972 -9493 -6908
rect -9620 -6988 -9493 -6972
rect -9620 -7052 -9573 -6988
rect -9509 -7052 -9493 -6988
rect -9620 -7068 -9493 -7052
rect -9620 -7132 -9573 -7068
rect -9509 -7132 -9493 -7068
rect -9620 -7148 -9493 -7132
rect -9620 -7212 -9573 -7148
rect -9509 -7212 -9493 -7148
rect -9620 -7228 -9493 -7212
rect -9620 -7292 -9573 -7228
rect -9509 -7292 -9493 -7228
rect -9620 -7308 -9493 -7292
rect -9620 -7372 -9573 -7308
rect -9509 -7372 -9493 -7308
rect -9620 -7388 -9493 -7372
rect -9620 -7452 -9573 -7388
rect -9509 -7452 -9493 -7388
rect -9620 -7468 -9493 -7452
rect -9620 -7532 -9573 -7468
rect -9509 -7532 -9493 -7468
rect -9620 -7548 -9493 -7532
rect -9620 -7612 -9573 -7548
rect -9509 -7612 -9493 -7548
rect -9620 -7628 -9493 -7612
rect -9620 -7692 -9573 -7628
rect -9509 -7692 -9493 -7628
rect -9620 -7708 -9493 -7692
rect -9620 -7772 -9573 -7708
rect -9509 -7772 -9493 -7708
rect -9620 -7788 -9493 -7772
rect -9620 -7852 -9573 -7788
rect -9509 -7852 -9493 -7788
rect -9620 -7868 -9493 -7852
rect -9620 -7932 -9573 -7868
rect -9509 -7932 -9493 -7868
rect -9620 -7948 -9493 -7932
rect -9620 -8012 -9573 -7948
rect -9509 -8012 -9493 -7948
rect -9620 -8028 -9493 -8012
rect -9620 -8092 -9573 -8028
rect -9509 -8092 -9493 -8028
rect -9620 -8108 -9493 -8092
rect -9620 -8172 -9573 -8108
rect -9509 -8172 -9493 -8108
rect -9620 -8188 -9493 -8172
rect -9620 -8252 -9573 -8188
rect -9509 -8252 -9493 -8188
rect -9620 -8268 -9493 -8252
rect -9620 -8332 -9573 -8268
rect -9509 -8332 -9493 -8268
rect -9620 -8348 -9493 -8332
rect -9620 -8412 -9573 -8348
rect -9509 -8412 -9493 -8348
rect -9620 -8428 -9493 -8412
rect -9620 -8492 -9573 -8428
rect -9509 -8492 -9493 -8428
rect -9620 -8508 -9493 -8492
rect -9620 -8572 -9573 -8508
rect -9509 -8572 -9493 -8508
rect -9620 -8588 -9493 -8572
rect -9620 -8652 -9573 -8588
rect -9509 -8652 -9493 -8588
rect -9620 -8668 -9493 -8652
rect -9620 -8732 -9573 -8668
rect -9509 -8732 -9493 -8668
rect -9620 -8748 -9493 -8732
rect -9620 -8812 -9573 -8748
rect -9509 -8812 -9493 -8748
rect -9620 -8828 -9493 -8812
rect -9620 -8892 -9573 -8828
rect -9509 -8892 -9493 -8828
rect -9620 -8908 -9493 -8892
rect -9620 -8972 -9573 -8908
rect -9509 -8972 -9493 -8908
rect -9620 -8988 -9493 -8972
rect -9620 -9052 -9573 -8988
rect -9509 -9052 -9493 -8988
rect -9620 -9068 -9493 -9052
rect -9620 -9132 -9573 -9068
rect -9509 -9132 -9493 -9068
rect -9620 -9148 -9493 -9132
rect -9620 -9212 -9573 -9148
rect -9509 -9212 -9493 -9148
rect -9620 -9228 -9493 -9212
rect -15939 -9308 -15812 -9292
rect -15939 -9372 -15892 -9308
rect -15828 -9372 -15812 -9308
rect -15939 -9388 -15812 -9372
rect -15939 -9512 -15835 -9388
rect -15939 -9528 -15812 -9512
rect -15939 -9592 -15892 -9528
rect -15828 -9592 -15812 -9528
rect -15939 -9608 -15812 -9592
rect -22258 -9688 -22131 -9672
rect -22258 -9752 -22211 -9688
rect -22147 -9752 -22131 -9688
rect -22258 -9768 -22131 -9752
rect -22258 -9832 -22211 -9768
rect -22147 -9832 -22131 -9768
rect -22258 -9848 -22131 -9832
rect -22258 -9912 -22211 -9848
rect -22147 -9912 -22131 -9848
rect -22258 -9928 -22131 -9912
rect -22258 -9992 -22211 -9928
rect -22147 -9992 -22131 -9928
rect -22258 -10008 -22131 -9992
rect -22258 -10072 -22211 -10008
rect -22147 -10072 -22131 -10008
rect -22258 -10088 -22131 -10072
rect -22258 -10152 -22211 -10088
rect -22147 -10152 -22131 -10088
rect -22258 -10168 -22131 -10152
rect -22258 -10232 -22211 -10168
rect -22147 -10232 -22131 -10168
rect -22258 -10248 -22131 -10232
rect -22258 -10312 -22211 -10248
rect -22147 -10312 -22131 -10248
rect -22258 -10328 -22131 -10312
rect -22258 -10392 -22211 -10328
rect -22147 -10392 -22131 -10328
rect -22258 -10408 -22131 -10392
rect -22258 -10472 -22211 -10408
rect -22147 -10472 -22131 -10408
rect -22258 -10488 -22131 -10472
rect -22258 -10552 -22211 -10488
rect -22147 -10552 -22131 -10488
rect -22258 -10568 -22131 -10552
rect -22258 -10632 -22211 -10568
rect -22147 -10632 -22131 -10568
rect -22258 -10648 -22131 -10632
rect -22258 -10712 -22211 -10648
rect -22147 -10712 -22131 -10648
rect -22258 -10728 -22131 -10712
rect -22258 -10792 -22211 -10728
rect -22147 -10792 -22131 -10728
rect -22258 -10808 -22131 -10792
rect -22258 -10872 -22211 -10808
rect -22147 -10872 -22131 -10808
rect -22258 -10888 -22131 -10872
rect -22258 -10952 -22211 -10888
rect -22147 -10952 -22131 -10888
rect -22258 -10968 -22131 -10952
rect -22258 -11032 -22211 -10968
rect -22147 -11032 -22131 -10968
rect -22258 -11048 -22131 -11032
rect -22258 -11112 -22211 -11048
rect -22147 -11112 -22131 -11048
rect -22258 -11128 -22131 -11112
rect -22258 -11192 -22211 -11128
rect -22147 -11192 -22131 -11128
rect -22258 -11208 -22131 -11192
rect -22258 -11272 -22211 -11208
rect -22147 -11272 -22131 -11208
rect -22258 -11288 -22131 -11272
rect -22258 -11352 -22211 -11288
rect -22147 -11352 -22131 -11288
rect -22258 -11368 -22131 -11352
rect -22258 -11432 -22211 -11368
rect -22147 -11432 -22131 -11368
rect -22258 -11448 -22131 -11432
rect -22258 -11512 -22211 -11448
rect -22147 -11512 -22131 -11448
rect -22258 -11528 -22131 -11512
rect -22258 -11592 -22211 -11528
rect -22147 -11592 -22131 -11528
rect -22258 -11608 -22131 -11592
rect -22258 -11672 -22211 -11608
rect -22147 -11672 -22131 -11608
rect -22258 -11688 -22131 -11672
rect -22258 -11752 -22211 -11688
rect -22147 -11752 -22131 -11688
rect -22258 -11768 -22131 -11752
rect -22258 -11832 -22211 -11768
rect -22147 -11832 -22131 -11768
rect -22258 -11848 -22131 -11832
rect -22258 -11912 -22211 -11848
rect -22147 -11912 -22131 -11848
rect -22258 -11928 -22131 -11912
rect -22258 -11992 -22211 -11928
rect -22147 -11992 -22131 -11928
rect -22258 -12008 -22131 -11992
rect -22258 -12072 -22211 -12008
rect -22147 -12072 -22131 -12008
rect -22258 -12088 -22131 -12072
rect -22258 -12152 -22211 -12088
rect -22147 -12152 -22131 -12088
rect -22258 -12168 -22131 -12152
rect -22258 -12232 -22211 -12168
rect -22147 -12232 -22131 -12168
rect -22258 -12248 -22131 -12232
rect -22258 -12312 -22211 -12248
rect -22147 -12312 -22131 -12248
rect -22258 -12328 -22131 -12312
rect -22258 -12392 -22211 -12328
rect -22147 -12392 -22131 -12328
rect -22258 -12408 -22131 -12392
rect -22258 -12472 -22211 -12408
rect -22147 -12472 -22131 -12408
rect -22258 -12488 -22131 -12472
rect -22258 -12552 -22211 -12488
rect -22147 -12552 -22131 -12488
rect -22258 -12568 -22131 -12552
rect -22258 -12632 -22211 -12568
rect -22147 -12632 -22131 -12568
rect -22258 -12648 -22131 -12632
rect -22258 -12712 -22211 -12648
rect -22147 -12712 -22131 -12648
rect -22258 -12728 -22131 -12712
rect -22258 -12792 -22211 -12728
rect -22147 -12792 -22131 -12728
rect -22258 -12808 -22131 -12792
rect -22258 -12872 -22211 -12808
rect -22147 -12872 -22131 -12808
rect -22258 -12888 -22131 -12872
rect -22258 -12952 -22211 -12888
rect -22147 -12952 -22131 -12888
rect -22258 -12968 -22131 -12952
rect -22258 -13032 -22211 -12968
rect -22147 -13032 -22131 -12968
rect -22258 -13048 -22131 -13032
rect -22258 -13112 -22211 -13048
rect -22147 -13112 -22131 -13048
rect -22258 -13128 -22131 -13112
rect -22258 -13192 -22211 -13128
rect -22147 -13192 -22131 -13128
rect -22258 -13208 -22131 -13192
rect -22258 -13272 -22211 -13208
rect -22147 -13272 -22131 -13208
rect -22258 -13288 -22131 -13272
rect -22258 -13352 -22211 -13288
rect -22147 -13352 -22131 -13288
rect -22258 -13368 -22131 -13352
rect -22258 -13432 -22211 -13368
rect -22147 -13432 -22131 -13368
rect -22258 -13448 -22131 -13432
rect -22258 -13512 -22211 -13448
rect -22147 -13512 -22131 -13448
rect -22258 -13528 -22131 -13512
rect -22258 -13592 -22211 -13528
rect -22147 -13592 -22131 -13528
rect -22258 -13608 -22131 -13592
rect -22258 -13672 -22211 -13608
rect -22147 -13672 -22131 -13608
rect -22258 -13688 -22131 -13672
rect -22258 -13752 -22211 -13688
rect -22147 -13752 -22131 -13688
rect -22258 -13768 -22131 -13752
rect -22258 -13832 -22211 -13768
rect -22147 -13832 -22131 -13768
rect -22258 -13848 -22131 -13832
rect -22258 -13912 -22211 -13848
rect -22147 -13912 -22131 -13848
rect -22258 -13928 -22131 -13912
rect -22258 -13992 -22211 -13928
rect -22147 -13992 -22131 -13928
rect -22258 -14008 -22131 -13992
rect -22258 -14072 -22211 -14008
rect -22147 -14072 -22131 -14008
rect -22258 -14088 -22131 -14072
rect -22258 -14152 -22211 -14088
rect -22147 -14152 -22131 -14088
rect -22258 -14168 -22131 -14152
rect -22258 -14232 -22211 -14168
rect -22147 -14232 -22131 -14168
rect -22258 -14248 -22131 -14232
rect -22258 -14312 -22211 -14248
rect -22147 -14312 -22131 -14248
rect -22258 -14328 -22131 -14312
rect -22258 -14392 -22211 -14328
rect -22147 -14392 -22131 -14328
rect -22258 -14408 -22131 -14392
rect -22258 -14472 -22211 -14408
rect -22147 -14472 -22131 -14408
rect -22258 -14488 -22131 -14472
rect -22258 -14552 -22211 -14488
rect -22147 -14552 -22131 -14488
rect -22258 -14568 -22131 -14552
rect -22258 -14632 -22211 -14568
rect -22147 -14632 -22131 -14568
rect -22258 -14648 -22131 -14632
rect -22258 -14712 -22211 -14648
rect -22147 -14712 -22131 -14648
rect -22258 -14728 -22131 -14712
rect -22258 -14792 -22211 -14728
rect -22147 -14792 -22131 -14728
rect -22258 -14808 -22131 -14792
rect -22258 -14872 -22211 -14808
rect -22147 -14872 -22131 -14808
rect -22258 -14888 -22131 -14872
rect -22258 -14952 -22211 -14888
rect -22147 -14952 -22131 -14888
rect -22258 -14968 -22131 -14952
rect -22258 -15032 -22211 -14968
rect -22147 -15032 -22131 -14968
rect -22258 -15048 -22131 -15032
rect -22258 -15112 -22211 -15048
rect -22147 -15112 -22131 -15048
rect -22258 -15128 -22131 -15112
rect -22258 -15192 -22211 -15128
rect -22147 -15192 -22131 -15128
rect -22258 -15208 -22131 -15192
rect -22258 -15272 -22211 -15208
rect -22147 -15272 -22131 -15208
rect -22258 -15288 -22131 -15272
rect -22258 -15352 -22211 -15288
rect -22147 -15352 -22131 -15288
rect -22258 -15368 -22131 -15352
rect -22258 -15432 -22211 -15368
rect -22147 -15432 -22131 -15368
rect -22258 -15448 -22131 -15432
rect -22258 -15512 -22211 -15448
rect -22147 -15512 -22131 -15448
rect -22258 -15528 -22131 -15512
rect -28577 -15608 -28450 -15592
rect -28577 -15672 -28530 -15608
rect -28466 -15672 -28450 -15608
rect -28577 -15688 -28450 -15672
rect -28577 -15812 -28473 -15688
rect -28577 -15828 -28450 -15812
rect -28577 -15892 -28530 -15828
rect -28466 -15892 -28450 -15828
rect -28577 -15908 -28450 -15892
rect -34896 -15988 -34769 -15972
rect -34896 -16052 -34849 -15988
rect -34785 -16052 -34769 -15988
rect -34896 -16068 -34769 -16052
rect -34896 -16132 -34849 -16068
rect -34785 -16132 -34769 -16068
rect -34896 -16148 -34769 -16132
rect -34896 -16212 -34849 -16148
rect -34785 -16212 -34769 -16148
rect -34896 -16228 -34769 -16212
rect -34896 -16292 -34849 -16228
rect -34785 -16292 -34769 -16228
rect -34896 -16308 -34769 -16292
rect -34896 -16372 -34849 -16308
rect -34785 -16372 -34769 -16308
rect -34896 -16388 -34769 -16372
rect -34896 -16452 -34849 -16388
rect -34785 -16452 -34769 -16388
rect -34896 -16468 -34769 -16452
rect -34896 -16532 -34849 -16468
rect -34785 -16532 -34769 -16468
rect -34896 -16548 -34769 -16532
rect -34896 -16612 -34849 -16548
rect -34785 -16612 -34769 -16548
rect -34896 -16628 -34769 -16612
rect -34896 -16692 -34849 -16628
rect -34785 -16692 -34769 -16628
rect -34896 -16708 -34769 -16692
rect -34896 -16772 -34849 -16708
rect -34785 -16772 -34769 -16708
rect -34896 -16788 -34769 -16772
rect -34896 -16852 -34849 -16788
rect -34785 -16852 -34769 -16788
rect -34896 -16868 -34769 -16852
rect -34896 -16932 -34849 -16868
rect -34785 -16932 -34769 -16868
rect -34896 -16948 -34769 -16932
rect -34896 -17012 -34849 -16948
rect -34785 -17012 -34769 -16948
rect -34896 -17028 -34769 -17012
rect -34896 -17092 -34849 -17028
rect -34785 -17092 -34769 -17028
rect -34896 -17108 -34769 -17092
rect -34896 -17172 -34849 -17108
rect -34785 -17172 -34769 -17108
rect -34896 -17188 -34769 -17172
rect -34896 -17252 -34849 -17188
rect -34785 -17252 -34769 -17188
rect -34896 -17268 -34769 -17252
rect -34896 -17332 -34849 -17268
rect -34785 -17332 -34769 -17268
rect -34896 -17348 -34769 -17332
rect -34896 -17412 -34849 -17348
rect -34785 -17412 -34769 -17348
rect -34896 -17428 -34769 -17412
rect -34896 -17492 -34849 -17428
rect -34785 -17492 -34769 -17428
rect -34896 -17508 -34769 -17492
rect -34896 -17572 -34849 -17508
rect -34785 -17572 -34769 -17508
rect -34896 -17588 -34769 -17572
rect -34896 -17652 -34849 -17588
rect -34785 -17652 -34769 -17588
rect -34896 -17668 -34769 -17652
rect -34896 -17732 -34849 -17668
rect -34785 -17732 -34769 -17668
rect -34896 -17748 -34769 -17732
rect -34896 -17812 -34849 -17748
rect -34785 -17812 -34769 -17748
rect -34896 -17828 -34769 -17812
rect -34896 -17892 -34849 -17828
rect -34785 -17892 -34769 -17828
rect -34896 -17908 -34769 -17892
rect -34896 -17972 -34849 -17908
rect -34785 -17972 -34769 -17908
rect -34896 -17988 -34769 -17972
rect -34896 -18052 -34849 -17988
rect -34785 -18052 -34769 -17988
rect -34896 -18068 -34769 -18052
rect -34896 -18132 -34849 -18068
rect -34785 -18132 -34769 -18068
rect -34896 -18148 -34769 -18132
rect -34896 -18212 -34849 -18148
rect -34785 -18212 -34769 -18148
rect -34896 -18228 -34769 -18212
rect -34896 -18292 -34849 -18228
rect -34785 -18292 -34769 -18228
rect -34896 -18308 -34769 -18292
rect -34896 -18372 -34849 -18308
rect -34785 -18372 -34769 -18308
rect -34896 -18388 -34769 -18372
rect -34896 -18452 -34849 -18388
rect -34785 -18452 -34769 -18388
rect -34896 -18468 -34769 -18452
rect -34896 -18532 -34849 -18468
rect -34785 -18532 -34769 -18468
rect -34896 -18548 -34769 -18532
rect -34896 -18612 -34849 -18548
rect -34785 -18612 -34769 -18548
rect -34896 -18628 -34769 -18612
rect -34896 -18692 -34849 -18628
rect -34785 -18692 -34769 -18628
rect -34896 -18708 -34769 -18692
rect -34896 -18772 -34849 -18708
rect -34785 -18772 -34769 -18708
rect -34896 -18788 -34769 -18772
rect -34896 -18852 -34849 -18788
rect -34785 -18852 -34769 -18788
rect -34896 -18868 -34769 -18852
rect -34896 -18932 -34849 -18868
rect -34785 -18932 -34769 -18868
rect -34896 -18948 -34769 -18932
rect -34896 -19012 -34849 -18948
rect -34785 -19012 -34769 -18948
rect -34896 -19028 -34769 -19012
rect -34896 -19092 -34849 -19028
rect -34785 -19092 -34769 -19028
rect -34896 -19108 -34769 -19092
rect -34896 -19172 -34849 -19108
rect -34785 -19172 -34769 -19108
rect -34896 -19188 -34769 -19172
rect -34896 -19252 -34849 -19188
rect -34785 -19252 -34769 -19188
rect -34896 -19268 -34769 -19252
rect -34896 -19332 -34849 -19268
rect -34785 -19332 -34769 -19268
rect -34896 -19348 -34769 -19332
rect -34896 -19412 -34849 -19348
rect -34785 -19412 -34769 -19348
rect -34896 -19428 -34769 -19412
rect -34896 -19492 -34849 -19428
rect -34785 -19492 -34769 -19428
rect -34896 -19508 -34769 -19492
rect -34896 -19572 -34849 -19508
rect -34785 -19572 -34769 -19508
rect -34896 -19588 -34769 -19572
rect -34896 -19652 -34849 -19588
rect -34785 -19652 -34769 -19588
rect -34896 -19668 -34769 -19652
rect -34896 -19732 -34849 -19668
rect -34785 -19732 -34769 -19668
rect -34896 -19748 -34769 -19732
rect -34896 -19812 -34849 -19748
rect -34785 -19812 -34769 -19748
rect -34896 -19828 -34769 -19812
rect -34896 -19892 -34849 -19828
rect -34785 -19892 -34769 -19828
rect -34896 -19908 -34769 -19892
rect -34896 -19972 -34849 -19908
rect -34785 -19972 -34769 -19908
rect -34896 -19988 -34769 -19972
rect -34896 -20052 -34849 -19988
rect -34785 -20052 -34769 -19988
rect -34896 -20068 -34769 -20052
rect -34896 -20132 -34849 -20068
rect -34785 -20132 -34769 -20068
rect -34896 -20148 -34769 -20132
rect -34896 -20212 -34849 -20148
rect -34785 -20212 -34769 -20148
rect -34896 -20228 -34769 -20212
rect -34896 -20292 -34849 -20228
rect -34785 -20292 -34769 -20228
rect -34896 -20308 -34769 -20292
rect -34896 -20372 -34849 -20308
rect -34785 -20372 -34769 -20308
rect -34896 -20388 -34769 -20372
rect -34896 -20452 -34849 -20388
rect -34785 -20452 -34769 -20388
rect -34896 -20468 -34769 -20452
rect -34896 -20532 -34849 -20468
rect -34785 -20532 -34769 -20468
rect -34896 -20548 -34769 -20532
rect -34896 -20612 -34849 -20548
rect -34785 -20612 -34769 -20548
rect -34896 -20628 -34769 -20612
rect -34896 -20692 -34849 -20628
rect -34785 -20692 -34769 -20628
rect -34896 -20708 -34769 -20692
rect -34896 -20772 -34849 -20708
rect -34785 -20772 -34769 -20708
rect -34896 -20788 -34769 -20772
rect -34896 -20852 -34849 -20788
rect -34785 -20852 -34769 -20788
rect -34896 -20868 -34769 -20852
rect -34896 -20932 -34849 -20868
rect -34785 -20932 -34769 -20868
rect -34896 -20948 -34769 -20932
rect -34896 -21012 -34849 -20948
rect -34785 -21012 -34769 -20948
rect -34896 -21028 -34769 -21012
rect -34896 -21092 -34849 -21028
rect -34785 -21092 -34769 -21028
rect -34896 -21108 -34769 -21092
rect -34896 -21172 -34849 -21108
rect -34785 -21172 -34769 -21108
rect -34896 -21188 -34769 -21172
rect -34896 -21252 -34849 -21188
rect -34785 -21252 -34769 -21188
rect -34896 -21268 -34769 -21252
rect -34896 -21332 -34849 -21268
rect -34785 -21332 -34769 -21268
rect -34896 -21348 -34769 -21332
rect -34896 -21412 -34849 -21348
rect -34785 -21412 -34769 -21348
rect -34896 -21428 -34769 -21412
rect -34896 -21492 -34849 -21428
rect -34785 -21492 -34769 -21428
rect -34896 -21508 -34769 -21492
rect -34896 -21572 -34849 -21508
rect -34785 -21572 -34769 -21508
rect -34896 -21588 -34769 -21572
rect -34896 -21652 -34849 -21588
rect -34785 -21652 -34769 -21588
rect -34896 -21668 -34769 -21652
rect -34896 -21732 -34849 -21668
rect -34785 -21732 -34769 -21668
rect -34896 -21748 -34769 -21732
rect -34896 -21812 -34849 -21748
rect -34785 -21812 -34769 -21748
rect -34896 -21828 -34769 -21812
rect -41215 -21908 -41088 -21892
rect -41215 -21972 -41168 -21908
rect -41104 -21972 -41088 -21908
rect -41215 -21988 -41088 -21972
rect -41215 -22112 -41111 -21988
rect -41215 -22128 -41088 -22112
rect -41215 -22192 -41168 -22128
rect -41104 -22192 -41088 -22128
rect -41215 -22208 -41088 -22192
rect -47244 -22248 -41322 -22239
rect -47244 -28152 -47235 -22248
rect -41331 -28152 -41322 -22248
rect -47244 -28161 -41322 -28152
rect -41215 -22272 -41168 -22208
rect -41104 -22272 -41088 -22208
rect -38016 -22239 -37912 -21861
rect -34896 -21892 -34849 -21828
rect -34785 -21892 -34769 -21828
rect -34606 -15948 -28684 -15939
rect -34606 -21852 -34597 -15948
rect -28693 -21852 -28684 -15948
rect -34606 -21861 -28684 -21852
rect -28577 -15972 -28530 -15908
rect -28466 -15972 -28450 -15908
rect -25378 -15939 -25274 -15561
rect -22258 -15592 -22211 -15528
rect -22147 -15592 -22131 -15528
rect -21968 -9648 -16046 -9639
rect -21968 -15552 -21959 -9648
rect -16055 -15552 -16046 -9648
rect -21968 -15561 -16046 -15552
rect -15939 -9672 -15892 -9608
rect -15828 -9672 -15812 -9608
rect -12740 -9639 -12636 -9261
rect -9620 -9292 -9573 -9228
rect -9509 -9292 -9493 -9228
rect -9330 -3348 -3408 -3339
rect -9330 -9252 -9321 -3348
rect -3417 -9252 -3408 -3348
rect -9330 -9261 -3408 -9252
rect -3301 -3372 -3254 -3308
rect -3190 -3372 -3174 -3308
rect -102 -3339 2 -2961
rect 3018 -2992 3065 -2928
rect 3129 -2992 3145 -2928
rect 3308 2952 9230 2961
rect 3308 -2952 3317 2952
rect 9221 -2952 9230 2952
rect 3308 -2961 9230 -2952
rect 9337 2928 9384 2992
rect 9448 2928 9464 2992
rect 12536 2961 12640 3339
rect 15656 3308 15703 3372
rect 15767 3308 15783 3372
rect 15946 9252 21868 9261
rect 15946 3348 15955 9252
rect 21859 3348 21868 9252
rect 15946 3339 21868 3348
rect 21975 9228 22022 9292
rect 22086 9228 22102 9292
rect 25174 9261 25278 9639
rect 28294 9608 28341 9672
rect 28405 9608 28421 9672
rect 28584 15552 34506 15561
rect 28584 9648 28593 15552
rect 34497 9648 34506 15552
rect 28584 9639 34506 9648
rect 34613 15528 34660 15592
rect 34724 15528 34740 15592
rect 37812 15561 37916 15939
rect 40932 15908 40979 15972
rect 41043 15908 41059 15972
rect 41222 21852 47144 21861
rect 41222 15948 41231 21852
rect 47135 15948 47144 21852
rect 41222 15939 47144 15948
rect 47251 21828 47298 21892
rect 47362 21828 47378 21892
rect 47251 21812 47378 21828
rect 47251 21748 47298 21812
rect 47362 21748 47378 21812
rect 47251 21732 47378 21748
rect 47251 21668 47298 21732
rect 47362 21668 47378 21732
rect 47251 21652 47378 21668
rect 47251 21588 47298 21652
rect 47362 21588 47378 21652
rect 47251 21572 47378 21588
rect 47251 21508 47298 21572
rect 47362 21508 47378 21572
rect 47251 21492 47378 21508
rect 47251 21428 47298 21492
rect 47362 21428 47378 21492
rect 47251 21412 47378 21428
rect 47251 21348 47298 21412
rect 47362 21348 47378 21412
rect 47251 21332 47378 21348
rect 47251 21268 47298 21332
rect 47362 21268 47378 21332
rect 47251 21252 47378 21268
rect 47251 21188 47298 21252
rect 47362 21188 47378 21252
rect 47251 21172 47378 21188
rect 47251 21108 47298 21172
rect 47362 21108 47378 21172
rect 47251 21092 47378 21108
rect 47251 21028 47298 21092
rect 47362 21028 47378 21092
rect 47251 21012 47378 21028
rect 47251 20948 47298 21012
rect 47362 20948 47378 21012
rect 47251 20932 47378 20948
rect 47251 20868 47298 20932
rect 47362 20868 47378 20932
rect 47251 20852 47378 20868
rect 47251 20788 47298 20852
rect 47362 20788 47378 20852
rect 47251 20772 47378 20788
rect 47251 20708 47298 20772
rect 47362 20708 47378 20772
rect 47251 20692 47378 20708
rect 47251 20628 47298 20692
rect 47362 20628 47378 20692
rect 47251 20612 47378 20628
rect 47251 20548 47298 20612
rect 47362 20548 47378 20612
rect 47251 20532 47378 20548
rect 47251 20468 47298 20532
rect 47362 20468 47378 20532
rect 47251 20452 47378 20468
rect 47251 20388 47298 20452
rect 47362 20388 47378 20452
rect 47251 20372 47378 20388
rect 47251 20308 47298 20372
rect 47362 20308 47378 20372
rect 47251 20292 47378 20308
rect 47251 20228 47298 20292
rect 47362 20228 47378 20292
rect 47251 20212 47378 20228
rect 47251 20148 47298 20212
rect 47362 20148 47378 20212
rect 47251 20132 47378 20148
rect 47251 20068 47298 20132
rect 47362 20068 47378 20132
rect 47251 20052 47378 20068
rect 47251 19988 47298 20052
rect 47362 19988 47378 20052
rect 47251 19972 47378 19988
rect 47251 19908 47298 19972
rect 47362 19908 47378 19972
rect 47251 19892 47378 19908
rect 47251 19828 47298 19892
rect 47362 19828 47378 19892
rect 47251 19812 47378 19828
rect 47251 19748 47298 19812
rect 47362 19748 47378 19812
rect 47251 19732 47378 19748
rect 47251 19668 47298 19732
rect 47362 19668 47378 19732
rect 47251 19652 47378 19668
rect 47251 19588 47298 19652
rect 47362 19588 47378 19652
rect 47251 19572 47378 19588
rect 47251 19508 47298 19572
rect 47362 19508 47378 19572
rect 47251 19492 47378 19508
rect 47251 19428 47298 19492
rect 47362 19428 47378 19492
rect 47251 19412 47378 19428
rect 47251 19348 47298 19412
rect 47362 19348 47378 19412
rect 47251 19332 47378 19348
rect 47251 19268 47298 19332
rect 47362 19268 47378 19332
rect 47251 19252 47378 19268
rect 47251 19188 47298 19252
rect 47362 19188 47378 19252
rect 47251 19172 47378 19188
rect 47251 19108 47298 19172
rect 47362 19108 47378 19172
rect 47251 19092 47378 19108
rect 47251 19028 47298 19092
rect 47362 19028 47378 19092
rect 47251 19012 47378 19028
rect 47251 18948 47298 19012
rect 47362 18948 47378 19012
rect 47251 18932 47378 18948
rect 47251 18868 47298 18932
rect 47362 18868 47378 18932
rect 47251 18852 47378 18868
rect 47251 18788 47298 18852
rect 47362 18788 47378 18852
rect 47251 18772 47378 18788
rect 47251 18708 47298 18772
rect 47362 18708 47378 18772
rect 47251 18692 47378 18708
rect 47251 18628 47298 18692
rect 47362 18628 47378 18692
rect 47251 18612 47378 18628
rect 47251 18548 47298 18612
rect 47362 18548 47378 18612
rect 47251 18532 47378 18548
rect 47251 18468 47298 18532
rect 47362 18468 47378 18532
rect 47251 18452 47378 18468
rect 47251 18388 47298 18452
rect 47362 18388 47378 18452
rect 47251 18372 47378 18388
rect 47251 18308 47298 18372
rect 47362 18308 47378 18372
rect 47251 18292 47378 18308
rect 47251 18228 47298 18292
rect 47362 18228 47378 18292
rect 47251 18212 47378 18228
rect 47251 18148 47298 18212
rect 47362 18148 47378 18212
rect 47251 18132 47378 18148
rect 47251 18068 47298 18132
rect 47362 18068 47378 18132
rect 47251 18052 47378 18068
rect 47251 17988 47298 18052
rect 47362 17988 47378 18052
rect 47251 17972 47378 17988
rect 47251 17908 47298 17972
rect 47362 17908 47378 17972
rect 47251 17892 47378 17908
rect 47251 17828 47298 17892
rect 47362 17828 47378 17892
rect 47251 17812 47378 17828
rect 47251 17748 47298 17812
rect 47362 17748 47378 17812
rect 47251 17732 47378 17748
rect 47251 17668 47298 17732
rect 47362 17668 47378 17732
rect 47251 17652 47378 17668
rect 47251 17588 47298 17652
rect 47362 17588 47378 17652
rect 47251 17572 47378 17588
rect 47251 17508 47298 17572
rect 47362 17508 47378 17572
rect 47251 17492 47378 17508
rect 47251 17428 47298 17492
rect 47362 17428 47378 17492
rect 47251 17412 47378 17428
rect 47251 17348 47298 17412
rect 47362 17348 47378 17412
rect 47251 17332 47378 17348
rect 47251 17268 47298 17332
rect 47362 17268 47378 17332
rect 47251 17252 47378 17268
rect 47251 17188 47298 17252
rect 47362 17188 47378 17252
rect 47251 17172 47378 17188
rect 47251 17108 47298 17172
rect 47362 17108 47378 17172
rect 47251 17092 47378 17108
rect 47251 17028 47298 17092
rect 47362 17028 47378 17092
rect 47251 17012 47378 17028
rect 47251 16948 47298 17012
rect 47362 16948 47378 17012
rect 47251 16932 47378 16948
rect 47251 16868 47298 16932
rect 47362 16868 47378 16932
rect 47251 16852 47378 16868
rect 47251 16788 47298 16852
rect 47362 16788 47378 16852
rect 47251 16772 47378 16788
rect 47251 16708 47298 16772
rect 47362 16708 47378 16772
rect 47251 16692 47378 16708
rect 47251 16628 47298 16692
rect 47362 16628 47378 16692
rect 47251 16612 47378 16628
rect 47251 16548 47298 16612
rect 47362 16548 47378 16612
rect 47251 16532 47378 16548
rect 47251 16468 47298 16532
rect 47362 16468 47378 16532
rect 47251 16452 47378 16468
rect 47251 16388 47298 16452
rect 47362 16388 47378 16452
rect 47251 16372 47378 16388
rect 47251 16308 47298 16372
rect 47362 16308 47378 16372
rect 47251 16292 47378 16308
rect 47251 16228 47298 16292
rect 47362 16228 47378 16292
rect 47251 16212 47378 16228
rect 47251 16148 47298 16212
rect 47362 16148 47378 16212
rect 47251 16132 47378 16148
rect 47251 16068 47298 16132
rect 47362 16068 47378 16132
rect 47251 16052 47378 16068
rect 47251 15988 47298 16052
rect 47362 15988 47378 16052
rect 47251 15972 47378 15988
rect 40932 15892 41059 15908
rect 40932 15828 40979 15892
rect 41043 15828 41059 15892
rect 40932 15812 41059 15828
rect 40932 15688 41036 15812
rect 40932 15672 41059 15688
rect 40932 15608 40979 15672
rect 41043 15608 41059 15672
rect 40932 15592 41059 15608
rect 34613 15512 34740 15528
rect 34613 15448 34660 15512
rect 34724 15448 34740 15512
rect 34613 15432 34740 15448
rect 34613 15368 34660 15432
rect 34724 15368 34740 15432
rect 34613 15352 34740 15368
rect 34613 15288 34660 15352
rect 34724 15288 34740 15352
rect 34613 15272 34740 15288
rect 34613 15208 34660 15272
rect 34724 15208 34740 15272
rect 34613 15192 34740 15208
rect 34613 15128 34660 15192
rect 34724 15128 34740 15192
rect 34613 15112 34740 15128
rect 34613 15048 34660 15112
rect 34724 15048 34740 15112
rect 34613 15032 34740 15048
rect 34613 14968 34660 15032
rect 34724 14968 34740 15032
rect 34613 14952 34740 14968
rect 34613 14888 34660 14952
rect 34724 14888 34740 14952
rect 34613 14872 34740 14888
rect 34613 14808 34660 14872
rect 34724 14808 34740 14872
rect 34613 14792 34740 14808
rect 34613 14728 34660 14792
rect 34724 14728 34740 14792
rect 34613 14712 34740 14728
rect 34613 14648 34660 14712
rect 34724 14648 34740 14712
rect 34613 14632 34740 14648
rect 34613 14568 34660 14632
rect 34724 14568 34740 14632
rect 34613 14552 34740 14568
rect 34613 14488 34660 14552
rect 34724 14488 34740 14552
rect 34613 14472 34740 14488
rect 34613 14408 34660 14472
rect 34724 14408 34740 14472
rect 34613 14392 34740 14408
rect 34613 14328 34660 14392
rect 34724 14328 34740 14392
rect 34613 14312 34740 14328
rect 34613 14248 34660 14312
rect 34724 14248 34740 14312
rect 34613 14232 34740 14248
rect 34613 14168 34660 14232
rect 34724 14168 34740 14232
rect 34613 14152 34740 14168
rect 34613 14088 34660 14152
rect 34724 14088 34740 14152
rect 34613 14072 34740 14088
rect 34613 14008 34660 14072
rect 34724 14008 34740 14072
rect 34613 13992 34740 14008
rect 34613 13928 34660 13992
rect 34724 13928 34740 13992
rect 34613 13912 34740 13928
rect 34613 13848 34660 13912
rect 34724 13848 34740 13912
rect 34613 13832 34740 13848
rect 34613 13768 34660 13832
rect 34724 13768 34740 13832
rect 34613 13752 34740 13768
rect 34613 13688 34660 13752
rect 34724 13688 34740 13752
rect 34613 13672 34740 13688
rect 34613 13608 34660 13672
rect 34724 13608 34740 13672
rect 34613 13592 34740 13608
rect 34613 13528 34660 13592
rect 34724 13528 34740 13592
rect 34613 13512 34740 13528
rect 34613 13448 34660 13512
rect 34724 13448 34740 13512
rect 34613 13432 34740 13448
rect 34613 13368 34660 13432
rect 34724 13368 34740 13432
rect 34613 13352 34740 13368
rect 34613 13288 34660 13352
rect 34724 13288 34740 13352
rect 34613 13272 34740 13288
rect 34613 13208 34660 13272
rect 34724 13208 34740 13272
rect 34613 13192 34740 13208
rect 34613 13128 34660 13192
rect 34724 13128 34740 13192
rect 34613 13112 34740 13128
rect 34613 13048 34660 13112
rect 34724 13048 34740 13112
rect 34613 13032 34740 13048
rect 34613 12968 34660 13032
rect 34724 12968 34740 13032
rect 34613 12952 34740 12968
rect 34613 12888 34660 12952
rect 34724 12888 34740 12952
rect 34613 12872 34740 12888
rect 34613 12808 34660 12872
rect 34724 12808 34740 12872
rect 34613 12792 34740 12808
rect 34613 12728 34660 12792
rect 34724 12728 34740 12792
rect 34613 12712 34740 12728
rect 34613 12648 34660 12712
rect 34724 12648 34740 12712
rect 34613 12632 34740 12648
rect 34613 12568 34660 12632
rect 34724 12568 34740 12632
rect 34613 12552 34740 12568
rect 34613 12488 34660 12552
rect 34724 12488 34740 12552
rect 34613 12472 34740 12488
rect 34613 12408 34660 12472
rect 34724 12408 34740 12472
rect 34613 12392 34740 12408
rect 34613 12328 34660 12392
rect 34724 12328 34740 12392
rect 34613 12312 34740 12328
rect 34613 12248 34660 12312
rect 34724 12248 34740 12312
rect 34613 12232 34740 12248
rect 34613 12168 34660 12232
rect 34724 12168 34740 12232
rect 34613 12152 34740 12168
rect 34613 12088 34660 12152
rect 34724 12088 34740 12152
rect 34613 12072 34740 12088
rect 34613 12008 34660 12072
rect 34724 12008 34740 12072
rect 34613 11992 34740 12008
rect 34613 11928 34660 11992
rect 34724 11928 34740 11992
rect 34613 11912 34740 11928
rect 34613 11848 34660 11912
rect 34724 11848 34740 11912
rect 34613 11832 34740 11848
rect 34613 11768 34660 11832
rect 34724 11768 34740 11832
rect 34613 11752 34740 11768
rect 34613 11688 34660 11752
rect 34724 11688 34740 11752
rect 34613 11672 34740 11688
rect 34613 11608 34660 11672
rect 34724 11608 34740 11672
rect 34613 11592 34740 11608
rect 34613 11528 34660 11592
rect 34724 11528 34740 11592
rect 34613 11512 34740 11528
rect 34613 11448 34660 11512
rect 34724 11448 34740 11512
rect 34613 11432 34740 11448
rect 34613 11368 34660 11432
rect 34724 11368 34740 11432
rect 34613 11352 34740 11368
rect 34613 11288 34660 11352
rect 34724 11288 34740 11352
rect 34613 11272 34740 11288
rect 34613 11208 34660 11272
rect 34724 11208 34740 11272
rect 34613 11192 34740 11208
rect 34613 11128 34660 11192
rect 34724 11128 34740 11192
rect 34613 11112 34740 11128
rect 34613 11048 34660 11112
rect 34724 11048 34740 11112
rect 34613 11032 34740 11048
rect 34613 10968 34660 11032
rect 34724 10968 34740 11032
rect 34613 10952 34740 10968
rect 34613 10888 34660 10952
rect 34724 10888 34740 10952
rect 34613 10872 34740 10888
rect 34613 10808 34660 10872
rect 34724 10808 34740 10872
rect 34613 10792 34740 10808
rect 34613 10728 34660 10792
rect 34724 10728 34740 10792
rect 34613 10712 34740 10728
rect 34613 10648 34660 10712
rect 34724 10648 34740 10712
rect 34613 10632 34740 10648
rect 34613 10568 34660 10632
rect 34724 10568 34740 10632
rect 34613 10552 34740 10568
rect 34613 10488 34660 10552
rect 34724 10488 34740 10552
rect 34613 10472 34740 10488
rect 34613 10408 34660 10472
rect 34724 10408 34740 10472
rect 34613 10392 34740 10408
rect 34613 10328 34660 10392
rect 34724 10328 34740 10392
rect 34613 10312 34740 10328
rect 34613 10248 34660 10312
rect 34724 10248 34740 10312
rect 34613 10232 34740 10248
rect 34613 10168 34660 10232
rect 34724 10168 34740 10232
rect 34613 10152 34740 10168
rect 34613 10088 34660 10152
rect 34724 10088 34740 10152
rect 34613 10072 34740 10088
rect 34613 10008 34660 10072
rect 34724 10008 34740 10072
rect 34613 9992 34740 10008
rect 34613 9928 34660 9992
rect 34724 9928 34740 9992
rect 34613 9912 34740 9928
rect 34613 9848 34660 9912
rect 34724 9848 34740 9912
rect 34613 9832 34740 9848
rect 34613 9768 34660 9832
rect 34724 9768 34740 9832
rect 34613 9752 34740 9768
rect 34613 9688 34660 9752
rect 34724 9688 34740 9752
rect 34613 9672 34740 9688
rect 28294 9592 28421 9608
rect 28294 9528 28341 9592
rect 28405 9528 28421 9592
rect 28294 9512 28421 9528
rect 28294 9388 28398 9512
rect 28294 9372 28421 9388
rect 28294 9308 28341 9372
rect 28405 9308 28421 9372
rect 28294 9292 28421 9308
rect 21975 9212 22102 9228
rect 21975 9148 22022 9212
rect 22086 9148 22102 9212
rect 21975 9132 22102 9148
rect 21975 9068 22022 9132
rect 22086 9068 22102 9132
rect 21975 9052 22102 9068
rect 21975 8988 22022 9052
rect 22086 8988 22102 9052
rect 21975 8972 22102 8988
rect 21975 8908 22022 8972
rect 22086 8908 22102 8972
rect 21975 8892 22102 8908
rect 21975 8828 22022 8892
rect 22086 8828 22102 8892
rect 21975 8812 22102 8828
rect 21975 8748 22022 8812
rect 22086 8748 22102 8812
rect 21975 8732 22102 8748
rect 21975 8668 22022 8732
rect 22086 8668 22102 8732
rect 21975 8652 22102 8668
rect 21975 8588 22022 8652
rect 22086 8588 22102 8652
rect 21975 8572 22102 8588
rect 21975 8508 22022 8572
rect 22086 8508 22102 8572
rect 21975 8492 22102 8508
rect 21975 8428 22022 8492
rect 22086 8428 22102 8492
rect 21975 8412 22102 8428
rect 21975 8348 22022 8412
rect 22086 8348 22102 8412
rect 21975 8332 22102 8348
rect 21975 8268 22022 8332
rect 22086 8268 22102 8332
rect 21975 8252 22102 8268
rect 21975 8188 22022 8252
rect 22086 8188 22102 8252
rect 21975 8172 22102 8188
rect 21975 8108 22022 8172
rect 22086 8108 22102 8172
rect 21975 8092 22102 8108
rect 21975 8028 22022 8092
rect 22086 8028 22102 8092
rect 21975 8012 22102 8028
rect 21975 7948 22022 8012
rect 22086 7948 22102 8012
rect 21975 7932 22102 7948
rect 21975 7868 22022 7932
rect 22086 7868 22102 7932
rect 21975 7852 22102 7868
rect 21975 7788 22022 7852
rect 22086 7788 22102 7852
rect 21975 7772 22102 7788
rect 21975 7708 22022 7772
rect 22086 7708 22102 7772
rect 21975 7692 22102 7708
rect 21975 7628 22022 7692
rect 22086 7628 22102 7692
rect 21975 7612 22102 7628
rect 21975 7548 22022 7612
rect 22086 7548 22102 7612
rect 21975 7532 22102 7548
rect 21975 7468 22022 7532
rect 22086 7468 22102 7532
rect 21975 7452 22102 7468
rect 21975 7388 22022 7452
rect 22086 7388 22102 7452
rect 21975 7372 22102 7388
rect 21975 7308 22022 7372
rect 22086 7308 22102 7372
rect 21975 7292 22102 7308
rect 21975 7228 22022 7292
rect 22086 7228 22102 7292
rect 21975 7212 22102 7228
rect 21975 7148 22022 7212
rect 22086 7148 22102 7212
rect 21975 7132 22102 7148
rect 21975 7068 22022 7132
rect 22086 7068 22102 7132
rect 21975 7052 22102 7068
rect 21975 6988 22022 7052
rect 22086 6988 22102 7052
rect 21975 6972 22102 6988
rect 21975 6908 22022 6972
rect 22086 6908 22102 6972
rect 21975 6892 22102 6908
rect 21975 6828 22022 6892
rect 22086 6828 22102 6892
rect 21975 6812 22102 6828
rect 21975 6748 22022 6812
rect 22086 6748 22102 6812
rect 21975 6732 22102 6748
rect 21975 6668 22022 6732
rect 22086 6668 22102 6732
rect 21975 6652 22102 6668
rect 21975 6588 22022 6652
rect 22086 6588 22102 6652
rect 21975 6572 22102 6588
rect 21975 6508 22022 6572
rect 22086 6508 22102 6572
rect 21975 6492 22102 6508
rect 21975 6428 22022 6492
rect 22086 6428 22102 6492
rect 21975 6412 22102 6428
rect 21975 6348 22022 6412
rect 22086 6348 22102 6412
rect 21975 6332 22102 6348
rect 21975 6268 22022 6332
rect 22086 6268 22102 6332
rect 21975 6252 22102 6268
rect 21975 6188 22022 6252
rect 22086 6188 22102 6252
rect 21975 6172 22102 6188
rect 21975 6108 22022 6172
rect 22086 6108 22102 6172
rect 21975 6092 22102 6108
rect 21975 6028 22022 6092
rect 22086 6028 22102 6092
rect 21975 6012 22102 6028
rect 21975 5948 22022 6012
rect 22086 5948 22102 6012
rect 21975 5932 22102 5948
rect 21975 5868 22022 5932
rect 22086 5868 22102 5932
rect 21975 5852 22102 5868
rect 21975 5788 22022 5852
rect 22086 5788 22102 5852
rect 21975 5772 22102 5788
rect 21975 5708 22022 5772
rect 22086 5708 22102 5772
rect 21975 5692 22102 5708
rect 21975 5628 22022 5692
rect 22086 5628 22102 5692
rect 21975 5612 22102 5628
rect 21975 5548 22022 5612
rect 22086 5548 22102 5612
rect 21975 5532 22102 5548
rect 21975 5468 22022 5532
rect 22086 5468 22102 5532
rect 21975 5452 22102 5468
rect 21975 5388 22022 5452
rect 22086 5388 22102 5452
rect 21975 5372 22102 5388
rect 21975 5308 22022 5372
rect 22086 5308 22102 5372
rect 21975 5292 22102 5308
rect 21975 5228 22022 5292
rect 22086 5228 22102 5292
rect 21975 5212 22102 5228
rect 21975 5148 22022 5212
rect 22086 5148 22102 5212
rect 21975 5132 22102 5148
rect 21975 5068 22022 5132
rect 22086 5068 22102 5132
rect 21975 5052 22102 5068
rect 21975 4988 22022 5052
rect 22086 4988 22102 5052
rect 21975 4972 22102 4988
rect 21975 4908 22022 4972
rect 22086 4908 22102 4972
rect 21975 4892 22102 4908
rect 21975 4828 22022 4892
rect 22086 4828 22102 4892
rect 21975 4812 22102 4828
rect 21975 4748 22022 4812
rect 22086 4748 22102 4812
rect 21975 4732 22102 4748
rect 21975 4668 22022 4732
rect 22086 4668 22102 4732
rect 21975 4652 22102 4668
rect 21975 4588 22022 4652
rect 22086 4588 22102 4652
rect 21975 4572 22102 4588
rect 21975 4508 22022 4572
rect 22086 4508 22102 4572
rect 21975 4492 22102 4508
rect 21975 4428 22022 4492
rect 22086 4428 22102 4492
rect 21975 4412 22102 4428
rect 21975 4348 22022 4412
rect 22086 4348 22102 4412
rect 21975 4332 22102 4348
rect 21975 4268 22022 4332
rect 22086 4268 22102 4332
rect 21975 4252 22102 4268
rect 21975 4188 22022 4252
rect 22086 4188 22102 4252
rect 21975 4172 22102 4188
rect 21975 4108 22022 4172
rect 22086 4108 22102 4172
rect 21975 4092 22102 4108
rect 21975 4028 22022 4092
rect 22086 4028 22102 4092
rect 21975 4012 22102 4028
rect 21975 3948 22022 4012
rect 22086 3948 22102 4012
rect 21975 3932 22102 3948
rect 21975 3868 22022 3932
rect 22086 3868 22102 3932
rect 21975 3852 22102 3868
rect 21975 3788 22022 3852
rect 22086 3788 22102 3852
rect 21975 3772 22102 3788
rect 21975 3708 22022 3772
rect 22086 3708 22102 3772
rect 21975 3692 22102 3708
rect 21975 3628 22022 3692
rect 22086 3628 22102 3692
rect 21975 3612 22102 3628
rect 21975 3548 22022 3612
rect 22086 3548 22102 3612
rect 21975 3532 22102 3548
rect 21975 3468 22022 3532
rect 22086 3468 22102 3532
rect 21975 3452 22102 3468
rect 21975 3388 22022 3452
rect 22086 3388 22102 3452
rect 21975 3372 22102 3388
rect 15656 3292 15783 3308
rect 15656 3228 15703 3292
rect 15767 3228 15783 3292
rect 15656 3212 15783 3228
rect 15656 3088 15760 3212
rect 15656 3072 15783 3088
rect 15656 3008 15703 3072
rect 15767 3008 15783 3072
rect 15656 2992 15783 3008
rect 9337 2912 9464 2928
rect 9337 2848 9384 2912
rect 9448 2848 9464 2912
rect 9337 2832 9464 2848
rect 9337 2768 9384 2832
rect 9448 2768 9464 2832
rect 9337 2752 9464 2768
rect 9337 2688 9384 2752
rect 9448 2688 9464 2752
rect 9337 2672 9464 2688
rect 9337 2608 9384 2672
rect 9448 2608 9464 2672
rect 9337 2592 9464 2608
rect 9337 2528 9384 2592
rect 9448 2528 9464 2592
rect 9337 2512 9464 2528
rect 9337 2448 9384 2512
rect 9448 2448 9464 2512
rect 9337 2432 9464 2448
rect 9337 2368 9384 2432
rect 9448 2368 9464 2432
rect 9337 2352 9464 2368
rect 9337 2288 9384 2352
rect 9448 2288 9464 2352
rect 9337 2272 9464 2288
rect 9337 2208 9384 2272
rect 9448 2208 9464 2272
rect 9337 2192 9464 2208
rect 9337 2128 9384 2192
rect 9448 2128 9464 2192
rect 9337 2112 9464 2128
rect 9337 2048 9384 2112
rect 9448 2048 9464 2112
rect 9337 2032 9464 2048
rect 9337 1968 9384 2032
rect 9448 1968 9464 2032
rect 9337 1952 9464 1968
rect 9337 1888 9384 1952
rect 9448 1888 9464 1952
rect 9337 1872 9464 1888
rect 9337 1808 9384 1872
rect 9448 1808 9464 1872
rect 9337 1792 9464 1808
rect 9337 1728 9384 1792
rect 9448 1728 9464 1792
rect 9337 1712 9464 1728
rect 9337 1648 9384 1712
rect 9448 1648 9464 1712
rect 9337 1632 9464 1648
rect 9337 1568 9384 1632
rect 9448 1568 9464 1632
rect 9337 1552 9464 1568
rect 9337 1488 9384 1552
rect 9448 1488 9464 1552
rect 9337 1472 9464 1488
rect 9337 1408 9384 1472
rect 9448 1408 9464 1472
rect 9337 1392 9464 1408
rect 9337 1328 9384 1392
rect 9448 1328 9464 1392
rect 9337 1312 9464 1328
rect 9337 1248 9384 1312
rect 9448 1248 9464 1312
rect 9337 1232 9464 1248
rect 9337 1168 9384 1232
rect 9448 1168 9464 1232
rect 9337 1152 9464 1168
rect 9337 1088 9384 1152
rect 9448 1088 9464 1152
rect 9337 1072 9464 1088
rect 9337 1008 9384 1072
rect 9448 1008 9464 1072
rect 9337 992 9464 1008
rect 9337 928 9384 992
rect 9448 928 9464 992
rect 9337 912 9464 928
rect 9337 848 9384 912
rect 9448 848 9464 912
rect 9337 832 9464 848
rect 9337 768 9384 832
rect 9448 768 9464 832
rect 9337 752 9464 768
rect 9337 688 9384 752
rect 9448 688 9464 752
rect 9337 672 9464 688
rect 9337 608 9384 672
rect 9448 608 9464 672
rect 9337 592 9464 608
rect 9337 528 9384 592
rect 9448 528 9464 592
rect 9337 512 9464 528
rect 9337 448 9384 512
rect 9448 448 9464 512
rect 9337 432 9464 448
rect 9337 368 9384 432
rect 9448 368 9464 432
rect 9337 352 9464 368
rect 9337 288 9384 352
rect 9448 288 9464 352
rect 9337 272 9464 288
rect 9337 208 9384 272
rect 9448 208 9464 272
rect 9337 192 9464 208
rect 9337 128 9384 192
rect 9448 128 9464 192
rect 9337 112 9464 128
rect 9337 48 9384 112
rect 9448 48 9464 112
rect 9337 32 9464 48
rect 9337 -32 9384 32
rect 9448 -32 9464 32
rect 9337 -48 9464 -32
rect 9337 -112 9384 -48
rect 9448 -112 9464 -48
rect 9337 -128 9464 -112
rect 9337 -192 9384 -128
rect 9448 -192 9464 -128
rect 9337 -208 9464 -192
rect 9337 -272 9384 -208
rect 9448 -272 9464 -208
rect 9337 -288 9464 -272
rect 9337 -352 9384 -288
rect 9448 -352 9464 -288
rect 9337 -368 9464 -352
rect 9337 -432 9384 -368
rect 9448 -432 9464 -368
rect 9337 -448 9464 -432
rect 9337 -512 9384 -448
rect 9448 -512 9464 -448
rect 9337 -528 9464 -512
rect 9337 -592 9384 -528
rect 9448 -592 9464 -528
rect 9337 -608 9464 -592
rect 9337 -672 9384 -608
rect 9448 -672 9464 -608
rect 9337 -688 9464 -672
rect 9337 -752 9384 -688
rect 9448 -752 9464 -688
rect 9337 -768 9464 -752
rect 9337 -832 9384 -768
rect 9448 -832 9464 -768
rect 9337 -848 9464 -832
rect 9337 -912 9384 -848
rect 9448 -912 9464 -848
rect 9337 -928 9464 -912
rect 9337 -992 9384 -928
rect 9448 -992 9464 -928
rect 9337 -1008 9464 -992
rect 9337 -1072 9384 -1008
rect 9448 -1072 9464 -1008
rect 9337 -1088 9464 -1072
rect 9337 -1152 9384 -1088
rect 9448 -1152 9464 -1088
rect 9337 -1168 9464 -1152
rect 9337 -1232 9384 -1168
rect 9448 -1232 9464 -1168
rect 9337 -1248 9464 -1232
rect 9337 -1312 9384 -1248
rect 9448 -1312 9464 -1248
rect 9337 -1328 9464 -1312
rect 9337 -1392 9384 -1328
rect 9448 -1392 9464 -1328
rect 9337 -1408 9464 -1392
rect 9337 -1472 9384 -1408
rect 9448 -1472 9464 -1408
rect 9337 -1488 9464 -1472
rect 9337 -1552 9384 -1488
rect 9448 -1552 9464 -1488
rect 9337 -1568 9464 -1552
rect 9337 -1632 9384 -1568
rect 9448 -1632 9464 -1568
rect 9337 -1648 9464 -1632
rect 9337 -1712 9384 -1648
rect 9448 -1712 9464 -1648
rect 9337 -1728 9464 -1712
rect 9337 -1792 9384 -1728
rect 9448 -1792 9464 -1728
rect 9337 -1808 9464 -1792
rect 9337 -1872 9384 -1808
rect 9448 -1872 9464 -1808
rect 9337 -1888 9464 -1872
rect 9337 -1952 9384 -1888
rect 9448 -1952 9464 -1888
rect 9337 -1968 9464 -1952
rect 9337 -2032 9384 -1968
rect 9448 -2032 9464 -1968
rect 9337 -2048 9464 -2032
rect 9337 -2112 9384 -2048
rect 9448 -2112 9464 -2048
rect 9337 -2128 9464 -2112
rect 9337 -2192 9384 -2128
rect 9448 -2192 9464 -2128
rect 9337 -2208 9464 -2192
rect 9337 -2272 9384 -2208
rect 9448 -2272 9464 -2208
rect 9337 -2288 9464 -2272
rect 9337 -2352 9384 -2288
rect 9448 -2352 9464 -2288
rect 9337 -2368 9464 -2352
rect 9337 -2432 9384 -2368
rect 9448 -2432 9464 -2368
rect 9337 -2448 9464 -2432
rect 9337 -2512 9384 -2448
rect 9448 -2512 9464 -2448
rect 9337 -2528 9464 -2512
rect 9337 -2592 9384 -2528
rect 9448 -2592 9464 -2528
rect 9337 -2608 9464 -2592
rect 9337 -2672 9384 -2608
rect 9448 -2672 9464 -2608
rect 9337 -2688 9464 -2672
rect 9337 -2752 9384 -2688
rect 9448 -2752 9464 -2688
rect 9337 -2768 9464 -2752
rect 9337 -2832 9384 -2768
rect 9448 -2832 9464 -2768
rect 9337 -2848 9464 -2832
rect 9337 -2912 9384 -2848
rect 9448 -2912 9464 -2848
rect 9337 -2928 9464 -2912
rect 3018 -3008 3145 -2992
rect 3018 -3072 3065 -3008
rect 3129 -3072 3145 -3008
rect 3018 -3088 3145 -3072
rect 3018 -3212 3122 -3088
rect 3018 -3228 3145 -3212
rect 3018 -3292 3065 -3228
rect 3129 -3292 3145 -3228
rect 3018 -3308 3145 -3292
rect -3301 -3388 -3174 -3372
rect -3301 -3452 -3254 -3388
rect -3190 -3452 -3174 -3388
rect -3301 -3468 -3174 -3452
rect -3301 -3532 -3254 -3468
rect -3190 -3532 -3174 -3468
rect -3301 -3548 -3174 -3532
rect -3301 -3612 -3254 -3548
rect -3190 -3612 -3174 -3548
rect -3301 -3628 -3174 -3612
rect -3301 -3692 -3254 -3628
rect -3190 -3692 -3174 -3628
rect -3301 -3708 -3174 -3692
rect -3301 -3772 -3254 -3708
rect -3190 -3772 -3174 -3708
rect -3301 -3788 -3174 -3772
rect -3301 -3852 -3254 -3788
rect -3190 -3852 -3174 -3788
rect -3301 -3868 -3174 -3852
rect -3301 -3932 -3254 -3868
rect -3190 -3932 -3174 -3868
rect -3301 -3948 -3174 -3932
rect -3301 -4012 -3254 -3948
rect -3190 -4012 -3174 -3948
rect -3301 -4028 -3174 -4012
rect -3301 -4092 -3254 -4028
rect -3190 -4092 -3174 -4028
rect -3301 -4108 -3174 -4092
rect -3301 -4172 -3254 -4108
rect -3190 -4172 -3174 -4108
rect -3301 -4188 -3174 -4172
rect -3301 -4252 -3254 -4188
rect -3190 -4252 -3174 -4188
rect -3301 -4268 -3174 -4252
rect -3301 -4332 -3254 -4268
rect -3190 -4332 -3174 -4268
rect -3301 -4348 -3174 -4332
rect -3301 -4412 -3254 -4348
rect -3190 -4412 -3174 -4348
rect -3301 -4428 -3174 -4412
rect -3301 -4492 -3254 -4428
rect -3190 -4492 -3174 -4428
rect -3301 -4508 -3174 -4492
rect -3301 -4572 -3254 -4508
rect -3190 -4572 -3174 -4508
rect -3301 -4588 -3174 -4572
rect -3301 -4652 -3254 -4588
rect -3190 -4652 -3174 -4588
rect -3301 -4668 -3174 -4652
rect -3301 -4732 -3254 -4668
rect -3190 -4732 -3174 -4668
rect -3301 -4748 -3174 -4732
rect -3301 -4812 -3254 -4748
rect -3190 -4812 -3174 -4748
rect -3301 -4828 -3174 -4812
rect -3301 -4892 -3254 -4828
rect -3190 -4892 -3174 -4828
rect -3301 -4908 -3174 -4892
rect -3301 -4972 -3254 -4908
rect -3190 -4972 -3174 -4908
rect -3301 -4988 -3174 -4972
rect -3301 -5052 -3254 -4988
rect -3190 -5052 -3174 -4988
rect -3301 -5068 -3174 -5052
rect -3301 -5132 -3254 -5068
rect -3190 -5132 -3174 -5068
rect -3301 -5148 -3174 -5132
rect -3301 -5212 -3254 -5148
rect -3190 -5212 -3174 -5148
rect -3301 -5228 -3174 -5212
rect -3301 -5292 -3254 -5228
rect -3190 -5292 -3174 -5228
rect -3301 -5308 -3174 -5292
rect -3301 -5372 -3254 -5308
rect -3190 -5372 -3174 -5308
rect -3301 -5388 -3174 -5372
rect -3301 -5452 -3254 -5388
rect -3190 -5452 -3174 -5388
rect -3301 -5468 -3174 -5452
rect -3301 -5532 -3254 -5468
rect -3190 -5532 -3174 -5468
rect -3301 -5548 -3174 -5532
rect -3301 -5612 -3254 -5548
rect -3190 -5612 -3174 -5548
rect -3301 -5628 -3174 -5612
rect -3301 -5692 -3254 -5628
rect -3190 -5692 -3174 -5628
rect -3301 -5708 -3174 -5692
rect -3301 -5772 -3254 -5708
rect -3190 -5772 -3174 -5708
rect -3301 -5788 -3174 -5772
rect -3301 -5852 -3254 -5788
rect -3190 -5852 -3174 -5788
rect -3301 -5868 -3174 -5852
rect -3301 -5932 -3254 -5868
rect -3190 -5932 -3174 -5868
rect -3301 -5948 -3174 -5932
rect -3301 -6012 -3254 -5948
rect -3190 -6012 -3174 -5948
rect -3301 -6028 -3174 -6012
rect -3301 -6092 -3254 -6028
rect -3190 -6092 -3174 -6028
rect -3301 -6108 -3174 -6092
rect -3301 -6172 -3254 -6108
rect -3190 -6172 -3174 -6108
rect -3301 -6188 -3174 -6172
rect -3301 -6252 -3254 -6188
rect -3190 -6252 -3174 -6188
rect -3301 -6268 -3174 -6252
rect -3301 -6332 -3254 -6268
rect -3190 -6332 -3174 -6268
rect -3301 -6348 -3174 -6332
rect -3301 -6412 -3254 -6348
rect -3190 -6412 -3174 -6348
rect -3301 -6428 -3174 -6412
rect -3301 -6492 -3254 -6428
rect -3190 -6492 -3174 -6428
rect -3301 -6508 -3174 -6492
rect -3301 -6572 -3254 -6508
rect -3190 -6572 -3174 -6508
rect -3301 -6588 -3174 -6572
rect -3301 -6652 -3254 -6588
rect -3190 -6652 -3174 -6588
rect -3301 -6668 -3174 -6652
rect -3301 -6732 -3254 -6668
rect -3190 -6732 -3174 -6668
rect -3301 -6748 -3174 -6732
rect -3301 -6812 -3254 -6748
rect -3190 -6812 -3174 -6748
rect -3301 -6828 -3174 -6812
rect -3301 -6892 -3254 -6828
rect -3190 -6892 -3174 -6828
rect -3301 -6908 -3174 -6892
rect -3301 -6972 -3254 -6908
rect -3190 -6972 -3174 -6908
rect -3301 -6988 -3174 -6972
rect -3301 -7052 -3254 -6988
rect -3190 -7052 -3174 -6988
rect -3301 -7068 -3174 -7052
rect -3301 -7132 -3254 -7068
rect -3190 -7132 -3174 -7068
rect -3301 -7148 -3174 -7132
rect -3301 -7212 -3254 -7148
rect -3190 -7212 -3174 -7148
rect -3301 -7228 -3174 -7212
rect -3301 -7292 -3254 -7228
rect -3190 -7292 -3174 -7228
rect -3301 -7308 -3174 -7292
rect -3301 -7372 -3254 -7308
rect -3190 -7372 -3174 -7308
rect -3301 -7388 -3174 -7372
rect -3301 -7452 -3254 -7388
rect -3190 -7452 -3174 -7388
rect -3301 -7468 -3174 -7452
rect -3301 -7532 -3254 -7468
rect -3190 -7532 -3174 -7468
rect -3301 -7548 -3174 -7532
rect -3301 -7612 -3254 -7548
rect -3190 -7612 -3174 -7548
rect -3301 -7628 -3174 -7612
rect -3301 -7692 -3254 -7628
rect -3190 -7692 -3174 -7628
rect -3301 -7708 -3174 -7692
rect -3301 -7772 -3254 -7708
rect -3190 -7772 -3174 -7708
rect -3301 -7788 -3174 -7772
rect -3301 -7852 -3254 -7788
rect -3190 -7852 -3174 -7788
rect -3301 -7868 -3174 -7852
rect -3301 -7932 -3254 -7868
rect -3190 -7932 -3174 -7868
rect -3301 -7948 -3174 -7932
rect -3301 -8012 -3254 -7948
rect -3190 -8012 -3174 -7948
rect -3301 -8028 -3174 -8012
rect -3301 -8092 -3254 -8028
rect -3190 -8092 -3174 -8028
rect -3301 -8108 -3174 -8092
rect -3301 -8172 -3254 -8108
rect -3190 -8172 -3174 -8108
rect -3301 -8188 -3174 -8172
rect -3301 -8252 -3254 -8188
rect -3190 -8252 -3174 -8188
rect -3301 -8268 -3174 -8252
rect -3301 -8332 -3254 -8268
rect -3190 -8332 -3174 -8268
rect -3301 -8348 -3174 -8332
rect -3301 -8412 -3254 -8348
rect -3190 -8412 -3174 -8348
rect -3301 -8428 -3174 -8412
rect -3301 -8492 -3254 -8428
rect -3190 -8492 -3174 -8428
rect -3301 -8508 -3174 -8492
rect -3301 -8572 -3254 -8508
rect -3190 -8572 -3174 -8508
rect -3301 -8588 -3174 -8572
rect -3301 -8652 -3254 -8588
rect -3190 -8652 -3174 -8588
rect -3301 -8668 -3174 -8652
rect -3301 -8732 -3254 -8668
rect -3190 -8732 -3174 -8668
rect -3301 -8748 -3174 -8732
rect -3301 -8812 -3254 -8748
rect -3190 -8812 -3174 -8748
rect -3301 -8828 -3174 -8812
rect -3301 -8892 -3254 -8828
rect -3190 -8892 -3174 -8828
rect -3301 -8908 -3174 -8892
rect -3301 -8972 -3254 -8908
rect -3190 -8972 -3174 -8908
rect -3301 -8988 -3174 -8972
rect -3301 -9052 -3254 -8988
rect -3190 -9052 -3174 -8988
rect -3301 -9068 -3174 -9052
rect -3301 -9132 -3254 -9068
rect -3190 -9132 -3174 -9068
rect -3301 -9148 -3174 -9132
rect -3301 -9212 -3254 -9148
rect -3190 -9212 -3174 -9148
rect -3301 -9228 -3174 -9212
rect -9620 -9308 -9493 -9292
rect -9620 -9372 -9573 -9308
rect -9509 -9372 -9493 -9308
rect -9620 -9388 -9493 -9372
rect -9620 -9512 -9516 -9388
rect -9620 -9528 -9493 -9512
rect -9620 -9592 -9573 -9528
rect -9509 -9592 -9493 -9528
rect -9620 -9608 -9493 -9592
rect -15939 -9688 -15812 -9672
rect -15939 -9752 -15892 -9688
rect -15828 -9752 -15812 -9688
rect -15939 -9768 -15812 -9752
rect -15939 -9832 -15892 -9768
rect -15828 -9832 -15812 -9768
rect -15939 -9848 -15812 -9832
rect -15939 -9912 -15892 -9848
rect -15828 -9912 -15812 -9848
rect -15939 -9928 -15812 -9912
rect -15939 -9992 -15892 -9928
rect -15828 -9992 -15812 -9928
rect -15939 -10008 -15812 -9992
rect -15939 -10072 -15892 -10008
rect -15828 -10072 -15812 -10008
rect -15939 -10088 -15812 -10072
rect -15939 -10152 -15892 -10088
rect -15828 -10152 -15812 -10088
rect -15939 -10168 -15812 -10152
rect -15939 -10232 -15892 -10168
rect -15828 -10232 -15812 -10168
rect -15939 -10248 -15812 -10232
rect -15939 -10312 -15892 -10248
rect -15828 -10312 -15812 -10248
rect -15939 -10328 -15812 -10312
rect -15939 -10392 -15892 -10328
rect -15828 -10392 -15812 -10328
rect -15939 -10408 -15812 -10392
rect -15939 -10472 -15892 -10408
rect -15828 -10472 -15812 -10408
rect -15939 -10488 -15812 -10472
rect -15939 -10552 -15892 -10488
rect -15828 -10552 -15812 -10488
rect -15939 -10568 -15812 -10552
rect -15939 -10632 -15892 -10568
rect -15828 -10632 -15812 -10568
rect -15939 -10648 -15812 -10632
rect -15939 -10712 -15892 -10648
rect -15828 -10712 -15812 -10648
rect -15939 -10728 -15812 -10712
rect -15939 -10792 -15892 -10728
rect -15828 -10792 -15812 -10728
rect -15939 -10808 -15812 -10792
rect -15939 -10872 -15892 -10808
rect -15828 -10872 -15812 -10808
rect -15939 -10888 -15812 -10872
rect -15939 -10952 -15892 -10888
rect -15828 -10952 -15812 -10888
rect -15939 -10968 -15812 -10952
rect -15939 -11032 -15892 -10968
rect -15828 -11032 -15812 -10968
rect -15939 -11048 -15812 -11032
rect -15939 -11112 -15892 -11048
rect -15828 -11112 -15812 -11048
rect -15939 -11128 -15812 -11112
rect -15939 -11192 -15892 -11128
rect -15828 -11192 -15812 -11128
rect -15939 -11208 -15812 -11192
rect -15939 -11272 -15892 -11208
rect -15828 -11272 -15812 -11208
rect -15939 -11288 -15812 -11272
rect -15939 -11352 -15892 -11288
rect -15828 -11352 -15812 -11288
rect -15939 -11368 -15812 -11352
rect -15939 -11432 -15892 -11368
rect -15828 -11432 -15812 -11368
rect -15939 -11448 -15812 -11432
rect -15939 -11512 -15892 -11448
rect -15828 -11512 -15812 -11448
rect -15939 -11528 -15812 -11512
rect -15939 -11592 -15892 -11528
rect -15828 -11592 -15812 -11528
rect -15939 -11608 -15812 -11592
rect -15939 -11672 -15892 -11608
rect -15828 -11672 -15812 -11608
rect -15939 -11688 -15812 -11672
rect -15939 -11752 -15892 -11688
rect -15828 -11752 -15812 -11688
rect -15939 -11768 -15812 -11752
rect -15939 -11832 -15892 -11768
rect -15828 -11832 -15812 -11768
rect -15939 -11848 -15812 -11832
rect -15939 -11912 -15892 -11848
rect -15828 -11912 -15812 -11848
rect -15939 -11928 -15812 -11912
rect -15939 -11992 -15892 -11928
rect -15828 -11992 -15812 -11928
rect -15939 -12008 -15812 -11992
rect -15939 -12072 -15892 -12008
rect -15828 -12072 -15812 -12008
rect -15939 -12088 -15812 -12072
rect -15939 -12152 -15892 -12088
rect -15828 -12152 -15812 -12088
rect -15939 -12168 -15812 -12152
rect -15939 -12232 -15892 -12168
rect -15828 -12232 -15812 -12168
rect -15939 -12248 -15812 -12232
rect -15939 -12312 -15892 -12248
rect -15828 -12312 -15812 -12248
rect -15939 -12328 -15812 -12312
rect -15939 -12392 -15892 -12328
rect -15828 -12392 -15812 -12328
rect -15939 -12408 -15812 -12392
rect -15939 -12472 -15892 -12408
rect -15828 -12472 -15812 -12408
rect -15939 -12488 -15812 -12472
rect -15939 -12552 -15892 -12488
rect -15828 -12552 -15812 -12488
rect -15939 -12568 -15812 -12552
rect -15939 -12632 -15892 -12568
rect -15828 -12632 -15812 -12568
rect -15939 -12648 -15812 -12632
rect -15939 -12712 -15892 -12648
rect -15828 -12712 -15812 -12648
rect -15939 -12728 -15812 -12712
rect -15939 -12792 -15892 -12728
rect -15828 -12792 -15812 -12728
rect -15939 -12808 -15812 -12792
rect -15939 -12872 -15892 -12808
rect -15828 -12872 -15812 -12808
rect -15939 -12888 -15812 -12872
rect -15939 -12952 -15892 -12888
rect -15828 -12952 -15812 -12888
rect -15939 -12968 -15812 -12952
rect -15939 -13032 -15892 -12968
rect -15828 -13032 -15812 -12968
rect -15939 -13048 -15812 -13032
rect -15939 -13112 -15892 -13048
rect -15828 -13112 -15812 -13048
rect -15939 -13128 -15812 -13112
rect -15939 -13192 -15892 -13128
rect -15828 -13192 -15812 -13128
rect -15939 -13208 -15812 -13192
rect -15939 -13272 -15892 -13208
rect -15828 -13272 -15812 -13208
rect -15939 -13288 -15812 -13272
rect -15939 -13352 -15892 -13288
rect -15828 -13352 -15812 -13288
rect -15939 -13368 -15812 -13352
rect -15939 -13432 -15892 -13368
rect -15828 -13432 -15812 -13368
rect -15939 -13448 -15812 -13432
rect -15939 -13512 -15892 -13448
rect -15828 -13512 -15812 -13448
rect -15939 -13528 -15812 -13512
rect -15939 -13592 -15892 -13528
rect -15828 -13592 -15812 -13528
rect -15939 -13608 -15812 -13592
rect -15939 -13672 -15892 -13608
rect -15828 -13672 -15812 -13608
rect -15939 -13688 -15812 -13672
rect -15939 -13752 -15892 -13688
rect -15828 -13752 -15812 -13688
rect -15939 -13768 -15812 -13752
rect -15939 -13832 -15892 -13768
rect -15828 -13832 -15812 -13768
rect -15939 -13848 -15812 -13832
rect -15939 -13912 -15892 -13848
rect -15828 -13912 -15812 -13848
rect -15939 -13928 -15812 -13912
rect -15939 -13992 -15892 -13928
rect -15828 -13992 -15812 -13928
rect -15939 -14008 -15812 -13992
rect -15939 -14072 -15892 -14008
rect -15828 -14072 -15812 -14008
rect -15939 -14088 -15812 -14072
rect -15939 -14152 -15892 -14088
rect -15828 -14152 -15812 -14088
rect -15939 -14168 -15812 -14152
rect -15939 -14232 -15892 -14168
rect -15828 -14232 -15812 -14168
rect -15939 -14248 -15812 -14232
rect -15939 -14312 -15892 -14248
rect -15828 -14312 -15812 -14248
rect -15939 -14328 -15812 -14312
rect -15939 -14392 -15892 -14328
rect -15828 -14392 -15812 -14328
rect -15939 -14408 -15812 -14392
rect -15939 -14472 -15892 -14408
rect -15828 -14472 -15812 -14408
rect -15939 -14488 -15812 -14472
rect -15939 -14552 -15892 -14488
rect -15828 -14552 -15812 -14488
rect -15939 -14568 -15812 -14552
rect -15939 -14632 -15892 -14568
rect -15828 -14632 -15812 -14568
rect -15939 -14648 -15812 -14632
rect -15939 -14712 -15892 -14648
rect -15828 -14712 -15812 -14648
rect -15939 -14728 -15812 -14712
rect -15939 -14792 -15892 -14728
rect -15828 -14792 -15812 -14728
rect -15939 -14808 -15812 -14792
rect -15939 -14872 -15892 -14808
rect -15828 -14872 -15812 -14808
rect -15939 -14888 -15812 -14872
rect -15939 -14952 -15892 -14888
rect -15828 -14952 -15812 -14888
rect -15939 -14968 -15812 -14952
rect -15939 -15032 -15892 -14968
rect -15828 -15032 -15812 -14968
rect -15939 -15048 -15812 -15032
rect -15939 -15112 -15892 -15048
rect -15828 -15112 -15812 -15048
rect -15939 -15128 -15812 -15112
rect -15939 -15192 -15892 -15128
rect -15828 -15192 -15812 -15128
rect -15939 -15208 -15812 -15192
rect -15939 -15272 -15892 -15208
rect -15828 -15272 -15812 -15208
rect -15939 -15288 -15812 -15272
rect -15939 -15352 -15892 -15288
rect -15828 -15352 -15812 -15288
rect -15939 -15368 -15812 -15352
rect -15939 -15432 -15892 -15368
rect -15828 -15432 -15812 -15368
rect -15939 -15448 -15812 -15432
rect -15939 -15512 -15892 -15448
rect -15828 -15512 -15812 -15448
rect -15939 -15528 -15812 -15512
rect -22258 -15608 -22131 -15592
rect -22258 -15672 -22211 -15608
rect -22147 -15672 -22131 -15608
rect -22258 -15688 -22131 -15672
rect -22258 -15812 -22154 -15688
rect -22258 -15828 -22131 -15812
rect -22258 -15892 -22211 -15828
rect -22147 -15892 -22131 -15828
rect -22258 -15908 -22131 -15892
rect -28577 -15988 -28450 -15972
rect -28577 -16052 -28530 -15988
rect -28466 -16052 -28450 -15988
rect -28577 -16068 -28450 -16052
rect -28577 -16132 -28530 -16068
rect -28466 -16132 -28450 -16068
rect -28577 -16148 -28450 -16132
rect -28577 -16212 -28530 -16148
rect -28466 -16212 -28450 -16148
rect -28577 -16228 -28450 -16212
rect -28577 -16292 -28530 -16228
rect -28466 -16292 -28450 -16228
rect -28577 -16308 -28450 -16292
rect -28577 -16372 -28530 -16308
rect -28466 -16372 -28450 -16308
rect -28577 -16388 -28450 -16372
rect -28577 -16452 -28530 -16388
rect -28466 -16452 -28450 -16388
rect -28577 -16468 -28450 -16452
rect -28577 -16532 -28530 -16468
rect -28466 -16532 -28450 -16468
rect -28577 -16548 -28450 -16532
rect -28577 -16612 -28530 -16548
rect -28466 -16612 -28450 -16548
rect -28577 -16628 -28450 -16612
rect -28577 -16692 -28530 -16628
rect -28466 -16692 -28450 -16628
rect -28577 -16708 -28450 -16692
rect -28577 -16772 -28530 -16708
rect -28466 -16772 -28450 -16708
rect -28577 -16788 -28450 -16772
rect -28577 -16852 -28530 -16788
rect -28466 -16852 -28450 -16788
rect -28577 -16868 -28450 -16852
rect -28577 -16932 -28530 -16868
rect -28466 -16932 -28450 -16868
rect -28577 -16948 -28450 -16932
rect -28577 -17012 -28530 -16948
rect -28466 -17012 -28450 -16948
rect -28577 -17028 -28450 -17012
rect -28577 -17092 -28530 -17028
rect -28466 -17092 -28450 -17028
rect -28577 -17108 -28450 -17092
rect -28577 -17172 -28530 -17108
rect -28466 -17172 -28450 -17108
rect -28577 -17188 -28450 -17172
rect -28577 -17252 -28530 -17188
rect -28466 -17252 -28450 -17188
rect -28577 -17268 -28450 -17252
rect -28577 -17332 -28530 -17268
rect -28466 -17332 -28450 -17268
rect -28577 -17348 -28450 -17332
rect -28577 -17412 -28530 -17348
rect -28466 -17412 -28450 -17348
rect -28577 -17428 -28450 -17412
rect -28577 -17492 -28530 -17428
rect -28466 -17492 -28450 -17428
rect -28577 -17508 -28450 -17492
rect -28577 -17572 -28530 -17508
rect -28466 -17572 -28450 -17508
rect -28577 -17588 -28450 -17572
rect -28577 -17652 -28530 -17588
rect -28466 -17652 -28450 -17588
rect -28577 -17668 -28450 -17652
rect -28577 -17732 -28530 -17668
rect -28466 -17732 -28450 -17668
rect -28577 -17748 -28450 -17732
rect -28577 -17812 -28530 -17748
rect -28466 -17812 -28450 -17748
rect -28577 -17828 -28450 -17812
rect -28577 -17892 -28530 -17828
rect -28466 -17892 -28450 -17828
rect -28577 -17908 -28450 -17892
rect -28577 -17972 -28530 -17908
rect -28466 -17972 -28450 -17908
rect -28577 -17988 -28450 -17972
rect -28577 -18052 -28530 -17988
rect -28466 -18052 -28450 -17988
rect -28577 -18068 -28450 -18052
rect -28577 -18132 -28530 -18068
rect -28466 -18132 -28450 -18068
rect -28577 -18148 -28450 -18132
rect -28577 -18212 -28530 -18148
rect -28466 -18212 -28450 -18148
rect -28577 -18228 -28450 -18212
rect -28577 -18292 -28530 -18228
rect -28466 -18292 -28450 -18228
rect -28577 -18308 -28450 -18292
rect -28577 -18372 -28530 -18308
rect -28466 -18372 -28450 -18308
rect -28577 -18388 -28450 -18372
rect -28577 -18452 -28530 -18388
rect -28466 -18452 -28450 -18388
rect -28577 -18468 -28450 -18452
rect -28577 -18532 -28530 -18468
rect -28466 -18532 -28450 -18468
rect -28577 -18548 -28450 -18532
rect -28577 -18612 -28530 -18548
rect -28466 -18612 -28450 -18548
rect -28577 -18628 -28450 -18612
rect -28577 -18692 -28530 -18628
rect -28466 -18692 -28450 -18628
rect -28577 -18708 -28450 -18692
rect -28577 -18772 -28530 -18708
rect -28466 -18772 -28450 -18708
rect -28577 -18788 -28450 -18772
rect -28577 -18852 -28530 -18788
rect -28466 -18852 -28450 -18788
rect -28577 -18868 -28450 -18852
rect -28577 -18932 -28530 -18868
rect -28466 -18932 -28450 -18868
rect -28577 -18948 -28450 -18932
rect -28577 -19012 -28530 -18948
rect -28466 -19012 -28450 -18948
rect -28577 -19028 -28450 -19012
rect -28577 -19092 -28530 -19028
rect -28466 -19092 -28450 -19028
rect -28577 -19108 -28450 -19092
rect -28577 -19172 -28530 -19108
rect -28466 -19172 -28450 -19108
rect -28577 -19188 -28450 -19172
rect -28577 -19252 -28530 -19188
rect -28466 -19252 -28450 -19188
rect -28577 -19268 -28450 -19252
rect -28577 -19332 -28530 -19268
rect -28466 -19332 -28450 -19268
rect -28577 -19348 -28450 -19332
rect -28577 -19412 -28530 -19348
rect -28466 -19412 -28450 -19348
rect -28577 -19428 -28450 -19412
rect -28577 -19492 -28530 -19428
rect -28466 -19492 -28450 -19428
rect -28577 -19508 -28450 -19492
rect -28577 -19572 -28530 -19508
rect -28466 -19572 -28450 -19508
rect -28577 -19588 -28450 -19572
rect -28577 -19652 -28530 -19588
rect -28466 -19652 -28450 -19588
rect -28577 -19668 -28450 -19652
rect -28577 -19732 -28530 -19668
rect -28466 -19732 -28450 -19668
rect -28577 -19748 -28450 -19732
rect -28577 -19812 -28530 -19748
rect -28466 -19812 -28450 -19748
rect -28577 -19828 -28450 -19812
rect -28577 -19892 -28530 -19828
rect -28466 -19892 -28450 -19828
rect -28577 -19908 -28450 -19892
rect -28577 -19972 -28530 -19908
rect -28466 -19972 -28450 -19908
rect -28577 -19988 -28450 -19972
rect -28577 -20052 -28530 -19988
rect -28466 -20052 -28450 -19988
rect -28577 -20068 -28450 -20052
rect -28577 -20132 -28530 -20068
rect -28466 -20132 -28450 -20068
rect -28577 -20148 -28450 -20132
rect -28577 -20212 -28530 -20148
rect -28466 -20212 -28450 -20148
rect -28577 -20228 -28450 -20212
rect -28577 -20292 -28530 -20228
rect -28466 -20292 -28450 -20228
rect -28577 -20308 -28450 -20292
rect -28577 -20372 -28530 -20308
rect -28466 -20372 -28450 -20308
rect -28577 -20388 -28450 -20372
rect -28577 -20452 -28530 -20388
rect -28466 -20452 -28450 -20388
rect -28577 -20468 -28450 -20452
rect -28577 -20532 -28530 -20468
rect -28466 -20532 -28450 -20468
rect -28577 -20548 -28450 -20532
rect -28577 -20612 -28530 -20548
rect -28466 -20612 -28450 -20548
rect -28577 -20628 -28450 -20612
rect -28577 -20692 -28530 -20628
rect -28466 -20692 -28450 -20628
rect -28577 -20708 -28450 -20692
rect -28577 -20772 -28530 -20708
rect -28466 -20772 -28450 -20708
rect -28577 -20788 -28450 -20772
rect -28577 -20852 -28530 -20788
rect -28466 -20852 -28450 -20788
rect -28577 -20868 -28450 -20852
rect -28577 -20932 -28530 -20868
rect -28466 -20932 -28450 -20868
rect -28577 -20948 -28450 -20932
rect -28577 -21012 -28530 -20948
rect -28466 -21012 -28450 -20948
rect -28577 -21028 -28450 -21012
rect -28577 -21092 -28530 -21028
rect -28466 -21092 -28450 -21028
rect -28577 -21108 -28450 -21092
rect -28577 -21172 -28530 -21108
rect -28466 -21172 -28450 -21108
rect -28577 -21188 -28450 -21172
rect -28577 -21252 -28530 -21188
rect -28466 -21252 -28450 -21188
rect -28577 -21268 -28450 -21252
rect -28577 -21332 -28530 -21268
rect -28466 -21332 -28450 -21268
rect -28577 -21348 -28450 -21332
rect -28577 -21412 -28530 -21348
rect -28466 -21412 -28450 -21348
rect -28577 -21428 -28450 -21412
rect -28577 -21492 -28530 -21428
rect -28466 -21492 -28450 -21428
rect -28577 -21508 -28450 -21492
rect -28577 -21572 -28530 -21508
rect -28466 -21572 -28450 -21508
rect -28577 -21588 -28450 -21572
rect -28577 -21652 -28530 -21588
rect -28466 -21652 -28450 -21588
rect -28577 -21668 -28450 -21652
rect -28577 -21732 -28530 -21668
rect -28466 -21732 -28450 -21668
rect -28577 -21748 -28450 -21732
rect -28577 -21812 -28530 -21748
rect -28466 -21812 -28450 -21748
rect -28577 -21828 -28450 -21812
rect -34896 -21908 -34769 -21892
rect -34896 -21972 -34849 -21908
rect -34785 -21972 -34769 -21908
rect -34896 -21988 -34769 -21972
rect -34896 -22112 -34792 -21988
rect -34896 -22128 -34769 -22112
rect -34896 -22192 -34849 -22128
rect -34785 -22192 -34769 -22128
rect -34896 -22208 -34769 -22192
rect -41215 -22288 -41088 -22272
rect -41215 -22352 -41168 -22288
rect -41104 -22352 -41088 -22288
rect -41215 -22368 -41088 -22352
rect -41215 -22432 -41168 -22368
rect -41104 -22432 -41088 -22368
rect -41215 -22448 -41088 -22432
rect -41215 -22512 -41168 -22448
rect -41104 -22512 -41088 -22448
rect -41215 -22528 -41088 -22512
rect -41215 -22592 -41168 -22528
rect -41104 -22592 -41088 -22528
rect -41215 -22608 -41088 -22592
rect -41215 -22672 -41168 -22608
rect -41104 -22672 -41088 -22608
rect -41215 -22688 -41088 -22672
rect -41215 -22752 -41168 -22688
rect -41104 -22752 -41088 -22688
rect -41215 -22768 -41088 -22752
rect -41215 -22832 -41168 -22768
rect -41104 -22832 -41088 -22768
rect -41215 -22848 -41088 -22832
rect -41215 -22912 -41168 -22848
rect -41104 -22912 -41088 -22848
rect -41215 -22928 -41088 -22912
rect -41215 -22992 -41168 -22928
rect -41104 -22992 -41088 -22928
rect -41215 -23008 -41088 -22992
rect -41215 -23072 -41168 -23008
rect -41104 -23072 -41088 -23008
rect -41215 -23088 -41088 -23072
rect -41215 -23152 -41168 -23088
rect -41104 -23152 -41088 -23088
rect -41215 -23168 -41088 -23152
rect -41215 -23232 -41168 -23168
rect -41104 -23232 -41088 -23168
rect -41215 -23248 -41088 -23232
rect -41215 -23312 -41168 -23248
rect -41104 -23312 -41088 -23248
rect -41215 -23328 -41088 -23312
rect -41215 -23392 -41168 -23328
rect -41104 -23392 -41088 -23328
rect -41215 -23408 -41088 -23392
rect -41215 -23472 -41168 -23408
rect -41104 -23472 -41088 -23408
rect -41215 -23488 -41088 -23472
rect -41215 -23552 -41168 -23488
rect -41104 -23552 -41088 -23488
rect -41215 -23568 -41088 -23552
rect -41215 -23632 -41168 -23568
rect -41104 -23632 -41088 -23568
rect -41215 -23648 -41088 -23632
rect -41215 -23712 -41168 -23648
rect -41104 -23712 -41088 -23648
rect -41215 -23728 -41088 -23712
rect -41215 -23792 -41168 -23728
rect -41104 -23792 -41088 -23728
rect -41215 -23808 -41088 -23792
rect -41215 -23872 -41168 -23808
rect -41104 -23872 -41088 -23808
rect -41215 -23888 -41088 -23872
rect -41215 -23952 -41168 -23888
rect -41104 -23952 -41088 -23888
rect -41215 -23968 -41088 -23952
rect -41215 -24032 -41168 -23968
rect -41104 -24032 -41088 -23968
rect -41215 -24048 -41088 -24032
rect -41215 -24112 -41168 -24048
rect -41104 -24112 -41088 -24048
rect -41215 -24128 -41088 -24112
rect -41215 -24192 -41168 -24128
rect -41104 -24192 -41088 -24128
rect -41215 -24208 -41088 -24192
rect -41215 -24272 -41168 -24208
rect -41104 -24272 -41088 -24208
rect -41215 -24288 -41088 -24272
rect -41215 -24352 -41168 -24288
rect -41104 -24352 -41088 -24288
rect -41215 -24368 -41088 -24352
rect -41215 -24432 -41168 -24368
rect -41104 -24432 -41088 -24368
rect -41215 -24448 -41088 -24432
rect -41215 -24512 -41168 -24448
rect -41104 -24512 -41088 -24448
rect -41215 -24528 -41088 -24512
rect -41215 -24592 -41168 -24528
rect -41104 -24592 -41088 -24528
rect -41215 -24608 -41088 -24592
rect -41215 -24672 -41168 -24608
rect -41104 -24672 -41088 -24608
rect -41215 -24688 -41088 -24672
rect -41215 -24752 -41168 -24688
rect -41104 -24752 -41088 -24688
rect -41215 -24768 -41088 -24752
rect -41215 -24832 -41168 -24768
rect -41104 -24832 -41088 -24768
rect -41215 -24848 -41088 -24832
rect -41215 -24912 -41168 -24848
rect -41104 -24912 -41088 -24848
rect -41215 -24928 -41088 -24912
rect -41215 -24992 -41168 -24928
rect -41104 -24992 -41088 -24928
rect -41215 -25008 -41088 -24992
rect -41215 -25072 -41168 -25008
rect -41104 -25072 -41088 -25008
rect -41215 -25088 -41088 -25072
rect -41215 -25152 -41168 -25088
rect -41104 -25152 -41088 -25088
rect -41215 -25168 -41088 -25152
rect -41215 -25232 -41168 -25168
rect -41104 -25232 -41088 -25168
rect -41215 -25248 -41088 -25232
rect -41215 -25312 -41168 -25248
rect -41104 -25312 -41088 -25248
rect -41215 -25328 -41088 -25312
rect -41215 -25392 -41168 -25328
rect -41104 -25392 -41088 -25328
rect -41215 -25408 -41088 -25392
rect -41215 -25472 -41168 -25408
rect -41104 -25472 -41088 -25408
rect -41215 -25488 -41088 -25472
rect -41215 -25552 -41168 -25488
rect -41104 -25552 -41088 -25488
rect -41215 -25568 -41088 -25552
rect -41215 -25632 -41168 -25568
rect -41104 -25632 -41088 -25568
rect -41215 -25648 -41088 -25632
rect -41215 -25712 -41168 -25648
rect -41104 -25712 -41088 -25648
rect -41215 -25728 -41088 -25712
rect -41215 -25792 -41168 -25728
rect -41104 -25792 -41088 -25728
rect -41215 -25808 -41088 -25792
rect -41215 -25872 -41168 -25808
rect -41104 -25872 -41088 -25808
rect -41215 -25888 -41088 -25872
rect -41215 -25952 -41168 -25888
rect -41104 -25952 -41088 -25888
rect -41215 -25968 -41088 -25952
rect -41215 -26032 -41168 -25968
rect -41104 -26032 -41088 -25968
rect -41215 -26048 -41088 -26032
rect -41215 -26112 -41168 -26048
rect -41104 -26112 -41088 -26048
rect -41215 -26128 -41088 -26112
rect -41215 -26192 -41168 -26128
rect -41104 -26192 -41088 -26128
rect -41215 -26208 -41088 -26192
rect -41215 -26272 -41168 -26208
rect -41104 -26272 -41088 -26208
rect -41215 -26288 -41088 -26272
rect -41215 -26352 -41168 -26288
rect -41104 -26352 -41088 -26288
rect -41215 -26368 -41088 -26352
rect -41215 -26432 -41168 -26368
rect -41104 -26432 -41088 -26368
rect -41215 -26448 -41088 -26432
rect -41215 -26512 -41168 -26448
rect -41104 -26512 -41088 -26448
rect -41215 -26528 -41088 -26512
rect -41215 -26592 -41168 -26528
rect -41104 -26592 -41088 -26528
rect -41215 -26608 -41088 -26592
rect -41215 -26672 -41168 -26608
rect -41104 -26672 -41088 -26608
rect -41215 -26688 -41088 -26672
rect -41215 -26752 -41168 -26688
rect -41104 -26752 -41088 -26688
rect -41215 -26768 -41088 -26752
rect -41215 -26832 -41168 -26768
rect -41104 -26832 -41088 -26768
rect -41215 -26848 -41088 -26832
rect -41215 -26912 -41168 -26848
rect -41104 -26912 -41088 -26848
rect -41215 -26928 -41088 -26912
rect -41215 -26992 -41168 -26928
rect -41104 -26992 -41088 -26928
rect -41215 -27008 -41088 -26992
rect -41215 -27072 -41168 -27008
rect -41104 -27072 -41088 -27008
rect -41215 -27088 -41088 -27072
rect -41215 -27152 -41168 -27088
rect -41104 -27152 -41088 -27088
rect -41215 -27168 -41088 -27152
rect -41215 -27232 -41168 -27168
rect -41104 -27232 -41088 -27168
rect -41215 -27248 -41088 -27232
rect -41215 -27312 -41168 -27248
rect -41104 -27312 -41088 -27248
rect -41215 -27328 -41088 -27312
rect -41215 -27392 -41168 -27328
rect -41104 -27392 -41088 -27328
rect -41215 -27408 -41088 -27392
rect -41215 -27472 -41168 -27408
rect -41104 -27472 -41088 -27408
rect -41215 -27488 -41088 -27472
rect -41215 -27552 -41168 -27488
rect -41104 -27552 -41088 -27488
rect -41215 -27568 -41088 -27552
rect -41215 -27632 -41168 -27568
rect -41104 -27632 -41088 -27568
rect -41215 -27648 -41088 -27632
rect -41215 -27712 -41168 -27648
rect -41104 -27712 -41088 -27648
rect -41215 -27728 -41088 -27712
rect -41215 -27792 -41168 -27728
rect -41104 -27792 -41088 -27728
rect -41215 -27808 -41088 -27792
rect -41215 -27872 -41168 -27808
rect -41104 -27872 -41088 -27808
rect -41215 -27888 -41088 -27872
rect -41215 -27952 -41168 -27888
rect -41104 -27952 -41088 -27888
rect -41215 -27968 -41088 -27952
rect -41215 -28032 -41168 -27968
rect -41104 -28032 -41088 -27968
rect -41215 -28048 -41088 -28032
rect -41215 -28112 -41168 -28048
rect -41104 -28112 -41088 -28048
rect -41215 -28128 -41088 -28112
rect -44335 -28539 -44231 -28161
rect -41215 -28192 -41168 -28128
rect -41104 -28192 -41088 -28128
rect -40925 -22248 -35003 -22239
rect -40925 -28152 -40916 -22248
rect -35012 -28152 -35003 -22248
rect -40925 -28161 -35003 -28152
rect -34896 -22272 -34849 -22208
rect -34785 -22272 -34769 -22208
rect -31697 -22239 -31593 -21861
rect -28577 -21892 -28530 -21828
rect -28466 -21892 -28450 -21828
rect -28287 -15948 -22365 -15939
rect -28287 -21852 -28278 -15948
rect -22374 -21852 -22365 -15948
rect -28287 -21861 -22365 -21852
rect -22258 -15972 -22211 -15908
rect -22147 -15972 -22131 -15908
rect -19059 -15939 -18955 -15561
rect -15939 -15592 -15892 -15528
rect -15828 -15592 -15812 -15528
rect -15649 -9648 -9727 -9639
rect -15649 -15552 -15640 -9648
rect -9736 -15552 -9727 -9648
rect -15649 -15561 -9727 -15552
rect -9620 -9672 -9573 -9608
rect -9509 -9672 -9493 -9608
rect -6421 -9639 -6317 -9261
rect -3301 -9292 -3254 -9228
rect -3190 -9292 -3174 -9228
rect -3011 -3348 2911 -3339
rect -3011 -9252 -3002 -3348
rect 2902 -9252 2911 -3348
rect -3011 -9261 2911 -9252
rect 3018 -3372 3065 -3308
rect 3129 -3372 3145 -3308
rect 6217 -3339 6321 -2961
rect 9337 -2992 9384 -2928
rect 9448 -2992 9464 -2928
rect 9627 2952 15549 2961
rect 9627 -2952 9636 2952
rect 15540 -2952 15549 2952
rect 9627 -2961 15549 -2952
rect 15656 2928 15703 2992
rect 15767 2928 15783 2992
rect 18855 2961 18959 3339
rect 21975 3308 22022 3372
rect 22086 3308 22102 3372
rect 22265 9252 28187 9261
rect 22265 3348 22274 9252
rect 28178 3348 28187 9252
rect 22265 3339 28187 3348
rect 28294 9228 28341 9292
rect 28405 9228 28421 9292
rect 31493 9261 31597 9639
rect 34613 9608 34660 9672
rect 34724 9608 34740 9672
rect 34903 15552 40825 15561
rect 34903 9648 34912 15552
rect 40816 9648 40825 15552
rect 34903 9639 40825 9648
rect 40932 15528 40979 15592
rect 41043 15528 41059 15592
rect 44131 15561 44235 15939
rect 47251 15908 47298 15972
rect 47362 15908 47378 15972
rect 47251 15892 47378 15908
rect 47251 15828 47298 15892
rect 47362 15828 47378 15892
rect 47251 15812 47378 15828
rect 47251 15688 47355 15812
rect 47251 15672 47378 15688
rect 47251 15608 47298 15672
rect 47362 15608 47378 15672
rect 47251 15592 47378 15608
rect 40932 15512 41059 15528
rect 40932 15448 40979 15512
rect 41043 15448 41059 15512
rect 40932 15432 41059 15448
rect 40932 15368 40979 15432
rect 41043 15368 41059 15432
rect 40932 15352 41059 15368
rect 40932 15288 40979 15352
rect 41043 15288 41059 15352
rect 40932 15272 41059 15288
rect 40932 15208 40979 15272
rect 41043 15208 41059 15272
rect 40932 15192 41059 15208
rect 40932 15128 40979 15192
rect 41043 15128 41059 15192
rect 40932 15112 41059 15128
rect 40932 15048 40979 15112
rect 41043 15048 41059 15112
rect 40932 15032 41059 15048
rect 40932 14968 40979 15032
rect 41043 14968 41059 15032
rect 40932 14952 41059 14968
rect 40932 14888 40979 14952
rect 41043 14888 41059 14952
rect 40932 14872 41059 14888
rect 40932 14808 40979 14872
rect 41043 14808 41059 14872
rect 40932 14792 41059 14808
rect 40932 14728 40979 14792
rect 41043 14728 41059 14792
rect 40932 14712 41059 14728
rect 40932 14648 40979 14712
rect 41043 14648 41059 14712
rect 40932 14632 41059 14648
rect 40932 14568 40979 14632
rect 41043 14568 41059 14632
rect 40932 14552 41059 14568
rect 40932 14488 40979 14552
rect 41043 14488 41059 14552
rect 40932 14472 41059 14488
rect 40932 14408 40979 14472
rect 41043 14408 41059 14472
rect 40932 14392 41059 14408
rect 40932 14328 40979 14392
rect 41043 14328 41059 14392
rect 40932 14312 41059 14328
rect 40932 14248 40979 14312
rect 41043 14248 41059 14312
rect 40932 14232 41059 14248
rect 40932 14168 40979 14232
rect 41043 14168 41059 14232
rect 40932 14152 41059 14168
rect 40932 14088 40979 14152
rect 41043 14088 41059 14152
rect 40932 14072 41059 14088
rect 40932 14008 40979 14072
rect 41043 14008 41059 14072
rect 40932 13992 41059 14008
rect 40932 13928 40979 13992
rect 41043 13928 41059 13992
rect 40932 13912 41059 13928
rect 40932 13848 40979 13912
rect 41043 13848 41059 13912
rect 40932 13832 41059 13848
rect 40932 13768 40979 13832
rect 41043 13768 41059 13832
rect 40932 13752 41059 13768
rect 40932 13688 40979 13752
rect 41043 13688 41059 13752
rect 40932 13672 41059 13688
rect 40932 13608 40979 13672
rect 41043 13608 41059 13672
rect 40932 13592 41059 13608
rect 40932 13528 40979 13592
rect 41043 13528 41059 13592
rect 40932 13512 41059 13528
rect 40932 13448 40979 13512
rect 41043 13448 41059 13512
rect 40932 13432 41059 13448
rect 40932 13368 40979 13432
rect 41043 13368 41059 13432
rect 40932 13352 41059 13368
rect 40932 13288 40979 13352
rect 41043 13288 41059 13352
rect 40932 13272 41059 13288
rect 40932 13208 40979 13272
rect 41043 13208 41059 13272
rect 40932 13192 41059 13208
rect 40932 13128 40979 13192
rect 41043 13128 41059 13192
rect 40932 13112 41059 13128
rect 40932 13048 40979 13112
rect 41043 13048 41059 13112
rect 40932 13032 41059 13048
rect 40932 12968 40979 13032
rect 41043 12968 41059 13032
rect 40932 12952 41059 12968
rect 40932 12888 40979 12952
rect 41043 12888 41059 12952
rect 40932 12872 41059 12888
rect 40932 12808 40979 12872
rect 41043 12808 41059 12872
rect 40932 12792 41059 12808
rect 40932 12728 40979 12792
rect 41043 12728 41059 12792
rect 40932 12712 41059 12728
rect 40932 12648 40979 12712
rect 41043 12648 41059 12712
rect 40932 12632 41059 12648
rect 40932 12568 40979 12632
rect 41043 12568 41059 12632
rect 40932 12552 41059 12568
rect 40932 12488 40979 12552
rect 41043 12488 41059 12552
rect 40932 12472 41059 12488
rect 40932 12408 40979 12472
rect 41043 12408 41059 12472
rect 40932 12392 41059 12408
rect 40932 12328 40979 12392
rect 41043 12328 41059 12392
rect 40932 12312 41059 12328
rect 40932 12248 40979 12312
rect 41043 12248 41059 12312
rect 40932 12232 41059 12248
rect 40932 12168 40979 12232
rect 41043 12168 41059 12232
rect 40932 12152 41059 12168
rect 40932 12088 40979 12152
rect 41043 12088 41059 12152
rect 40932 12072 41059 12088
rect 40932 12008 40979 12072
rect 41043 12008 41059 12072
rect 40932 11992 41059 12008
rect 40932 11928 40979 11992
rect 41043 11928 41059 11992
rect 40932 11912 41059 11928
rect 40932 11848 40979 11912
rect 41043 11848 41059 11912
rect 40932 11832 41059 11848
rect 40932 11768 40979 11832
rect 41043 11768 41059 11832
rect 40932 11752 41059 11768
rect 40932 11688 40979 11752
rect 41043 11688 41059 11752
rect 40932 11672 41059 11688
rect 40932 11608 40979 11672
rect 41043 11608 41059 11672
rect 40932 11592 41059 11608
rect 40932 11528 40979 11592
rect 41043 11528 41059 11592
rect 40932 11512 41059 11528
rect 40932 11448 40979 11512
rect 41043 11448 41059 11512
rect 40932 11432 41059 11448
rect 40932 11368 40979 11432
rect 41043 11368 41059 11432
rect 40932 11352 41059 11368
rect 40932 11288 40979 11352
rect 41043 11288 41059 11352
rect 40932 11272 41059 11288
rect 40932 11208 40979 11272
rect 41043 11208 41059 11272
rect 40932 11192 41059 11208
rect 40932 11128 40979 11192
rect 41043 11128 41059 11192
rect 40932 11112 41059 11128
rect 40932 11048 40979 11112
rect 41043 11048 41059 11112
rect 40932 11032 41059 11048
rect 40932 10968 40979 11032
rect 41043 10968 41059 11032
rect 40932 10952 41059 10968
rect 40932 10888 40979 10952
rect 41043 10888 41059 10952
rect 40932 10872 41059 10888
rect 40932 10808 40979 10872
rect 41043 10808 41059 10872
rect 40932 10792 41059 10808
rect 40932 10728 40979 10792
rect 41043 10728 41059 10792
rect 40932 10712 41059 10728
rect 40932 10648 40979 10712
rect 41043 10648 41059 10712
rect 40932 10632 41059 10648
rect 40932 10568 40979 10632
rect 41043 10568 41059 10632
rect 40932 10552 41059 10568
rect 40932 10488 40979 10552
rect 41043 10488 41059 10552
rect 40932 10472 41059 10488
rect 40932 10408 40979 10472
rect 41043 10408 41059 10472
rect 40932 10392 41059 10408
rect 40932 10328 40979 10392
rect 41043 10328 41059 10392
rect 40932 10312 41059 10328
rect 40932 10248 40979 10312
rect 41043 10248 41059 10312
rect 40932 10232 41059 10248
rect 40932 10168 40979 10232
rect 41043 10168 41059 10232
rect 40932 10152 41059 10168
rect 40932 10088 40979 10152
rect 41043 10088 41059 10152
rect 40932 10072 41059 10088
rect 40932 10008 40979 10072
rect 41043 10008 41059 10072
rect 40932 9992 41059 10008
rect 40932 9928 40979 9992
rect 41043 9928 41059 9992
rect 40932 9912 41059 9928
rect 40932 9848 40979 9912
rect 41043 9848 41059 9912
rect 40932 9832 41059 9848
rect 40932 9768 40979 9832
rect 41043 9768 41059 9832
rect 40932 9752 41059 9768
rect 40932 9688 40979 9752
rect 41043 9688 41059 9752
rect 40932 9672 41059 9688
rect 34613 9592 34740 9608
rect 34613 9528 34660 9592
rect 34724 9528 34740 9592
rect 34613 9512 34740 9528
rect 34613 9388 34717 9512
rect 34613 9372 34740 9388
rect 34613 9308 34660 9372
rect 34724 9308 34740 9372
rect 34613 9292 34740 9308
rect 28294 9212 28421 9228
rect 28294 9148 28341 9212
rect 28405 9148 28421 9212
rect 28294 9132 28421 9148
rect 28294 9068 28341 9132
rect 28405 9068 28421 9132
rect 28294 9052 28421 9068
rect 28294 8988 28341 9052
rect 28405 8988 28421 9052
rect 28294 8972 28421 8988
rect 28294 8908 28341 8972
rect 28405 8908 28421 8972
rect 28294 8892 28421 8908
rect 28294 8828 28341 8892
rect 28405 8828 28421 8892
rect 28294 8812 28421 8828
rect 28294 8748 28341 8812
rect 28405 8748 28421 8812
rect 28294 8732 28421 8748
rect 28294 8668 28341 8732
rect 28405 8668 28421 8732
rect 28294 8652 28421 8668
rect 28294 8588 28341 8652
rect 28405 8588 28421 8652
rect 28294 8572 28421 8588
rect 28294 8508 28341 8572
rect 28405 8508 28421 8572
rect 28294 8492 28421 8508
rect 28294 8428 28341 8492
rect 28405 8428 28421 8492
rect 28294 8412 28421 8428
rect 28294 8348 28341 8412
rect 28405 8348 28421 8412
rect 28294 8332 28421 8348
rect 28294 8268 28341 8332
rect 28405 8268 28421 8332
rect 28294 8252 28421 8268
rect 28294 8188 28341 8252
rect 28405 8188 28421 8252
rect 28294 8172 28421 8188
rect 28294 8108 28341 8172
rect 28405 8108 28421 8172
rect 28294 8092 28421 8108
rect 28294 8028 28341 8092
rect 28405 8028 28421 8092
rect 28294 8012 28421 8028
rect 28294 7948 28341 8012
rect 28405 7948 28421 8012
rect 28294 7932 28421 7948
rect 28294 7868 28341 7932
rect 28405 7868 28421 7932
rect 28294 7852 28421 7868
rect 28294 7788 28341 7852
rect 28405 7788 28421 7852
rect 28294 7772 28421 7788
rect 28294 7708 28341 7772
rect 28405 7708 28421 7772
rect 28294 7692 28421 7708
rect 28294 7628 28341 7692
rect 28405 7628 28421 7692
rect 28294 7612 28421 7628
rect 28294 7548 28341 7612
rect 28405 7548 28421 7612
rect 28294 7532 28421 7548
rect 28294 7468 28341 7532
rect 28405 7468 28421 7532
rect 28294 7452 28421 7468
rect 28294 7388 28341 7452
rect 28405 7388 28421 7452
rect 28294 7372 28421 7388
rect 28294 7308 28341 7372
rect 28405 7308 28421 7372
rect 28294 7292 28421 7308
rect 28294 7228 28341 7292
rect 28405 7228 28421 7292
rect 28294 7212 28421 7228
rect 28294 7148 28341 7212
rect 28405 7148 28421 7212
rect 28294 7132 28421 7148
rect 28294 7068 28341 7132
rect 28405 7068 28421 7132
rect 28294 7052 28421 7068
rect 28294 6988 28341 7052
rect 28405 6988 28421 7052
rect 28294 6972 28421 6988
rect 28294 6908 28341 6972
rect 28405 6908 28421 6972
rect 28294 6892 28421 6908
rect 28294 6828 28341 6892
rect 28405 6828 28421 6892
rect 28294 6812 28421 6828
rect 28294 6748 28341 6812
rect 28405 6748 28421 6812
rect 28294 6732 28421 6748
rect 28294 6668 28341 6732
rect 28405 6668 28421 6732
rect 28294 6652 28421 6668
rect 28294 6588 28341 6652
rect 28405 6588 28421 6652
rect 28294 6572 28421 6588
rect 28294 6508 28341 6572
rect 28405 6508 28421 6572
rect 28294 6492 28421 6508
rect 28294 6428 28341 6492
rect 28405 6428 28421 6492
rect 28294 6412 28421 6428
rect 28294 6348 28341 6412
rect 28405 6348 28421 6412
rect 28294 6332 28421 6348
rect 28294 6268 28341 6332
rect 28405 6268 28421 6332
rect 28294 6252 28421 6268
rect 28294 6188 28341 6252
rect 28405 6188 28421 6252
rect 28294 6172 28421 6188
rect 28294 6108 28341 6172
rect 28405 6108 28421 6172
rect 28294 6092 28421 6108
rect 28294 6028 28341 6092
rect 28405 6028 28421 6092
rect 28294 6012 28421 6028
rect 28294 5948 28341 6012
rect 28405 5948 28421 6012
rect 28294 5932 28421 5948
rect 28294 5868 28341 5932
rect 28405 5868 28421 5932
rect 28294 5852 28421 5868
rect 28294 5788 28341 5852
rect 28405 5788 28421 5852
rect 28294 5772 28421 5788
rect 28294 5708 28341 5772
rect 28405 5708 28421 5772
rect 28294 5692 28421 5708
rect 28294 5628 28341 5692
rect 28405 5628 28421 5692
rect 28294 5612 28421 5628
rect 28294 5548 28341 5612
rect 28405 5548 28421 5612
rect 28294 5532 28421 5548
rect 28294 5468 28341 5532
rect 28405 5468 28421 5532
rect 28294 5452 28421 5468
rect 28294 5388 28341 5452
rect 28405 5388 28421 5452
rect 28294 5372 28421 5388
rect 28294 5308 28341 5372
rect 28405 5308 28421 5372
rect 28294 5292 28421 5308
rect 28294 5228 28341 5292
rect 28405 5228 28421 5292
rect 28294 5212 28421 5228
rect 28294 5148 28341 5212
rect 28405 5148 28421 5212
rect 28294 5132 28421 5148
rect 28294 5068 28341 5132
rect 28405 5068 28421 5132
rect 28294 5052 28421 5068
rect 28294 4988 28341 5052
rect 28405 4988 28421 5052
rect 28294 4972 28421 4988
rect 28294 4908 28341 4972
rect 28405 4908 28421 4972
rect 28294 4892 28421 4908
rect 28294 4828 28341 4892
rect 28405 4828 28421 4892
rect 28294 4812 28421 4828
rect 28294 4748 28341 4812
rect 28405 4748 28421 4812
rect 28294 4732 28421 4748
rect 28294 4668 28341 4732
rect 28405 4668 28421 4732
rect 28294 4652 28421 4668
rect 28294 4588 28341 4652
rect 28405 4588 28421 4652
rect 28294 4572 28421 4588
rect 28294 4508 28341 4572
rect 28405 4508 28421 4572
rect 28294 4492 28421 4508
rect 28294 4428 28341 4492
rect 28405 4428 28421 4492
rect 28294 4412 28421 4428
rect 28294 4348 28341 4412
rect 28405 4348 28421 4412
rect 28294 4332 28421 4348
rect 28294 4268 28341 4332
rect 28405 4268 28421 4332
rect 28294 4252 28421 4268
rect 28294 4188 28341 4252
rect 28405 4188 28421 4252
rect 28294 4172 28421 4188
rect 28294 4108 28341 4172
rect 28405 4108 28421 4172
rect 28294 4092 28421 4108
rect 28294 4028 28341 4092
rect 28405 4028 28421 4092
rect 28294 4012 28421 4028
rect 28294 3948 28341 4012
rect 28405 3948 28421 4012
rect 28294 3932 28421 3948
rect 28294 3868 28341 3932
rect 28405 3868 28421 3932
rect 28294 3852 28421 3868
rect 28294 3788 28341 3852
rect 28405 3788 28421 3852
rect 28294 3772 28421 3788
rect 28294 3708 28341 3772
rect 28405 3708 28421 3772
rect 28294 3692 28421 3708
rect 28294 3628 28341 3692
rect 28405 3628 28421 3692
rect 28294 3612 28421 3628
rect 28294 3548 28341 3612
rect 28405 3548 28421 3612
rect 28294 3532 28421 3548
rect 28294 3468 28341 3532
rect 28405 3468 28421 3532
rect 28294 3452 28421 3468
rect 28294 3388 28341 3452
rect 28405 3388 28421 3452
rect 28294 3372 28421 3388
rect 21975 3292 22102 3308
rect 21975 3228 22022 3292
rect 22086 3228 22102 3292
rect 21975 3212 22102 3228
rect 21975 3088 22079 3212
rect 21975 3072 22102 3088
rect 21975 3008 22022 3072
rect 22086 3008 22102 3072
rect 21975 2992 22102 3008
rect 15656 2912 15783 2928
rect 15656 2848 15703 2912
rect 15767 2848 15783 2912
rect 15656 2832 15783 2848
rect 15656 2768 15703 2832
rect 15767 2768 15783 2832
rect 15656 2752 15783 2768
rect 15656 2688 15703 2752
rect 15767 2688 15783 2752
rect 15656 2672 15783 2688
rect 15656 2608 15703 2672
rect 15767 2608 15783 2672
rect 15656 2592 15783 2608
rect 15656 2528 15703 2592
rect 15767 2528 15783 2592
rect 15656 2512 15783 2528
rect 15656 2448 15703 2512
rect 15767 2448 15783 2512
rect 15656 2432 15783 2448
rect 15656 2368 15703 2432
rect 15767 2368 15783 2432
rect 15656 2352 15783 2368
rect 15656 2288 15703 2352
rect 15767 2288 15783 2352
rect 15656 2272 15783 2288
rect 15656 2208 15703 2272
rect 15767 2208 15783 2272
rect 15656 2192 15783 2208
rect 15656 2128 15703 2192
rect 15767 2128 15783 2192
rect 15656 2112 15783 2128
rect 15656 2048 15703 2112
rect 15767 2048 15783 2112
rect 15656 2032 15783 2048
rect 15656 1968 15703 2032
rect 15767 1968 15783 2032
rect 15656 1952 15783 1968
rect 15656 1888 15703 1952
rect 15767 1888 15783 1952
rect 15656 1872 15783 1888
rect 15656 1808 15703 1872
rect 15767 1808 15783 1872
rect 15656 1792 15783 1808
rect 15656 1728 15703 1792
rect 15767 1728 15783 1792
rect 15656 1712 15783 1728
rect 15656 1648 15703 1712
rect 15767 1648 15783 1712
rect 15656 1632 15783 1648
rect 15656 1568 15703 1632
rect 15767 1568 15783 1632
rect 15656 1552 15783 1568
rect 15656 1488 15703 1552
rect 15767 1488 15783 1552
rect 15656 1472 15783 1488
rect 15656 1408 15703 1472
rect 15767 1408 15783 1472
rect 15656 1392 15783 1408
rect 15656 1328 15703 1392
rect 15767 1328 15783 1392
rect 15656 1312 15783 1328
rect 15656 1248 15703 1312
rect 15767 1248 15783 1312
rect 15656 1232 15783 1248
rect 15656 1168 15703 1232
rect 15767 1168 15783 1232
rect 15656 1152 15783 1168
rect 15656 1088 15703 1152
rect 15767 1088 15783 1152
rect 15656 1072 15783 1088
rect 15656 1008 15703 1072
rect 15767 1008 15783 1072
rect 15656 992 15783 1008
rect 15656 928 15703 992
rect 15767 928 15783 992
rect 15656 912 15783 928
rect 15656 848 15703 912
rect 15767 848 15783 912
rect 15656 832 15783 848
rect 15656 768 15703 832
rect 15767 768 15783 832
rect 15656 752 15783 768
rect 15656 688 15703 752
rect 15767 688 15783 752
rect 15656 672 15783 688
rect 15656 608 15703 672
rect 15767 608 15783 672
rect 15656 592 15783 608
rect 15656 528 15703 592
rect 15767 528 15783 592
rect 15656 512 15783 528
rect 15656 448 15703 512
rect 15767 448 15783 512
rect 15656 432 15783 448
rect 15656 368 15703 432
rect 15767 368 15783 432
rect 15656 352 15783 368
rect 15656 288 15703 352
rect 15767 288 15783 352
rect 15656 272 15783 288
rect 15656 208 15703 272
rect 15767 208 15783 272
rect 15656 192 15783 208
rect 15656 128 15703 192
rect 15767 128 15783 192
rect 15656 112 15783 128
rect 15656 48 15703 112
rect 15767 48 15783 112
rect 15656 32 15783 48
rect 15656 -32 15703 32
rect 15767 -32 15783 32
rect 15656 -48 15783 -32
rect 15656 -112 15703 -48
rect 15767 -112 15783 -48
rect 15656 -128 15783 -112
rect 15656 -192 15703 -128
rect 15767 -192 15783 -128
rect 15656 -208 15783 -192
rect 15656 -272 15703 -208
rect 15767 -272 15783 -208
rect 15656 -288 15783 -272
rect 15656 -352 15703 -288
rect 15767 -352 15783 -288
rect 15656 -368 15783 -352
rect 15656 -432 15703 -368
rect 15767 -432 15783 -368
rect 15656 -448 15783 -432
rect 15656 -512 15703 -448
rect 15767 -512 15783 -448
rect 15656 -528 15783 -512
rect 15656 -592 15703 -528
rect 15767 -592 15783 -528
rect 15656 -608 15783 -592
rect 15656 -672 15703 -608
rect 15767 -672 15783 -608
rect 15656 -688 15783 -672
rect 15656 -752 15703 -688
rect 15767 -752 15783 -688
rect 15656 -768 15783 -752
rect 15656 -832 15703 -768
rect 15767 -832 15783 -768
rect 15656 -848 15783 -832
rect 15656 -912 15703 -848
rect 15767 -912 15783 -848
rect 15656 -928 15783 -912
rect 15656 -992 15703 -928
rect 15767 -992 15783 -928
rect 15656 -1008 15783 -992
rect 15656 -1072 15703 -1008
rect 15767 -1072 15783 -1008
rect 15656 -1088 15783 -1072
rect 15656 -1152 15703 -1088
rect 15767 -1152 15783 -1088
rect 15656 -1168 15783 -1152
rect 15656 -1232 15703 -1168
rect 15767 -1232 15783 -1168
rect 15656 -1248 15783 -1232
rect 15656 -1312 15703 -1248
rect 15767 -1312 15783 -1248
rect 15656 -1328 15783 -1312
rect 15656 -1392 15703 -1328
rect 15767 -1392 15783 -1328
rect 15656 -1408 15783 -1392
rect 15656 -1472 15703 -1408
rect 15767 -1472 15783 -1408
rect 15656 -1488 15783 -1472
rect 15656 -1552 15703 -1488
rect 15767 -1552 15783 -1488
rect 15656 -1568 15783 -1552
rect 15656 -1632 15703 -1568
rect 15767 -1632 15783 -1568
rect 15656 -1648 15783 -1632
rect 15656 -1712 15703 -1648
rect 15767 -1712 15783 -1648
rect 15656 -1728 15783 -1712
rect 15656 -1792 15703 -1728
rect 15767 -1792 15783 -1728
rect 15656 -1808 15783 -1792
rect 15656 -1872 15703 -1808
rect 15767 -1872 15783 -1808
rect 15656 -1888 15783 -1872
rect 15656 -1952 15703 -1888
rect 15767 -1952 15783 -1888
rect 15656 -1968 15783 -1952
rect 15656 -2032 15703 -1968
rect 15767 -2032 15783 -1968
rect 15656 -2048 15783 -2032
rect 15656 -2112 15703 -2048
rect 15767 -2112 15783 -2048
rect 15656 -2128 15783 -2112
rect 15656 -2192 15703 -2128
rect 15767 -2192 15783 -2128
rect 15656 -2208 15783 -2192
rect 15656 -2272 15703 -2208
rect 15767 -2272 15783 -2208
rect 15656 -2288 15783 -2272
rect 15656 -2352 15703 -2288
rect 15767 -2352 15783 -2288
rect 15656 -2368 15783 -2352
rect 15656 -2432 15703 -2368
rect 15767 -2432 15783 -2368
rect 15656 -2448 15783 -2432
rect 15656 -2512 15703 -2448
rect 15767 -2512 15783 -2448
rect 15656 -2528 15783 -2512
rect 15656 -2592 15703 -2528
rect 15767 -2592 15783 -2528
rect 15656 -2608 15783 -2592
rect 15656 -2672 15703 -2608
rect 15767 -2672 15783 -2608
rect 15656 -2688 15783 -2672
rect 15656 -2752 15703 -2688
rect 15767 -2752 15783 -2688
rect 15656 -2768 15783 -2752
rect 15656 -2832 15703 -2768
rect 15767 -2832 15783 -2768
rect 15656 -2848 15783 -2832
rect 15656 -2912 15703 -2848
rect 15767 -2912 15783 -2848
rect 15656 -2928 15783 -2912
rect 9337 -3008 9464 -2992
rect 9337 -3072 9384 -3008
rect 9448 -3072 9464 -3008
rect 9337 -3088 9464 -3072
rect 9337 -3212 9441 -3088
rect 9337 -3228 9464 -3212
rect 9337 -3292 9384 -3228
rect 9448 -3292 9464 -3228
rect 9337 -3308 9464 -3292
rect 3018 -3388 3145 -3372
rect 3018 -3452 3065 -3388
rect 3129 -3452 3145 -3388
rect 3018 -3468 3145 -3452
rect 3018 -3532 3065 -3468
rect 3129 -3532 3145 -3468
rect 3018 -3548 3145 -3532
rect 3018 -3612 3065 -3548
rect 3129 -3612 3145 -3548
rect 3018 -3628 3145 -3612
rect 3018 -3692 3065 -3628
rect 3129 -3692 3145 -3628
rect 3018 -3708 3145 -3692
rect 3018 -3772 3065 -3708
rect 3129 -3772 3145 -3708
rect 3018 -3788 3145 -3772
rect 3018 -3852 3065 -3788
rect 3129 -3852 3145 -3788
rect 3018 -3868 3145 -3852
rect 3018 -3932 3065 -3868
rect 3129 -3932 3145 -3868
rect 3018 -3948 3145 -3932
rect 3018 -4012 3065 -3948
rect 3129 -4012 3145 -3948
rect 3018 -4028 3145 -4012
rect 3018 -4092 3065 -4028
rect 3129 -4092 3145 -4028
rect 3018 -4108 3145 -4092
rect 3018 -4172 3065 -4108
rect 3129 -4172 3145 -4108
rect 3018 -4188 3145 -4172
rect 3018 -4252 3065 -4188
rect 3129 -4252 3145 -4188
rect 3018 -4268 3145 -4252
rect 3018 -4332 3065 -4268
rect 3129 -4332 3145 -4268
rect 3018 -4348 3145 -4332
rect 3018 -4412 3065 -4348
rect 3129 -4412 3145 -4348
rect 3018 -4428 3145 -4412
rect 3018 -4492 3065 -4428
rect 3129 -4492 3145 -4428
rect 3018 -4508 3145 -4492
rect 3018 -4572 3065 -4508
rect 3129 -4572 3145 -4508
rect 3018 -4588 3145 -4572
rect 3018 -4652 3065 -4588
rect 3129 -4652 3145 -4588
rect 3018 -4668 3145 -4652
rect 3018 -4732 3065 -4668
rect 3129 -4732 3145 -4668
rect 3018 -4748 3145 -4732
rect 3018 -4812 3065 -4748
rect 3129 -4812 3145 -4748
rect 3018 -4828 3145 -4812
rect 3018 -4892 3065 -4828
rect 3129 -4892 3145 -4828
rect 3018 -4908 3145 -4892
rect 3018 -4972 3065 -4908
rect 3129 -4972 3145 -4908
rect 3018 -4988 3145 -4972
rect 3018 -5052 3065 -4988
rect 3129 -5052 3145 -4988
rect 3018 -5068 3145 -5052
rect 3018 -5132 3065 -5068
rect 3129 -5132 3145 -5068
rect 3018 -5148 3145 -5132
rect 3018 -5212 3065 -5148
rect 3129 -5212 3145 -5148
rect 3018 -5228 3145 -5212
rect 3018 -5292 3065 -5228
rect 3129 -5292 3145 -5228
rect 3018 -5308 3145 -5292
rect 3018 -5372 3065 -5308
rect 3129 -5372 3145 -5308
rect 3018 -5388 3145 -5372
rect 3018 -5452 3065 -5388
rect 3129 -5452 3145 -5388
rect 3018 -5468 3145 -5452
rect 3018 -5532 3065 -5468
rect 3129 -5532 3145 -5468
rect 3018 -5548 3145 -5532
rect 3018 -5612 3065 -5548
rect 3129 -5612 3145 -5548
rect 3018 -5628 3145 -5612
rect 3018 -5692 3065 -5628
rect 3129 -5692 3145 -5628
rect 3018 -5708 3145 -5692
rect 3018 -5772 3065 -5708
rect 3129 -5772 3145 -5708
rect 3018 -5788 3145 -5772
rect 3018 -5852 3065 -5788
rect 3129 -5852 3145 -5788
rect 3018 -5868 3145 -5852
rect 3018 -5932 3065 -5868
rect 3129 -5932 3145 -5868
rect 3018 -5948 3145 -5932
rect 3018 -6012 3065 -5948
rect 3129 -6012 3145 -5948
rect 3018 -6028 3145 -6012
rect 3018 -6092 3065 -6028
rect 3129 -6092 3145 -6028
rect 3018 -6108 3145 -6092
rect 3018 -6172 3065 -6108
rect 3129 -6172 3145 -6108
rect 3018 -6188 3145 -6172
rect 3018 -6252 3065 -6188
rect 3129 -6252 3145 -6188
rect 3018 -6268 3145 -6252
rect 3018 -6332 3065 -6268
rect 3129 -6332 3145 -6268
rect 3018 -6348 3145 -6332
rect 3018 -6412 3065 -6348
rect 3129 -6412 3145 -6348
rect 3018 -6428 3145 -6412
rect 3018 -6492 3065 -6428
rect 3129 -6492 3145 -6428
rect 3018 -6508 3145 -6492
rect 3018 -6572 3065 -6508
rect 3129 -6572 3145 -6508
rect 3018 -6588 3145 -6572
rect 3018 -6652 3065 -6588
rect 3129 -6652 3145 -6588
rect 3018 -6668 3145 -6652
rect 3018 -6732 3065 -6668
rect 3129 -6732 3145 -6668
rect 3018 -6748 3145 -6732
rect 3018 -6812 3065 -6748
rect 3129 -6812 3145 -6748
rect 3018 -6828 3145 -6812
rect 3018 -6892 3065 -6828
rect 3129 -6892 3145 -6828
rect 3018 -6908 3145 -6892
rect 3018 -6972 3065 -6908
rect 3129 -6972 3145 -6908
rect 3018 -6988 3145 -6972
rect 3018 -7052 3065 -6988
rect 3129 -7052 3145 -6988
rect 3018 -7068 3145 -7052
rect 3018 -7132 3065 -7068
rect 3129 -7132 3145 -7068
rect 3018 -7148 3145 -7132
rect 3018 -7212 3065 -7148
rect 3129 -7212 3145 -7148
rect 3018 -7228 3145 -7212
rect 3018 -7292 3065 -7228
rect 3129 -7292 3145 -7228
rect 3018 -7308 3145 -7292
rect 3018 -7372 3065 -7308
rect 3129 -7372 3145 -7308
rect 3018 -7388 3145 -7372
rect 3018 -7452 3065 -7388
rect 3129 -7452 3145 -7388
rect 3018 -7468 3145 -7452
rect 3018 -7532 3065 -7468
rect 3129 -7532 3145 -7468
rect 3018 -7548 3145 -7532
rect 3018 -7612 3065 -7548
rect 3129 -7612 3145 -7548
rect 3018 -7628 3145 -7612
rect 3018 -7692 3065 -7628
rect 3129 -7692 3145 -7628
rect 3018 -7708 3145 -7692
rect 3018 -7772 3065 -7708
rect 3129 -7772 3145 -7708
rect 3018 -7788 3145 -7772
rect 3018 -7852 3065 -7788
rect 3129 -7852 3145 -7788
rect 3018 -7868 3145 -7852
rect 3018 -7932 3065 -7868
rect 3129 -7932 3145 -7868
rect 3018 -7948 3145 -7932
rect 3018 -8012 3065 -7948
rect 3129 -8012 3145 -7948
rect 3018 -8028 3145 -8012
rect 3018 -8092 3065 -8028
rect 3129 -8092 3145 -8028
rect 3018 -8108 3145 -8092
rect 3018 -8172 3065 -8108
rect 3129 -8172 3145 -8108
rect 3018 -8188 3145 -8172
rect 3018 -8252 3065 -8188
rect 3129 -8252 3145 -8188
rect 3018 -8268 3145 -8252
rect 3018 -8332 3065 -8268
rect 3129 -8332 3145 -8268
rect 3018 -8348 3145 -8332
rect 3018 -8412 3065 -8348
rect 3129 -8412 3145 -8348
rect 3018 -8428 3145 -8412
rect 3018 -8492 3065 -8428
rect 3129 -8492 3145 -8428
rect 3018 -8508 3145 -8492
rect 3018 -8572 3065 -8508
rect 3129 -8572 3145 -8508
rect 3018 -8588 3145 -8572
rect 3018 -8652 3065 -8588
rect 3129 -8652 3145 -8588
rect 3018 -8668 3145 -8652
rect 3018 -8732 3065 -8668
rect 3129 -8732 3145 -8668
rect 3018 -8748 3145 -8732
rect 3018 -8812 3065 -8748
rect 3129 -8812 3145 -8748
rect 3018 -8828 3145 -8812
rect 3018 -8892 3065 -8828
rect 3129 -8892 3145 -8828
rect 3018 -8908 3145 -8892
rect 3018 -8972 3065 -8908
rect 3129 -8972 3145 -8908
rect 3018 -8988 3145 -8972
rect 3018 -9052 3065 -8988
rect 3129 -9052 3145 -8988
rect 3018 -9068 3145 -9052
rect 3018 -9132 3065 -9068
rect 3129 -9132 3145 -9068
rect 3018 -9148 3145 -9132
rect 3018 -9212 3065 -9148
rect 3129 -9212 3145 -9148
rect 3018 -9228 3145 -9212
rect -3301 -9308 -3174 -9292
rect -3301 -9372 -3254 -9308
rect -3190 -9372 -3174 -9308
rect -3301 -9388 -3174 -9372
rect -3301 -9512 -3197 -9388
rect -3301 -9528 -3174 -9512
rect -3301 -9592 -3254 -9528
rect -3190 -9592 -3174 -9528
rect -3301 -9608 -3174 -9592
rect -9620 -9688 -9493 -9672
rect -9620 -9752 -9573 -9688
rect -9509 -9752 -9493 -9688
rect -9620 -9768 -9493 -9752
rect -9620 -9832 -9573 -9768
rect -9509 -9832 -9493 -9768
rect -9620 -9848 -9493 -9832
rect -9620 -9912 -9573 -9848
rect -9509 -9912 -9493 -9848
rect -9620 -9928 -9493 -9912
rect -9620 -9992 -9573 -9928
rect -9509 -9992 -9493 -9928
rect -9620 -10008 -9493 -9992
rect -9620 -10072 -9573 -10008
rect -9509 -10072 -9493 -10008
rect -9620 -10088 -9493 -10072
rect -9620 -10152 -9573 -10088
rect -9509 -10152 -9493 -10088
rect -9620 -10168 -9493 -10152
rect -9620 -10232 -9573 -10168
rect -9509 -10232 -9493 -10168
rect -9620 -10248 -9493 -10232
rect -9620 -10312 -9573 -10248
rect -9509 -10312 -9493 -10248
rect -9620 -10328 -9493 -10312
rect -9620 -10392 -9573 -10328
rect -9509 -10392 -9493 -10328
rect -9620 -10408 -9493 -10392
rect -9620 -10472 -9573 -10408
rect -9509 -10472 -9493 -10408
rect -9620 -10488 -9493 -10472
rect -9620 -10552 -9573 -10488
rect -9509 -10552 -9493 -10488
rect -9620 -10568 -9493 -10552
rect -9620 -10632 -9573 -10568
rect -9509 -10632 -9493 -10568
rect -9620 -10648 -9493 -10632
rect -9620 -10712 -9573 -10648
rect -9509 -10712 -9493 -10648
rect -9620 -10728 -9493 -10712
rect -9620 -10792 -9573 -10728
rect -9509 -10792 -9493 -10728
rect -9620 -10808 -9493 -10792
rect -9620 -10872 -9573 -10808
rect -9509 -10872 -9493 -10808
rect -9620 -10888 -9493 -10872
rect -9620 -10952 -9573 -10888
rect -9509 -10952 -9493 -10888
rect -9620 -10968 -9493 -10952
rect -9620 -11032 -9573 -10968
rect -9509 -11032 -9493 -10968
rect -9620 -11048 -9493 -11032
rect -9620 -11112 -9573 -11048
rect -9509 -11112 -9493 -11048
rect -9620 -11128 -9493 -11112
rect -9620 -11192 -9573 -11128
rect -9509 -11192 -9493 -11128
rect -9620 -11208 -9493 -11192
rect -9620 -11272 -9573 -11208
rect -9509 -11272 -9493 -11208
rect -9620 -11288 -9493 -11272
rect -9620 -11352 -9573 -11288
rect -9509 -11352 -9493 -11288
rect -9620 -11368 -9493 -11352
rect -9620 -11432 -9573 -11368
rect -9509 -11432 -9493 -11368
rect -9620 -11448 -9493 -11432
rect -9620 -11512 -9573 -11448
rect -9509 -11512 -9493 -11448
rect -9620 -11528 -9493 -11512
rect -9620 -11592 -9573 -11528
rect -9509 -11592 -9493 -11528
rect -9620 -11608 -9493 -11592
rect -9620 -11672 -9573 -11608
rect -9509 -11672 -9493 -11608
rect -9620 -11688 -9493 -11672
rect -9620 -11752 -9573 -11688
rect -9509 -11752 -9493 -11688
rect -9620 -11768 -9493 -11752
rect -9620 -11832 -9573 -11768
rect -9509 -11832 -9493 -11768
rect -9620 -11848 -9493 -11832
rect -9620 -11912 -9573 -11848
rect -9509 -11912 -9493 -11848
rect -9620 -11928 -9493 -11912
rect -9620 -11992 -9573 -11928
rect -9509 -11992 -9493 -11928
rect -9620 -12008 -9493 -11992
rect -9620 -12072 -9573 -12008
rect -9509 -12072 -9493 -12008
rect -9620 -12088 -9493 -12072
rect -9620 -12152 -9573 -12088
rect -9509 -12152 -9493 -12088
rect -9620 -12168 -9493 -12152
rect -9620 -12232 -9573 -12168
rect -9509 -12232 -9493 -12168
rect -9620 -12248 -9493 -12232
rect -9620 -12312 -9573 -12248
rect -9509 -12312 -9493 -12248
rect -9620 -12328 -9493 -12312
rect -9620 -12392 -9573 -12328
rect -9509 -12392 -9493 -12328
rect -9620 -12408 -9493 -12392
rect -9620 -12472 -9573 -12408
rect -9509 -12472 -9493 -12408
rect -9620 -12488 -9493 -12472
rect -9620 -12552 -9573 -12488
rect -9509 -12552 -9493 -12488
rect -9620 -12568 -9493 -12552
rect -9620 -12632 -9573 -12568
rect -9509 -12632 -9493 -12568
rect -9620 -12648 -9493 -12632
rect -9620 -12712 -9573 -12648
rect -9509 -12712 -9493 -12648
rect -9620 -12728 -9493 -12712
rect -9620 -12792 -9573 -12728
rect -9509 -12792 -9493 -12728
rect -9620 -12808 -9493 -12792
rect -9620 -12872 -9573 -12808
rect -9509 -12872 -9493 -12808
rect -9620 -12888 -9493 -12872
rect -9620 -12952 -9573 -12888
rect -9509 -12952 -9493 -12888
rect -9620 -12968 -9493 -12952
rect -9620 -13032 -9573 -12968
rect -9509 -13032 -9493 -12968
rect -9620 -13048 -9493 -13032
rect -9620 -13112 -9573 -13048
rect -9509 -13112 -9493 -13048
rect -9620 -13128 -9493 -13112
rect -9620 -13192 -9573 -13128
rect -9509 -13192 -9493 -13128
rect -9620 -13208 -9493 -13192
rect -9620 -13272 -9573 -13208
rect -9509 -13272 -9493 -13208
rect -9620 -13288 -9493 -13272
rect -9620 -13352 -9573 -13288
rect -9509 -13352 -9493 -13288
rect -9620 -13368 -9493 -13352
rect -9620 -13432 -9573 -13368
rect -9509 -13432 -9493 -13368
rect -9620 -13448 -9493 -13432
rect -9620 -13512 -9573 -13448
rect -9509 -13512 -9493 -13448
rect -9620 -13528 -9493 -13512
rect -9620 -13592 -9573 -13528
rect -9509 -13592 -9493 -13528
rect -9620 -13608 -9493 -13592
rect -9620 -13672 -9573 -13608
rect -9509 -13672 -9493 -13608
rect -9620 -13688 -9493 -13672
rect -9620 -13752 -9573 -13688
rect -9509 -13752 -9493 -13688
rect -9620 -13768 -9493 -13752
rect -9620 -13832 -9573 -13768
rect -9509 -13832 -9493 -13768
rect -9620 -13848 -9493 -13832
rect -9620 -13912 -9573 -13848
rect -9509 -13912 -9493 -13848
rect -9620 -13928 -9493 -13912
rect -9620 -13992 -9573 -13928
rect -9509 -13992 -9493 -13928
rect -9620 -14008 -9493 -13992
rect -9620 -14072 -9573 -14008
rect -9509 -14072 -9493 -14008
rect -9620 -14088 -9493 -14072
rect -9620 -14152 -9573 -14088
rect -9509 -14152 -9493 -14088
rect -9620 -14168 -9493 -14152
rect -9620 -14232 -9573 -14168
rect -9509 -14232 -9493 -14168
rect -9620 -14248 -9493 -14232
rect -9620 -14312 -9573 -14248
rect -9509 -14312 -9493 -14248
rect -9620 -14328 -9493 -14312
rect -9620 -14392 -9573 -14328
rect -9509 -14392 -9493 -14328
rect -9620 -14408 -9493 -14392
rect -9620 -14472 -9573 -14408
rect -9509 -14472 -9493 -14408
rect -9620 -14488 -9493 -14472
rect -9620 -14552 -9573 -14488
rect -9509 -14552 -9493 -14488
rect -9620 -14568 -9493 -14552
rect -9620 -14632 -9573 -14568
rect -9509 -14632 -9493 -14568
rect -9620 -14648 -9493 -14632
rect -9620 -14712 -9573 -14648
rect -9509 -14712 -9493 -14648
rect -9620 -14728 -9493 -14712
rect -9620 -14792 -9573 -14728
rect -9509 -14792 -9493 -14728
rect -9620 -14808 -9493 -14792
rect -9620 -14872 -9573 -14808
rect -9509 -14872 -9493 -14808
rect -9620 -14888 -9493 -14872
rect -9620 -14952 -9573 -14888
rect -9509 -14952 -9493 -14888
rect -9620 -14968 -9493 -14952
rect -9620 -15032 -9573 -14968
rect -9509 -15032 -9493 -14968
rect -9620 -15048 -9493 -15032
rect -9620 -15112 -9573 -15048
rect -9509 -15112 -9493 -15048
rect -9620 -15128 -9493 -15112
rect -9620 -15192 -9573 -15128
rect -9509 -15192 -9493 -15128
rect -9620 -15208 -9493 -15192
rect -9620 -15272 -9573 -15208
rect -9509 -15272 -9493 -15208
rect -9620 -15288 -9493 -15272
rect -9620 -15352 -9573 -15288
rect -9509 -15352 -9493 -15288
rect -9620 -15368 -9493 -15352
rect -9620 -15432 -9573 -15368
rect -9509 -15432 -9493 -15368
rect -9620 -15448 -9493 -15432
rect -9620 -15512 -9573 -15448
rect -9509 -15512 -9493 -15448
rect -9620 -15528 -9493 -15512
rect -15939 -15608 -15812 -15592
rect -15939 -15672 -15892 -15608
rect -15828 -15672 -15812 -15608
rect -15939 -15688 -15812 -15672
rect -15939 -15812 -15835 -15688
rect -15939 -15828 -15812 -15812
rect -15939 -15892 -15892 -15828
rect -15828 -15892 -15812 -15828
rect -15939 -15908 -15812 -15892
rect -22258 -15988 -22131 -15972
rect -22258 -16052 -22211 -15988
rect -22147 -16052 -22131 -15988
rect -22258 -16068 -22131 -16052
rect -22258 -16132 -22211 -16068
rect -22147 -16132 -22131 -16068
rect -22258 -16148 -22131 -16132
rect -22258 -16212 -22211 -16148
rect -22147 -16212 -22131 -16148
rect -22258 -16228 -22131 -16212
rect -22258 -16292 -22211 -16228
rect -22147 -16292 -22131 -16228
rect -22258 -16308 -22131 -16292
rect -22258 -16372 -22211 -16308
rect -22147 -16372 -22131 -16308
rect -22258 -16388 -22131 -16372
rect -22258 -16452 -22211 -16388
rect -22147 -16452 -22131 -16388
rect -22258 -16468 -22131 -16452
rect -22258 -16532 -22211 -16468
rect -22147 -16532 -22131 -16468
rect -22258 -16548 -22131 -16532
rect -22258 -16612 -22211 -16548
rect -22147 -16612 -22131 -16548
rect -22258 -16628 -22131 -16612
rect -22258 -16692 -22211 -16628
rect -22147 -16692 -22131 -16628
rect -22258 -16708 -22131 -16692
rect -22258 -16772 -22211 -16708
rect -22147 -16772 -22131 -16708
rect -22258 -16788 -22131 -16772
rect -22258 -16852 -22211 -16788
rect -22147 -16852 -22131 -16788
rect -22258 -16868 -22131 -16852
rect -22258 -16932 -22211 -16868
rect -22147 -16932 -22131 -16868
rect -22258 -16948 -22131 -16932
rect -22258 -17012 -22211 -16948
rect -22147 -17012 -22131 -16948
rect -22258 -17028 -22131 -17012
rect -22258 -17092 -22211 -17028
rect -22147 -17092 -22131 -17028
rect -22258 -17108 -22131 -17092
rect -22258 -17172 -22211 -17108
rect -22147 -17172 -22131 -17108
rect -22258 -17188 -22131 -17172
rect -22258 -17252 -22211 -17188
rect -22147 -17252 -22131 -17188
rect -22258 -17268 -22131 -17252
rect -22258 -17332 -22211 -17268
rect -22147 -17332 -22131 -17268
rect -22258 -17348 -22131 -17332
rect -22258 -17412 -22211 -17348
rect -22147 -17412 -22131 -17348
rect -22258 -17428 -22131 -17412
rect -22258 -17492 -22211 -17428
rect -22147 -17492 -22131 -17428
rect -22258 -17508 -22131 -17492
rect -22258 -17572 -22211 -17508
rect -22147 -17572 -22131 -17508
rect -22258 -17588 -22131 -17572
rect -22258 -17652 -22211 -17588
rect -22147 -17652 -22131 -17588
rect -22258 -17668 -22131 -17652
rect -22258 -17732 -22211 -17668
rect -22147 -17732 -22131 -17668
rect -22258 -17748 -22131 -17732
rect -22258 -17812 -22211 -17748
rect -22147 -17812 -22131 -17748
rect -22258 -17828 -22131 -17812
rect -22258 -17892 -22211 -17828
rect -22147 -17892 -22131 -17828
rect -22258 -17908 -22131 -17892
rect -22258 -17972 -22211 -17908
rect -22147 -17972 -22131 -17908
rect -22258 -17988 -22131 -17972
rect -22258 -18052 -22211 -17988
rect -22147 -18052 -22131 -17988
rect -22258 -18068 -22131 -18052
rect -22258 -18132 -22211 -18068
rect -22147 -18132 -22131 -18068
rect -22258 -18148 -22131 -18132
rect -22258 -18212 -22211 -18148
rect -22147 -18212 -22131 -18148
rect -22258 -18228 -22131 -18212
rect -22258 -18292 -22211 -18228
rect -22147 -18292 -22131 -18228
rect -22258 -18308 -22131 -18292
rect -22258 -18372 -22211 -18308
rect -22147 -18372 -22131 -18308
rect -22258 -18388 -22131 -18372
rect -22258 -18452 -22211 -18388
rect -22147 -18452 -22131 -18388
rect -22258 -18468 -22131 -18452
rect -22258 -18532 -22211 -18468
rect -22147 -18532 -22131 -18468
rect -22258 -18548 -22131 -18532
rect -22258 -18612 -22211 -18548
rect -22147 -18612 -22131 -18548
rect -22258 -18628 -22131 -18612
rect -22258 -18692 -22211 -18628
rect -22147 -18692 -22131 -18628
rect -22258 -18708 -22131 -18692
rect -22258 -18772 -22211 -18708
rect -22147 -18772 -22131 -18708
rect -22258 -18788 -22131 -18772
rect -22258 -18852 -22211 -18788
rect -22147 -18852 -22131 -18788
rect -22258 -18868 -22131 -18852
rect -22258 -18932 -22211 -18868
rect -22147 -18932 -22131 -18868
rect -22258 -18948 -22131 -18932
rect -22258 -19012 -22211 -18948
rect -22147 -19012 -22131 -18948
rect -22258 -19028 -22131 -19012
rect -22258 -19092 -22211 -19028
rect -22147 -19092 -22131 -19028
rect -22258 -19108 -22131 -19092
rect -22258 -19172 -22211 -19108
rect -22147 -19172 -22131 -19108
rect -22258 -19188 -22131 -19172
rect -22258 -19252 -22211 -19188
rect -22147 -19252 -22131 -19188
rect -22258 -19268 -22131 -19252
rect -22258 -19332 -22211 -19268
rect -22147 -19332 -22131 -19268
rect -22258 -19348 -22131 -19332
rect -22258 -19412 -22211 -19348
rect -22147 -19412 -22131 -19348
rect -22258 -19428 -22131 -19412
rect -22258 -19492 -22211 -19428
rect -22147 -19492 -22131 -19428
rect -22258 -19508 -22131 -19492
rect -22258 -19572 -22211 -19508
rect -22147 -19572 -22131 -19508
rect -22258 -19588 -22131 -19572
rect -22258 -19652 -22211 -19588
rect -22147 -19652 -22131 -19588
rect -22258 -19668 -22131 -19652
rect -22258 -19732 -22211 -19668
rect -22147 -19732 -22131 -19668
rect -22258 -19748 -22131 -19732
rect -22258 -19812 -22211 -19748
rect -22147 -19812 -22131 -19748
rect -22258 -19828 -22131 -19812
rect -22258 -19892 -22211 -19828
rect -22147 -19892 -22131 -19828
rect -22258 -19908 -22131 -19892
rect -22258 -19972 -22211 -19908
rect -22147 -19972 -22131 -19908
rect -22258 -19988 -22131 -19972
rect -22258 -20052 -22211 -19988
rect -22147 -20052 -22131 -19988
rect -22258 -20068 -22131 -20052
rect -22258 -20132 -22211 -20068
rect -22147 -20132 -22131 -20068
rect -22258 -20148 -22131 -20132
rect -22258 -20212 -22211 -20148
rect -22147 -20212 -22131 -20148
rect -22258 -20228 -22131 -20212
rect -22258 -20292 -22211 -20228
rect -22147 -20292 -22131 -20228
rect -22258 -20308 -22131 -20292
rect -22258 -20372 -22211 -20308
rect -22147 -20372 -22131 -20308
rect -22258 -20388 -22131 -20372
rect -22258 -20452 -22211 -20388
rect -22147 -20452 -22131 -20388
rect -22258 -20468 -22131 -20452
rect -22258 -20532 -22211 -20468
rect -22147 -20532 -22131 -20468
rect -22258 -20548 -22131 -20532
rect -22258 -20612 -22211 -20548
rect -22147 -20612 -22131 -20548
rect -22258 -20628 -22131 -20612
rect -22258 -20692 -22211 -20628
rect -22147 -20692 -22131 -20628
rect -22258 -20708 -22131 -20692
rect -22258 -20772 -22211 -20708
rect -22147 -20772 -22131 -20708
rect -22258 -20788 -22131 -20772
rect -22258 -20852 -22211 -20788
rect -22147 -20852 -22131 -20788
rect -22258 -20868 -22131 -20852
rect -22258 -20932 -22211 -20868
rect -22147 -20932 -22131 -20868
rect -22258 -20948 -22131 -20932
rect -22258 -21012 -22211 -20948
rect -22147 -21012 -22131 -20948
rect -22258 -21028 -22131 -21012
rect -22258 -21092 -22211 -21028
rect -22147 -21092 -22131 -21028
rect -22258 -21108 -22131 -21092
rect -22258 -21172 -22211 -21108
rect -22147 -21172 -22131 -21108
rect -22258 -21188 -22131 -21172
rect -22258 -21252 -22211 -21188
rect -22147 -21252 -22131 -21188
rect -22258 -21268 -22131 -21252
rect -22258 -21332 -22211 -21268
rect -22147 -21332 -22131 -21268
rect -22258 -21348 -22131 -21332
rect -22258 -21412 -22211 -21348
rect -22147 -21412 -22131 -21348
rect -22258 -21428 -22131 -21412
rect -22258 -21492 -22211 -21428
rect -22147 -21492 -22131 -21428
rect -22258 -21508 -22131 -21492
rect -22258 -21572 -22211 -21508
rect -22147 -21572 -22131 -21508
rect -22258 -21588 -22131 -21572
rect -22258 -21652 -22211 -21588
rect -22147 -21652 -22131 -21588
rect -22258 -21668 -22131 -21652
rect -22258 -21732 -22211 -21668
rect -22147 -21732 -22131 -21668
rect -22258 -21748 -22131 -21732
rect -22258 -21812 -22211 -21748
rect -22147 -21812 -22131 -21748
rect -22258 -21828 -22131 -21812
rect -28577 -21908 -28450 -21892
rect -28577 -21972 -28530 -21908
rect -28466 -21972 -28450 -21908
rect -28577 -21988 -28450 -21972
rect -28577 -22112 -28473 -21988
rect -28577 -22128 -28450 -22112
rect -28577 -22192 -28530 -22128
rect -28466 -22192 -28450 -22128
rect -28577 -22208 -28450 -22192
rect -34896 -22288 -34769 -22272
rect -34896 -22352 -34849 -22288
rect -34785 -22352 -34769 -22288
rect -34896 -22368 -34769 -22352
rect -34896 -22432 -34849 -22368
rect -34785 -22432 -34769 -22368
rect -34896 -22448 -34769 -22432
rect -34896 -22512 -34849 -22448
rect -34785 -22512 -34769 -22448
rect -34896 -22528 -34769 -22512
rect -34896 -22592 -34849 -22528
rect -34785 -22592 -34769 -22528
rect -34896 -22608 -34769 -22592
rect -34896 -22672 -34849 -22608
rect -34785 -22672 -34769 -22608
rect -34896 -22688 -34769 -22672
rect -34896 -22752 -34849 -22688
rect -34785 -22752 -34769 -22688
rect -34896 -22768 -34769 -22752
rect -34896 -22832 -34849 -22768
rect -34785 -22832 -34769 -22768
rect -34896 -22848 -34769 -22832
rect -34896 -22912 -34849 -22848
rect -34785 -22912 -34769 -22848
rect -34896 -22928 -34769 -22912
rect -34896 -22992 -34849 -22928
rect -34785 -22992 -34769 -22928
rect -34896 -23008 -34769 -22992
rect -34896 -23072 -34849 -23008
rect -34785 -23072 -34769 -23008
rect -34896 -23088 -34769 -23072
rect -34896 -23152 -34849 -23088
rect -34785 -23152 -34769 -23088
rect -34896 -23168 -34769 -23152
rect -34896 -23232 -34849 -23168
rect -34785 -23232 -34769 -23168
rect -34896 -23248 -34769 -23232
rect -34896 -23312 -34849 -23248
rect -34785 -23312 -34769 -23248
rect -34896 -23328 -34769 -23312
rect -34896 -23392 -34849 -23328
rect -34785 -23392 -34769 -23328
rect -34896 -23408 -34769 -23392
rect -34896 -23472 -34849 -23408
rect -34785 -23472 -34769 -23408
rect -34896 -23488 -34769 -23472
rect -34896 -23552 -34849 -23488
rect -34785 -23552 -34769 -23488
rect -34896 -23568 -34769 -23552
rect -34896 -23632 -34849 -23568
rect -34785 -23632 -34769 -23568
rect -34896 -23648 -34769 -23632
rect -34896 -23712 -34849 -23648
rect -34785 -23712 -34769 -23648
rect -34896 -23728 -34769 -23712
rect -34896 -23792 -34849 -23728
rect -34785 -23792 -34769 -23728
rect -34896 -23808 -34769 -23792
rect -34896 -23872 -34849 -23808
rect -34785 -23872 -34769 -23808
rect -34896 -23888 -34769 -23872
rect -34896 -23952 -34849 -23888
rect -34785 -23952 -34769 -23888
rect -34896 -23968 -34769 -23952
rect -34896 -24032 -34849 -23968
rect -34785 -24032 -34769 -23968
rect -34896 -24048 -34769 -24032
rect -34896 -24112 -34849 -24048
rect -34785 -24112 -34769 -24048
rect -34896 -24128 -34769 -24112
rect -34896 -24192 -34849 -24128
rect -34785 -24192 -34769 -24128
rect -34896 -24208 -34769 -24192
rect -34896 -24272 -34849 -24208
rect -34785 -24272 -34769 -24208
rect -34896 -24288 -34769 -24272
rect -34896 -24352 -34849 -24288
rect -34785 -24352 -34769 -24288
rect -34896 -24368 -34769 -24352
rect -34896 -24432 -34849 -24368
rect -34785 -24432 -34769 -24368
rect -34896 -24448 -34769 -24432
rect -34896 -24512 -34849 -24448
rect -34785 -24512 -34769 -24448
rect -34896 -24528 -34769 -24512
rect -34896 -24592 -34849 -24528
rect -34785 -24592 -34769 -24528
rect -34896 -24608 -34769 -24592
rect -34896 -24672 -34849 -24608
rect -34785 -24672 -34769 -24608
rect -34896 -24688 -34769 -24672
rect -34896 -24752 -34849 -24688
rect -34785 -24752 -34769 -24688
rect -34896 -24768 -34769 -24752
rect -34896 -24832 -34849 -24768
rect -34785 -24832 -34769 -24768
rect -34896 -24848 -34769 -24832
rect -34896 -24912 -34849 -24848
rect -34785 -24912 -34769 -24848
rect -34896 -24928 -34769 -24912
rect -34896 -24992 -34849 -24928
rect -34785 -24992 -34769 -24928
rect -34896 -25008 -34769 -24992
rect -34896 -25072 -34849 -25008
rect -34785 -25072 -34769 -25008
rect -34896 -25088 -34769 -25072
rect -34896 -25152 -34849 -25088
rect -34785 -25152 -34769 -25088
rect -34896 -25168 -34769 -25152
rect -34896 -25232 -34849 -25168
rect -34785 -25232 -34769 -25168
rect -34896 -25248 -34769 -25232
rect -34896 -25312 -34849 -25248
rect -34785 -25312 -34769 -25248
rect -34896 -25328 -34769 -25312
rect -34896 -25392 -34849 -25328
rect -34785 -25392 -34769 -25328
rect -34896 -25408 -34769 -25392
rect -34896 -25472 -34849 -25408
rect -34785 -25472 -34769 -25408
rect -34896 -25488 -34769 -25472
rect -34896 -25552 -34849 -25488
rect -34785 -25552 -34769 -25488
rect -34896 -25568 -34769 -25552
rect -34896 -25632 -34849 -25568
rect -34785 -25632 -34769 -25568
rect -34896 -25648 -34769 -25632
rect -34896 -25712 -34849 -25648
rect -34785 -25712 -34769 -25648
rect -34896 -25728 -34769 -25712
rect -34896 -25792 -34849 -25728
rect -34785 -25792 -34769 -25728
rect -34896 -25808 -34769 -25792
rect -34896 -25872 -34849 -25808
rect -34785 -25872 -34769 -25808
rect -34896 -25888 -34769 -25872
rect -34896 -25952 -34849 -25888
rect -34785 -25952 -34769 -25888
rect -34896 -25968 -34769 -25952
rect -34896 -26032 -34849 -25968
rect -34785 -26032 -34769 -25968
rect -34896 -26048 -34769 -26032
rect -34896 -26112 -34849 -26048
rect -34785 -26112 -34769 -26048
rect -34896 -26128 -34769 -26112
rect -34896 -26192 -34849 -26128
rect -34785 -26192 -34769 -26128
rect -34896 -26208 -34769 -26192
rect -34896 -26272 -34849 -26208
rect -34785 -26272 -34769 -26208
rect -34896 -26288 -34769 -26272
rect -34896 -26352 -34849 -26288
rect -34785 -26352 -34769 -26288
rect -34896 -26368 -34769 -26352
rect -34896 -26432 -34849 -26368
rect -34785 -26432 -34769 -26368
rect -34896 -26448 -34769 -26432
rect -34896 -26512 -34849 -26448
rect -34785 -26512 -34769 -26448
rect -34896 -26528 -34769 -26512
rect -34896 -26592 -34849 -26528
rect -34785 -26592 -34769 -26528
rect -34896 -26608 -34769 -26592
rect -34896 -26672 -34849 -26608
rect -34785 -26672 -34769 -26608
rect -34896 -26688 -34769 -26672
rect -34896 -26752 -34849 -26688
rect -34785 -26752 -34769 -26688
rect -34896 -26768 -34769 -26752
rect -34896 -26832 -34849 -26768
rect -34785 -26832 -34769 -26768
rect -34896 -26848 -34769 -26832
rect -34896 -26912 -34849 -26848
rect -34785 -26912 -34769 -26848
rect -34896 -26928 -34769 -26912
rect -34896 -26992 -34849 -26928
rect -34785 -26992 -34769 -26928
rect -34896 -27008 -34769 -26992
rect -34896 -27072 -34849 -27008
rect -34785 -27072 -34769 -27008
rect -34896 -27088 -34769 -27072
rect -34896 -27152 -34849 -27088
rect -34785 -27152 -34769 -27088
rect -34896 -27168 -34769 -27152
rect -34896 -27232 -34849 -27168
rect -34785 -27232 -34769 -27168
rect -34896 -27248 -34769 -27232
rect -34896 -27312 -34849 -27248
rect -34785 -27312 -34769 -27248
rect -34896 -27328 -34769 -27312
rect -34896 -27392 -34849 -27328
rect -34785 -27392 -34769 -27328
rect -34896 -27408 -34769 -27392
rect -34896 -27472 -34849 -27408
rect -34785 -27472 -34769 -27408
rect -34896 -27488 -34769 -27472
rect -34896 -27552 -34849 -27488
rect -34785 -27552 -34769 -27488
rect -34896 -27568 -34769 -27552
rect -34896 -27632 -34849 -27568
rect -34785 -27632 -34769 -27568
rect -34896 -27648 -34769 -27632
rect -34896 -27712 -34849 -27648
rect -34785 -27712 -34769 -27648
rect -34896 -27728 -34769 -27712
rect -34896 -27792 -34849 -27728
rect -34785 -27792 -34769 -27728
rect -34896 -27808 -34769 -27792
rect -34896 -27872 -34849 -27808
rect -34785 -27872 -34769 -27808
rect -34896 -27888 -34769 -27872
rect -34896 -27952 -34849 -27888
rect -34785 -27952 -34769 -27888
rect -34896 -27968 -34769 -27952
rect -34896 -28032 -34849 -27968
rect -34785 -28032 -34769 -27968
rect -34896 -28048 -34769 -28032
rect -34896 -28112 -34849 -28048
rect -34785 -28112 -34769 -28048
rect -34896 -28128 -34769 -28112
rect -41215 -28208 -41088 -28192
rect -41215 -28272 -41168 -28208
rect -41104 -28272 -41088 -28208
rect -41215 -28288 -41088 -28272
rect -41215 -28412 -41111 -28288
rect -41215 -28428 -41088 -28412
rect -41215 -28492 -41168 -28428
rect -41104 -28492 -41088 -28428
rect -41215 -28508 -41088 -28492
rect -47244 -28548 -41322 -28539
rect -47244 -34452 -47235 -28548
rect -41331 -34452 -41322 -28548
rect -47244 -34461 -41322 -34452
rect -41215 -28572 -41168 -28508
rect -41104 -28572 -41088 -28508
rect -38016 -28539 -37912 -28161
rect -34896 -28192 -34849 -28128
rect -34785 -28192 -34769 -28128
rect -34606 -22248 -28684 -22239
rect -34606 -28152 -34597 -22248
rect -28693 -28152 -28684 -22248
rect -34606 -28161 -28684 -28152
rect -28577 -22272 -28530 -22208
rect -28466 -22272 -28450 -22208
rect -25378 -22239 -25274 -21861
rect -22258 -21892 -22211 -21828
rect -22147 -21892 -22131 -21828
rect -21968 -15948 -16046 -15939
rect -21968 -21852 -21959 -15948
rect -16055 -21852 -16046 -15948
rect -21968 -21861 -16046 -21852
rect -15939 -15972 -15892 -15908
rect -15828 -15972 -15812 -15908
rect -12740 -15939 -12636 -15561
rect -9620 -15592 -9573 -15528
rect -9509 -15592 -9493 -15528
rect -9330 -9648 -3408 -9639
rect -9330 -15552 -9321 -9648
rect -3417 -15552 -3408 -9648
rect -9330 -15561 -3408 -15552
rect -3301 -9672 -3254 -9608
rect -3190 -9672 -3174 -9608
rect -102 -9639 2 -9261
rect 3018 -9292 3065 -9228
rect 3129 -9292 3145 -9228
rect 3308 -3348 9230 -3339
rect 3308 -9252 3317 -3348
rect 9221 -9252 9230 -3348
rect 3308 -9261 9230 -9252
rect 9337 -3372 9384 -3308
rect 9448 -3372 9464 -3308
rect 12536 -3339 12640 -2961
rect 15656 -2992 15703 -2928
rect 15767 -2992 15783 -2928
rect 15946 2952 21868 2961
rect 15946 -2952 15955 2952
rect 21859 -2952 21868 2952
rect 15946 -2961 21868 -2952
rect 21975 2928 22022 2992
rect 22086 2928 22102 2992
rect 25174 2961 25278 3339
rect 28294 3308 28341 3372
rect 28405 3308 28421 3372
rect 28584 9252 34506 9261
rect 28584 3348 28593 9252
rect 34497 3348 34506 9252
rect 28584 3339 34506 3348
rect 34613 9228 34660 9292
rect 34724 9228 34740 9292
rect 37812 9261 37916 9639
rect 40932 9608 40979 9672
rect 41043 9608 41059 9672
rect 41222 15552 47144 15561
rect 41222 9648 41231 15552
rect 47135 9648 47144 15552
rect 41222 9639 47144 9648
rect 47251 15528 47298 15592
rect 47362 15528 47378 15592
rect 47251 15512 47378 15528
rect 47251 15448 47298 15512
rect 47362 15448 47378 15512
rect 47251 15432 47378 15448
rect 47251 15368 47298 15432
rect 47362 15368 47378 15432
rect 47251 15352 47378 15368
rect 47251 15288 47298 15352
rect 47362 15288 47378 15352
rect 47251 15272 47378 15288
rect 47251 15208 47298 15272
rect 47362 15208 47378 15272
rect 47251 15192 47378 15208
rect 47251 15128 47298 15192
rect 47362 15128 47378 15192
rect 47251 15112 47378 15128
rect 47251 15048 47298 15112
rect 47362 15048 47378 15112
rect 47251 15032 47378 15048
rect 47251 14968 47298 15032
rect 47362 14968 47378 15032
rect 47251 14952 47378 14968
rect 47251 14888 47298 14952
rect 47362 14888 47378 14952
rect 47251 14872 47378 14888
rect 47251 14808 47298 14872
rect 47362 14808 47378 14872
rect 47251 14792 47378 14808
rect 47251 14728 47298 14792
rect 47362 14728 47378 14792
rect 47251 14712 47378 14728
rect 47251 14648 47298 14712
rect 47362 14648 47378 14712
rect 47251 14632 47378 14648
rect 47251 14568 47298 14632
rect 47362 14568 47378 14632
rect 47251 14552 47378 14568
rect 47251 14488 47298 14552
rect 47362 14488 47378 14552
rect 47251 14472 47378 14488
rect 47251 14408 47298 14472
rect 47362 14408 47378 14472
rect 47251 14392 47378 14408
rect 47251 14328 47298 14392
rect 47362 14328 47378 14392
rect 47251 14312 47378 14328
rect 47251 14248 47298 14312
rect 47362 14248 47378 14312
rect 47251 14232 47378 14248
rect 47251 14168 47298 14232
rect 47362 14168 47378 14232
rect 47251 14152 47378 14168
rect 47251 14088 47298 14152
rect 47362 14088 47378 14152
rect 47251 14072 47378 14088
rect 47251 14008 47298 14072
rect 47362 14008 47378 14072
rect 47251 13992 47378 14008
rect 47251 13928 47298 13992
rect 47362 13928 47378 13992
rect 47251 13912 47378 13928
rect 47251 13848 47298 13912
rect 47362 13848 47378 13912
rect 47251 13832 47378 13848
rect 47251 13768 47298 13832
rect 47362 13768 47378 13832
rect 47251 13752 47378 13768
rect 47251 13688 47298 13752
rect 47362 13688 47378 13752
rect 47251 13672 47378 13688
rect 47251 13608 47298 13672
rect 47362 13608 47378 13672
rect 47251 13592 47378 13608
rect 47251 13528 47298 13592
rect 47362 13528 47378 13592
rect 47251 13512 47378 13528
rect 47251 13448 47298 13512
rect 47362 13448 47378 13512
rect 47251 13432 47378 13448
rect 47251 13368 47298 13432
rect 47362 13368 47378 13432
rect 47251 13352 47378 13368
rect 47251 13288 47298 13352
rect 47362 13288 47378 13352
rect 47251 13272 47378 13288
rect 47251 13208 47298 13272
rect 47362 13208 47378 13272
rect 47251 13192 47378 13208
rect 47251 13128 47298 13192
rect 47362 13128 47378 13192
rect 47251 13112 47378 13128
rect 47251 13048 47298 13112
rect 47362 13048 47378 13112
rect 47251 13032 47378 13048
rect 47251 12968 47298 13032
rect 47362 12968 47378 13032
rect 47251 12952 47378 12968
rect 47251 12888 47298 12952
rect 47362 12888 47378 12952
rect 47251 12872 47378 12888
rect 47251 12808 47298 12872
rect 47362 12808 47378 12872
rect 47251 12792 47378 12808
rect 47251 12728 47298 12792
rect 47362 12728 47378 12792
rect 47251 12712 47378 12728
rect 47251 12648 47298 12712
rect 47362 12648 47378 12712
rect 47251 12632 47378 12648
rect 47251 12568 47298 12632
rect 47362 12568 47378 12632
rect 47251 12552 47378 12568
rect 47251 12488 47298 12552
rect 47362 12488 47378 12552
rect 47251 12472 47378 12488
rect 47251 12408 47298 12472
rect 47362 12408 47378 12472
rect 47251 12392 47378 12408
rect 47251 12328 47298 12392
rect 47362 12328 47378 12392
rect 47251 12312 47378 12328
rect 47251 12248 47298 12312
rect 47362 12248 47378 12312
rect 47251 12232 47378 12248
rect 47251 12168 47298 12232
rect 47362 12168 47378 12232
rect 47251 12152 47378 12168
rect 47251 12088 47298 12152
rect 47362 12088 47378 12152
rect 47251 12072 47378 12088
rect 47251 12008 47298 12072
rect 47362 12008 47378 12072
rect 47251 11992 47378 12008
rect 47251 11928 47298 11992
rect 47362 11928 47378 11992
rect 47251 11912 47378 11928
rect 47251 11848 47298 11912
rect 47362 11848 47378 11912
rect 47251 11832 47378 11848
rect 47251 11768 47298 11832
rect 47362 11768 47378 11832
rect 47251 11752 47378 11768
rect 47251 11688 47298 11752
rect 47362 11688 47378 11752
rect 47251 11672 47378 11688
rect 47251 11608 47298 11672
rect 47362 11608 47378 11672
rect 47251 11592 47378 11608
rect 47251 11528 47298 11592
rect 47362 11528 47378 11592
rect 47251 11512 47378 11528
rect 47251 11448 47298 11512
rect 47362 11448 47378 11512
rect 47251 11432 47378 11448
rect 47251 11368 47298 11432
rect 47362 11368 47378 11432
rect 47251 11352 47378 11368
rect 47251 11288 47298 11352
rect 47362 11288 47378 11352
rect 47251 11272 47378 11288
rect 47251 11208 47298 11272
rect 47362 11208 47378 11272
rect 47251 11192 47378 11208
rect 47251 11128 47298 11192
rect 47362 11128 47378 11192
rect 47251 11112 47378 11128
rect 47251 11048 47298 11112
rect 47362 11048 47378 11112
rect 47251 11032 47378 11048
rect 47251 10968 47298 11032
rect 47362 10968 47378 11032
rect 47251 10952 47378 10968
rect 47251 10888 47298 10952
rect 47362 10888 47378 10952
rect 47251 10872 47378 10888
rect 47251 10808 47298 10872
rect 47362 10808 47378 10872
rect 47251 10792 47378 10808
rect 47251 10728 47298 10792
rect 47362 10728 47378 10792
rect 47251 10712 47378 10728
rect 47251 10648 47298 10712
rect 47362 10648 47378 10712
rect 47251 10632 47378 10648
rect 47251 10568 47298 10632
rect 47362 10568 47378 10632
rect 47251 10552 47378 10568
rect 47251 10488 47298 10552
rect 47362 10488 47378 10552
rect 47251 10472 47378 10488
rect 47251 10408 47298 10472
rect 47362 10408 47378 10472
rect 47251 10392 47378 10408
rect 47251 10328 47298 10392
rect 47362 10328 47378 10392
rect 47251 10312 47378 10328
rect 47251 10248 47298 10312
rect 47362 10248 47378 10312
rect 47251 10232 47378 10248
rect 47251 10168 47298 10232
rect 47362 10168 47378 10232
rect 47251 10152 47378 10168
rect 47251 10088 47298 10152
rect 47362 10088 47378 10152
rect 47251 10072 47378 10088
rect 47251 10008 47298 10072
rect 47362 10008 47378 10072
rect 47251 9992 47378 10008
rect 47251 9928 47298 9992
rect 47362 9928 47378 9992
rect 47251 9912 47378 9928
rect 47251 9848 47298 9912
rect 47362 9848 47378 9912
rect 47251 9832 47378 9848
rect 47251 9768 47298 9832
rect 47362 9768 47378 9832
rect 47251 9752 47378 9768
rect 47251 9688 47298 9752
rect 47362 9688 47378 9752
rect 47251 9672 47378 9688
rect 40932 9592 41059 9608
rect 40932 9528 40979 9592
rect 41043 9528 41059 9592
rect 40932 9512 41059 9528
rect 40932 9388 41036 9512
rect 40932 9372 41059 9388
rect 40932 9308 40979 9372
rect 41043 9308 41059 9372
rect 40932 9292 41059 9308
rect 34613 9212 34740 9228
rect 34613 9148 34660 9212
rect 34724 9148 34740 9212
rect 34613 9132 34740 9148
rect 34613 9068 34660 9132
rect 34724 9068 34740 9132
rect 34613 9052 34740 9068
rect 34613 8988 34660 9052
rect 34724 8988 34740 9052
rect 34613 8972 34740 8988
rect 34613 8908 34660 8972
rect 34724 8908 34740 8972
rect 34613 8892 34740 8908
rect 34613 8828 34660 8892
rect 34724 8828 34740 8892
rect 34613 8812 34740 8828
rect 34613 8748 34660 8812
rect 34724 8748 34740 8812
rect 34613 8732 34740 8748
rect 34613 8668 34660 8732
rect 34724 8668 34740 8732
rect 34613 8652 34740 8668
rect 34613 8588 34660 8652
rect 34724 8588 34740 8652
rect 34613 8572 34740 8588
rect 34613 8508 34660 8572
rect 34724 8508 34740 8572
rect 34613 8492 34740 8508
rect 34613 8428 34660 8492
rect 34724 8428 34740 8492
rect 34613 8412 34740 8428
rect 34613 8348 34660 8412
rect 34724 8348 34740 8412
rect 34613 8332 34740 8348
rect 34613 8268 34660 8332
rect 34724 8268 34740 8332
rect 34613 8252 34740 8268
rect 34613 8188 34660 8252
rect 34724 8188 34740 8252
rect 34613 8172 34740 8188
rect 34613 8108 34660 8172
rect 34724 8108 34740 8172
rect 34613 8092 34740 8108
rect 34613 8028 34660 8092
rect 34724 8028 34740 8092
rect 34613 8012 34740 8028
rect 34613 7948 34660 8012
rect 34724 7948 34740 8012
rect 34613 7932 34740 7948
rect 34613 7868 34660 7932
rect 34724 7868 34740 7932
rect 34613 7852 34740 7868
rect 34613 7788 34660 7852
rect 34724 7788 34740 7852
rect 34613 7772 34740 7788
rect 34613 7708 34660 7772
rect 34724 7708 34740 7772
rect 34613 7692 34740 7708
rect 34613 7628 34660 7692
rect 34724 7628 34740 7692
rect 34613 7612 34740 7628
rect 34613 7548 34660 7612
rect 34724 7548 34740 7612
rect 34613 7532 34740 7548
rect 34613 7468 34660 7532
rect 34724 7468 34740 7532
rect 34613 7452 34740 7468
rect 34613 7388 34660 7452
rect 34724 7388 34740 7452
rect 34613 7372 34740 7388
rect 34613 7308 34660 7372
rect 34724 7308 34740 7372
rect 34613 7292 34740 7308
rect 34613 7228 34660 7292
rect 34724 7228 34740 7292
rect 34613 7212 34740 7228
rect 34613 7148 34660 7212
rect 34724 7148 34740 7212
rect 34613 7132 34740 7148
rect 34613 7068 34660 7132
rect 34724 7068 34740 7132
rect 34613 7052 34740 7068
rect 34613 6988 34660 7052
rect 34724 6988 34740 7052
rect 34613 6972 34740 6988
rect 34613 6908 34660 6972
rect 34724 6908 34740 6972
rect 34613 6892 34740 6908
rect 34613 6828 34660 6892
rect 34724 6828 34740 6892
rect 34613 6812 34740 6828
rect 34613 6748 34660 6812
rect 34724 6748 34740 6812
rect 34613 6732 34740 6748
rect 34613 6668 34660 6732
rect 34724 6668 34740 6732
rect 34613 6652 34740 6668
rect 34613 6588 34660 6652
rect 34724 6588 34740 6652
rect 34613 6572 34740 6588
rect 34613 6508 34660 6572
rect 34724 6508 34740 6572
rect 34613 6492 34740 6508
rect 34613 6428 34660 6492
rect 34724 6428 34740 6492
rect 34613 6412 34740 6428
rect 34613 6348 34660 6412
rect 34724 6348 34740 6412
rect 34613 6332 34740 6348
rect 34613 6268 34660 6332
rect 34724 6268 34740 6332
rect 34613 6252 34740 6268
rect 34613 6188 34660 6252
rect 34724 6188 34740 6252
rect 34613 6172 34740 6188
rect 34613 6108 34660 6172
rect 34724 6108 34740 6172
rect 34613 6092 34740 6108
rect 34613 6028 34660 6092
rect 34724 6028 34740 6092
rect 34613 6012 34740 6028
rect 34613 5948 34660 6012
rect 34724 5948 34740 6012
rect 34613 5932 34740 5948
rect 34613 5868 34660 5932
rect 34724 5868 34740 5932
rect 34613 5852 34740 5868
rect 34613 5788 34660 5852
rect 34724 5788 34740 5852
rect 34613 5772 34740 5788
rect 34613 5708 34660 5772
rect 34724 5708 34740 5772
rect 34613 5692 34740 5708
rect 34613 5628 34660 5692
rect 34724 5628 34740 5692
rect 34613 5612 34740 5628
rect 34613 5548 34660 5612
rect 34724 5548 34740 5612
rect 34613 5532 34740 5548
rect 34613 5468 34660 5532
rect 34724 5468 34740 5532
rect 34613 5452 34740 5468
rect 34613 5388 34660 5452
rect 34724 5388 34740 5452
rect 34613 5372 34740 5388
rect 34613 5308 34660 5372
rect 34724 5308 34740 5372
rect 34613 5292 34740 5308
rect 34613 5228 34660 5292
rect 34724 5228 34740 5292
rect 34613 5212 34740 5228
rect 34613 5148 34660 5212
rect 34724 5148 34740 5212
rect 34613 5132 34740 5148
rect 34613 5068 34660 5132
rect 34724 5068 34740 5132
rect 34613 5052 34740 5068
rect 34613 4988 34660 5052
rect 34724 4988 34740 5052
rect 34613 4972 34740 4988
rect 34613 4908 34660 4972
rect 34724 4908 34740 4972
rect 34613 4892 34740 4908
rect 34613 4828 34660 4892
rect 34724 4828 34740 4892
rect 34613 4812 34740 4828
rect 34613 4748 34660 4812
rect 34724 4748 34740 4812
rect 34613 4732 34740 4748
rect 34613 4668 34660 4732
rect 34724 4668 34740 4732
rect 34613 4652 34740 4668
rect 34613 4588 34660 4652
rect 34724 4588 34740 4652
rect 34613 4572 34740 4588
rect 34613 4508 34660 4572
rect 34724 4508 34740 4572
rect 34613 4492 34740 4508
rect 34613 4428 34660 4492
rect 34724 4428 34740 4492
rect 34613 4412 34740 4428
rect 34613 4348 34660 4412
rect 34724 4348 34740 4412
rect 34613 4332 34740 4348
rect 34613 4268 34660 4332
rect 34724 4268 34740 4332
rect 34613 4252 34740 4268
rect 34613 4188 34660 4252
rect 34724 4188 34740 4252
rect 34613 4172 34740 4188
rect 34613 4108 34660 4172
rect 34724 4108 34740 4172
rect 34613 4092 34740 4108
rect 34613 4028 34660 4092
rect 34724 4028 34740 4092
rect 34613 4012 34740 4028
rect 34613 3948 34660 4012
rect 34724 3948 34740 4012
rect 34613 3932 34740 3948
rect 34613 3868 34660 3932
rect 34724 3868 34740 3932
rect 34613 3852 34740 3868
rect 34613 3788 34660 3852
rect 34724 3788 34740 3852
rect 34613 3772 34740 3788
rect 34613 3708 34660 3772
rect 34724 3708 34740 3772
rect 34613 3692 34740 3708
rect 34613 3628 34660 3692
rect 34724 3628 34740 3692
rect 34613 3612 34740 3628
rect 34613 3548 34660 3612
rect 34724 3548 34740 3612
rect 34613 3532 34740 3548
rect 34613 3468 34660 3532
rect 34724 3468 34740 3532
rect 34613 3452 34740 3468
rect 34613 3388 34660 3452
rect 34724 3388 34740 3452
rect 34613 3372 34740 3388
rect 28294 3292 28421 3308
rect 28294 3228 28341 3292
rect 28405 3228 28421 3292
rect 28294 3212 28421 3228
rect 28294 3088 28398 3212
rect 28294 3072 28421 3088
rect 28294 3008 28341 3072
rect 28405 3008 28421 3072
rect 28294 2992 28421 3008
rect 21975 2912 22102 2928
rect 21975 2848 22022 2912
rect 22086 2848 22102 2912
rect 21975 2832 22102 2848
rect 21975 2768 22022 2832
rect 22086 2768 22102 2832
rect 21975 2752 22102 2768
rect 21975 2688 22022 2752
rect 22086 2688 22102 2752
rect 21975 2672 22102 2688
rect 21975 2608 22022 2672
rect 22086 2608 22102 2672
rect 21975 2592 22102 2608
rect 21975 2528 22022 2592
rect 22086 2528 22102 2592
rect 21975 2512 22102 2528
rect 21975 2448 22022 2512
rect 22086 2448 22102 2512
rect 21975 2432 22102 2448
rect 21975 2368 22022 2432
rect 22086 2368 22102 2432
rect 21975 2352 22102 2368
rect 21975 2288 22022 2352
rect 22086 2288 22102 2352
rect 21975 2272 22102 2288
rect 21975 2208 22022 2272
rect 22086 2208 22102 2272
rect 21975 2192 22102 2208
rect 21975 2128 22022 2192
rect 22086 2128 22102 2192
rect 21975 2112 22102 2128
rect 21975 2048 22022 2112
rect 22086 2048 22102 2112
rect 21975 2032 22102 2048
rect 21975 1968 22022 2032
rect 22086 1968 22102 2032
rect 21975 1952 22102 1968
rect 21975 1888 22022 1952
rect 22086 1888 22102 1952
rect 21975 1872 22102 1888
rect 21975 1808 22022 1872
rect 22086 1808 22102 1872
rect 21975 1792 22102 1808
rect 21975 1728 22022 1792
rect 22086 1728 22102 1792
rect 21975 1712 22102 1728
rect 21975 1648 22022 1712
rect 22086 1648 22102 1712
rect 21975 1632 22102 1648
rect 21975 1568 22022 1632
rect 22086 1568 22102 1632
rect 21975 1552 22102 1568
rect 21975 1488 22022 1552
rect 22086 1488 22102 1552
rect 21975 1472 22102 1488
rect 21975 1408 22022 1472
rect 22086 1408 22102 1472
rect 21975 1392 22102 1408
rect 21975 1328 22022 1392
rect 22086 1328 22102 1392
rect 21975 1312 22102 1328
rect 21975 1248 22022 1312
rect 22086 1248 22102 1312
rect 21975 1232 22102 1248
rect 21975 1168 22022 1232
rect 22086 1168 22102 1232
rect 21975 1152 22102 1168
rect 21975 1088 22022 1152
rect 22086 1088 22102 1152
rect 21975 1072 22102 1088
rect 21975 1008 22022 1072
rect 22086 1008 22102 1072
rect 21975 992 22102 1008
rect 21975 928 22022 992
rect 22086 928 22102 992
rect 21975 912 22102 928
rect 21975 848 22022 912
rect 22086 848 22102 912
rect 21975 832 22102 848
rect 21975 768 22022 832
rect 22086 768 22102 832
rect 21975 752 22102 768
rect 21975 688 22022 752
rect 22086 688 22102 752
rect 21975 672 22102 688
rect 21975 608 22022 672
rect 22086 608 22102 672
rect 21975 592 22102 608
rect 21975 528 22022 592
rect 22086 528 22102 592
rect 21975 512 22102 528
rect 21975 448 22022 512
rect 22086 448 22102 512
rect 21975 432 22102 448
rect 21975 368 22022 432
rect 22086 368 22102 432
rect 21975 352 22102 368
rect 21975 288 22022 352
rect 22086 288 22102 352
rect 21975 272 22102 288
rect 21975 208 22022 272
rect 22086 208 22102 272
rect 21975 192 22102 208
rect 21975 128 22022 192
rect 22086 128 22102 192
rect 21975 112 22102 128
rect 21975 48 22022 112
rect 22086 48 22102 112
rect 21975 32 22102 48
rect 21975 -32 22022 32
rect 22086 -32 22102 32
rect 21975 -48 22102 -32
rect 21975 -112 22022 -48
rect 22086 -112 22102 -48
rect 21975 -128 22102 -112
rect 21975 -192 22022 -128
rect 22086 -192 22102 -128
rect 21975 -208 22102 -192
rect 21975 -272 22022 -208
rect 22086 -272 22102 -208
rect 21975 -288 22102 -272
rect 21975 -352 22022 -288
rect 22086 -352 22102 -288
rect 21975 -368 22102 -352
rect 21975 -432 22022 -368
rect 22086 -432 22102 -368
rect 21975 -448 22102 -432
rect 21975 -512 22022 -448
rect 22086 -512 22102 -448
rect 21975 -528 22102 -512
rect 21975 -592 22022 -528
rect 22086 -592 22102 -528
rect 21975 -608 22102 -592
rect 21975 -672 22022 -608
rect 22086 -672 22102 -608
rect 21975 -688 22102 -672
rect 21975 -752 22022 -688
rect 22086 -752 22102 -688
rect 21975 -768 22102 -752
rect 21975 -832 22022 -768
rect 22086 -832 22102 -768
rect 21975 -848 22102 -832
rect 21975 -912 22022 -848
rect 22086 -912 22102 -848
rect 21975 -928 22102 -912
rect 21975 -992 22022 -928
rect 22086 -992 22102 -928
rect 21975 -1008 22102 -992
rect 21975 -1072 22022 -1008
rect 22086 -1072 22102 -1008
rect 21975 -1088 22102 -1072
rect 21975 -1152 22022 -1088
rect 22086 -1152 22102 -1088
rect 21975 -1168 22102 -1152
rect 21975 -1232 22022 -1168
rect 22086 -1232 22102 -1168
rect 21975 -1248 22102 -1232
rect 21975 -1312 22022 -1248
rect 22086 -1312 22102 -1248
rect 21975 -1328 22102 -1312
rect 21975 -1392 22022 -1328
rect 22086 -1392 22102 -1328
rect 21975 -1408 22102 -1392
rect 21975 -1472 22022 -1408
rect 22086 -1472 22102 -1408
rect 21975 -1488 22102 -1472
rect 21975 -1552 22022 -1488
rect 22086 -1552 22102 -1488
rect 21975 -1568 22102 -1552
rect 21975 -1632 22022 -1568
rect 22086 -1632 22102 -1568
rect 21975 -1648 22102 -1632
rect 21975 -1712 22022 -1648
rect 22086 -1712 22102 -1648
rect 21975 -1728 22102 -1712
rect 21975 -1792 22022 -1728
rect 22086 -1792 22102 -1728
rect 21975 -1808 22102 -1792
rect 21975 -1872 22022 -1808
rect 22086 -1872 22102 -1808
rect 21975 -1888 22102 -1872
rect 21975 -1952 22022 -1888
rect 22086 -1952 22102 -1888
rect 21975 -1968 22102 -1952
rect 21975 -2032 22022 -1968
rect 22086 -2032 22102 -1968
rect 21975 -2048 22102 -2032
rect 21975 -2112 22022 -2048
rect 22086 -2112 22102 -2048
rect 21975 -2128 22102 -2112
rect 21975 -2192 22022 -2128
rect 22086 -2192 22102 -2128
rect 21975 -2208 22102 -2192
rect 21975 -2272 22022 -2208
rect 22086 -2272 22102 -2208
rect 21975 -2288 22102 -2272
rect 21975 -2352 22022 -2288
rect 22086 -2352 22102 -2288
rect 21975 -2368 22102 -2352
rect 21975 -2432 22022 -2368
rect 22086 -2432 22102 -2368
rect 21975 -2448 22102 -2432
rect 21975 -2512 22022 -2448
rect 22086 -2512 22102 -2448
rect 21975 -2528 22102 -2512
rect 21975 -2592 22022 -2528
rect 22086 -2592 22102 -2528
rect 21975 -2608 22102 -2592
rect 21975 -2672 22022 -2608
rect 22086 -2672 22102 -2608
rect 21975 -2688 22102 -2672
rect 21975 -2752 22022 -2688
rect 22086 -2752 22102 -2688
rect 21975 -2768 22102 -2752
rect 21975 -2832 22022 -2768
rect 22086 -2832 22102 -2768
rect 21975 -2848 22102 -2832
rect 21975 -2912 22022 -2848
rect 22086 -2912 22102 -2848
rect 21975 -2928 22102 -2912
rect 15656 -3008 15783 -2992
rect 15656 -3072 15703 -3008
rect 15767 -3072 15783 -3008
rect 15656 -3088 15783 -3072
rect 15656 -3212 15760 -3088
rect 15656 -3228 15783 -3212
rect 15656 -3292 15703 -3228
rect 15767 -3292 15783 -3228
rect 15656 -3308 15783 -3292
rect 9337 -3388 9464 -3372
rect 9337 -3452 9384 -3388
rect 9448 -3452 9464 -3388
rect 9337 -3468 9464 -3452
rect 9337 -3532 9384 -3468
rect 9448 -3532 9464 -3468
rect 9337 -3548 9464 -3532
rect 9337 -3612 9384 -3548
rect 9448 -3612 9464 -3548
rect 9337 -3628 9464 -3612
rect 9337 -3692 9384 -3628
rect 9448 -3692 9464 -3628
rect 9337 -3708 9464 -3692
rect 9337 -3772 9384 -3708
rect 9448 -3772 9464 -3708
rect 9337 -3788 9464 -3772
rect 9337 -3852 9384 -3788
rect 9448 -3852 9464 -3788
rect 9337 -3868 9464 -3852
rect 9337 -3932 9384 -3868
rect 9448 -3932 9464 -3868
rect 9337 -3948 9464 -3932
rect 9337 -4012 9384 -3948
rect 9448 -4012 9464 -3948
rect 9337 -4028 9464 -4012
rect 9337 -4092 9384 -4028
rect 9448 -4092 9464 -4028
rect 9337 -4108 9464 -4092
rect 9337 -4172 9384 -4108
rect 9448 -4172 9464 -4108
rect 9337 -4188 9464 -4172
rect 9337 -4252 9384 -4188
rect 9448 -4252 9464 -4188
rect 9337 -4268 9464 -4252
rect 9337 -4332 9384 -4268
rect 9448 -4332 9464 -4268
rect 9337 -4348 9464 -4332
rect 9337 -4412 9384 -4348
rect 9448 -4412 9464 -4348
rect 9337 -4428 9464 -4412
rect 9337 -4492 9384 -4428
rect 9448 -4492 9464 -4428
rect 9337 -4508 9464 -4492
rect 9337 -4572 9384 -4508
rect 9448 -4572 9464 -4508
rect 9337 -4588 9464 -4572
rect 9337 -4652 9384 -4588
rect 9448 -4652 9464 -4588
rect 9337 -4668 9464 -4652
rect 9337 -4732 9384 -4668
rect 9448 -4732 9464 -4668
rect 9337 -4748 9464 -4732
rect 9337 -4812 9384 -4748
rect 9448 -4812 9464 -4748
rect 9337 -4828 9464 -4812
rect 9337 -4892 9384 -4828
rect 9448 -4892 9464 -4828
rect 9337 -4908 9464 -4892
rect 9337 -4972 9384 -4908
rect 9448 -4972 9464 -4908
rect 9337 -4988 9464 -4972
rect 9337 -5052 9384 -4988
rect 9448 -5052 9464 -4988
rect 9337 -5068 9464 -5052
rect 9337 -5132 9384 -5068
rect 9448 -5132 9464 -5068
rect 9337 -5148 9464 -5132
rect 9337 -5212 9384 -5148
rect 9448 -5212 9464 -5148
rect 9337 -5228 9464 -5212
rect 9337 -5292 9384 -5228
rect 9448 -5292 9464 -5228
rect 9337 -5308 9464 -5292
rect 9337 -5372 9384 -5308
rect 9448 -5372 9464 -5308
rect 9337 -5388 9464 -5372
rect 9337 -5452 9384 -5388
rect 9448 -5452 9464 -5388
rect 9337 -5468 9464 -5452
rect 9337 -5532 9384 -5468
rect 9448 -5532 9464 -5468
rect 9337 -5548 9464 -5532
rect 9337 -5612 9384 -5548
rect 9448 -5612 9464 -5548
rect 9337 -5628 9464 -5612
rect 9337 -5692 9384 -5628
rect 9448 -5692 9464 -5628
rect 9337 -5708 9464 -5692
rect 9337 -5772 9384 -5708
rect 9448 -5772 9464 -5708
rect 9337 -5788 9464 -5772
rect 9337 -5852 9384 -5788
rect 9448 -5852 9464 -5788
rect 9337 -5868 9464 -5852
rect 9337 -5932 9384 -5868
rect 9448 -5932 9464 -5868
rect 9337 -5948 9464 -5932
rect 9337 -6012 9384 -5948
rect 9448 -6012 9464 -5948
rect 9337 -6028 9464 -6012
rect 9337 -6092 9384 -6028
rect 9448 -6092 9464 -6028
rect 9337 -6108 9464 -6092
rect 9337 -6172 9384 -6108
rect 9448 -6172 9464 -6108
rect 9337 -6188 9464 -6172
rect 9337 -6252 9384 -6188
rect 9448 -6252 9464 -6188
rect 9337 -6268 9464 -6252
rect 9337 -6332 9384 -6268
rect 9448 -6332 9464 -6268
rect 9337 -6348 9464 -6332
rect 9337 -6412 9384 -6348
rect 9448 -6412 9464 -6348
rect 9337 -6428 9464 -6412
rect 9337 -6492 9384 -6428
rect 9448 -6492 9464 -6428
rect 9337 -6508 9464 -6492
rect 9337 -6572 9384 -6508
rect 9448 -6572 9464 -6508
rect 9337 -6588 9464 -6572
rect 9337 -6652 9384 -6588
rect 9448 -6652 9464 -6588
rect 9337 -6668 9464 -6652
rect 9337 -6732 9384 -6668
rect 9448 -6732 9464 -6668
rect 9337 -6748 9464 -6732
rect 9337 -6812 9384 -6748
rect 9448 -6812 9464 -6748
rect 9337 -6828 9464 -6812
rect 9337 -6892 9384 -6828
rect 9448 -6892 9464 -6828
rect 9337 -6908 9464 -6892
rect 9337 -6972 9384 -6908
rect 9448 -6972 9464 -6908
rect 9337 -6988 9464 -6972
rect 9337 -7052 9384 -6988
rect 9448 -7052 9464 -6988
rect 9337 -7068 9464 -7052
rect 9337 -7132 9384 -7068
rect 9448 -7132 9464 -7068
rect 9337 -7148 9464 -7132
rect 9337 -7212 9384 -7148
rect 9448 -7212 9464 -7148
rect 9337 -7228 9464 -7212
rect 9337 -7292 9384 -7228
rect 9448 -7292 9464 -7228
rect 9337 -7308 9464 -7292
rect 9337 -7372 9384 -7308
rect 9448 -7372 9464 -7308
rect 9337 -7388 9464 -7372
rect 9337 -7452 9384 -7388
rect 9448 -7452 9464 -7388
rect 9337 -7468 9464 -7452
rect 9337 -7532 9384 -7468
rect 9448 -7532 9464 -7468
rect 9337 -7548 9464 -7532
rect 9337 -7612 9384 -7548
rect 9448 -7612 9464 -7548
rect 9337 -7628 9464 -7612
rect 9337 -7692 9384 -7628
rect 9448 -7692 9464 -7628
rect 9337 -7708 9464 -7692
rect 9337 -7772 9384 -7708
rect 9448 -7772 9464 -7708
rect 9337 -7788 9464 -7772
rect 9337 -7852 9384 -7788
rect 9448 -7852 9464 -7788
rect 9337 -7868 9464 -7852
rect 9337 -7932 9384 -7868
rect 9448 -7932 9464 -7868
rect 9337 -7948 9464 -7932
rect 9337 -8012 9384 -7948
rect 9448 -8012 9464 -7948
rect 9337 -8028 9464 -8012
rect 9337 -8092 9384 -8028
rect 9448 -8092 9464 -8028
rect 9337 -8108 9464 -8092
rect 9337 -8172 9384 -8108
rect 9448 -8172 9464 -8108
rect 9337 -8188 9464 -8172
rect 9337 -8252 9384 -8188
rect 9448 -8252 9464 -8188
rect 9337 -8268 9464 -8252
rect 9337 -8332 9384 -8268
rect 9448 -8332 9464 -8268
rect 9337 -8348 9464 -8332
rect 9337 -8412 9384 -8348
rect 9448 -8412 9464 -8348
rect 9337 -8428 9464 -8412
rect 9337 -8492 9384 -8428
rect 9448 -8492 9464 -8428
rect 9337 -8508 9464 -8492
rect 9337 -8572 9384 -8508
rect 9448 -8572 9464 -8508
rect 9337 -8588 9464 -8572
rect 9337 -8652 9384 -8588
rect 9448 -8652 9464 -8588
rect 9337 -8668 9464 -8652
rect 9337 -8732 9384 -8668
rect 9448 -8732 9464 -8668
rect 9337 -8748 9464 -8732
rect 9337 -8812 9384 -8748
rect 9448 -8812 9464 -8748
rect 9337 -8828 9464 -8812
rect 9337 -8892 9384 -8828
rect 9448 -8892 9464 -8828
rect 9337 -8908 9464 -8892
rect 9337 -8972 9384 -8908
rect 9448 -8972 9464 -8908
rect 9337 -8988 9464 -8972
rect 9337 -9052 9384 -8988
rect 9448 -9052 9464 -8988
rect 9337 -9068 9464 -9052
rect 9337 -9132 9384 -9068
rect 9448 -9132 9464 -9068
rect 9337 -9148 9464 -9132
rect 9337 -9212 9384 -9148
rect 9448 -9212 9464 -9148
rect 9337 -9228 9464 -9212
rect 3018 -9308 3145 -9292
rect 3018 -9372 3065 -9308
rect 3129 -9372 3145 -9308
rect 3018 -9388 3145 -9372
rect 3018 -9512 3122 -9388
rect 3018 -9528 3145 -9512
rect 3018 -9592 3065 -9528
rect 3129 -9592 3145 -9528
rect 3018 -9608 3145 -9592
rect -3301 -9688 -3174 -9672
rect -3301 -9752 -3254 -9688
rect -3190 -9752 -3174 -9688
rect -3301 -9768 -3174 -9752
rect -3301 -9832 -3254 -9768
rect -3190 -9832 -3174 -9768
rect -3301 -9848 -3174 -9832
rect -3301 -9912 -3254 -9848
rect -3190 -9912 -3174 -9848
rect -3301 -9928 -3174 -9912
rect -3301 -9992 -3254 -9928
rect -3190 -9992 -3174 -9928
rect -3301 -10008 -3174 -9992
rect -3301 -10072 -3254 -10008
rect -3190 -10072 -3174 -10008
rect -3301 -10088 -3174 -10072
rect -3301 -10152 -3254 -10088
rect -3190 -10152 -3174 -10088
rect -3301 -10168 -3174 -10152
rect -3301 -10232 -3254 -10168
rect -3190 -10232 -3174 -10168
rect -3301 -10248 -3174 -10232
rect -3301 -10312 -3254 -10248
rect -3190 -10312 -3174 -10248
rect -3301 -10328 -3174 -10312
rect -3301 -10392 -3254 -10328
rect -3190 -10392 -3174 -10328
rect -3301 -10408 -3174 -10392
rect -3301 -10472 -3254 -10408
rect -3190 -10472 -3174 -10408
rect -3301 -10488 -3174 -10472
rect -3301 -10552 -3254 -10488
rect -3190 -10552 -3174 -10488
rect -3301 -10568 -3174 -10552
rect -3301 -10632 -3254 -10568
rect -3190 -10632 -3174 -10568
rect -3301 -10648 -3174 -10632
rect -3301 -10712 -3254 -10648
rect -3190 -10712 -3174 -10648
rect -3301 -10728 -3174 -10712
rect -3301 -10792 -3254 -10728
rect -3190 -10792 -3174 -10728
rect -3301 -10808 -3174 -10792
rect -3301 -10872 -3254 -10808
rect -3190 -10872 -3174 -10808
rect -3301 -10888 -3174 -10872
rect -3301 -10952 -3254 -10888
rect -3190 -10952 -3174 -10888
rect -3301 -10968 -3174 -10952
rect -3301 -11032 -3254 -10968
rect -3190 -11032 -3174 -10968
rect -3301 -11048 -3174 -11032
rect -3301 -11112 -3254 -11048
rect -3190 -11112 -3174 -11048
rect -3301 -11128 -3174 -11112
rect -3301 -11192 -3254 -11128
rect -3190 -11192 -3174 -11128
rect -3301 -11208 -3174 -11192
rect -3301 -11272 -3254 -11208
rect -3190 -11272 -3174 -11208
rect -3301 -11288 -3174 -11272
rect -3301 -11352 -3254 -11288
rect -3190 -11352 -3174 -11288
rect -3301 -11368 -3174 -11352
rect -3301 -11432 -3254 -11368
rect -3190 -11432 -3174 -11368
rect -3301 -11448 -3174 -11432
rect -3301 -11512 -3254 -11448
rect -3190 -11512 -3174 -11448
rect -3301 -11528 -3174 -11512
rect -3301 -11592 -3254 -11528
rect -3190 -11592 -3174 -11528
rect -3301 -11608 -3174 -11592
rect -3301 -11672 -3254 -11608
rect -3190 -11672 -3174 -11608
rect -3301 -11688 -3174 -11672
rect -3301 -11752 -3254 -11688
rect -3190 -11752 -3174 -11688
rect -3301 -11768 -3174 -11752
rect -3301 -11832 -3254 -11768
rect -3190 -11832 -3174 -11768
rect -3301 -11848 -3174 -11832
rect -3301 -11912 -3254 -11848
rect -3190 -11912 -3174 -11848
rect -3301 -11928 -3174 -11912
rect -3301 -11992 -3254 -11928
rect -3190 -11992 -3174 -11928
rect -3301 -12008 -3174 -11992
rect -3301 -12072 -3254 -12008
rect -3190 -12072 -3174 -12008
rect -3301 -12088 -3174 -12072
rect -3301 -12152 -3254 -12088
rect -3190 -12152 -3174 -12088
rect -3301 -12168 -3174 -12152
rect -3301 -12232 -3254 -12168
rect -3190 -12232 -3174 -12168
rect -3301 -12248 -3174 -12232
rect -3301 -12312 -3254 -12248
rect -3190 -12312 -3174 -12248
rect -3301 -12328 -3174 -12312
rect -3301 -12392 -3254 -12328
rect -3190 -12392 -3174 -12328
rect -3301 -12408 -3174 -12392
rect -3301 -12472 -3254 -12408
rect -3190 -12472 -3174 -12408
rect -3301 -12488 -3174 -12472
rect -3301 -12552 -3254 -12488
rect -3190 -12552 -3174 -12488
rect -3301 -12568 -3174 -12552
rect -3301 -12632 -3254 -12568
rect -3190 -12632 -3174 -12568
rect -3301 -12648 -3174 -12632
rect -3301 -12712 -3254 -12648
rect -3190 -12712 -3174 -12648
rect -3301 -12728 -3174 -12712
rect -3301 -12792 -3254 -12728
rect -3190 -12792 -3174 -12728
rect -3301 -12808 -3174 -12792
rect -3301 -12872 -3254 -12808
rect -3190 -12872 -3174 -12808
rect -3301 -12888 -3174 -12872
rect -3301 -12952 -3254 -12888
rect -3190 -12952 -3174 -12888
rect -3301 -12968 -3174 -12952
rect -3301 -13032 -3254 -12968
rect -3190 -13032 -3174 -12968
rect -3301 -13048 -3174 -13032
rect -3301 -13112 -3254 -13048
rect -3190 -13112 -3174 -13048
rect -3301 -13128 -3174 -13112
rect -3301 -13192 -3254 -13128
rect -3190 -13192 -3174 -13128
rect -3301 -13208 -3174 -13192
rect -3301 -13272 -3254 -13208
rect -3190 -13272 -3174 -13208
rect -3301 -13288 -3174 -13272
rect -3301 -13352 -3254 -13288
rect -3190 -13352 -3174 -13288
rect -3301 -13368 -3174 -13352
rect -3301 -13432 -3254 -13368
rect -3190 -13432 -3174 -13368
rect -3301 -13448 -3174 -13432
rect -3301 -13512 -3254 -13448
rect -3190 -13512 -3174 -13448
rect -3301 -13528 -3174 -13512
rect -3301 -13592 -3254 -13528
rect -3190 -13592 -3174 -13528
rect -3301 -13608 -3174 -13592
rect -3301 -13672 -3254 -13608
rect -3190 -13672 -3174 -13608
rect -3301 -13688 -3174 -13672
rect -3301 -13752 -3254 -13688
rect -3190 -13752 -3174 -13688
rect -3301 -13768 -3174 -13752
rect -3301 -13832 -3254 -13768
rect -3190 -13832 -3174 -13768
rect -3301 -13848 -3174 -13832
rect -3301 -13912 -3254 -13848
rect -3190 -13912 -3174 -13848
rect -3301 -13928 -3174 -13912
rect -3301 -13992 -3254 -13928
rect -3190 -13992 -3174 -13928
rect -3301 -14008 -3174 -13992
rect -3301 -14072 -3254 -14008
rect -3190 -14072 -3174 -14008
rect -3301 -14088 -3174 -14072
rect -3301 -14152 -3254 -14088
rect -3190 -14152 -3174 -14088
rect -3301 -14168 -3174 -14152
rect -3301 -14232 -3254 -14168
rect -3190 -14232 -3174 -14168
rect -3301 -14248 -3174 -14232
rect -3301 -14312 -3254 -14248
rect -3190 -14312 -3174 -14248
rect -3301 -14328 -3174 -14312
rect -3301 -14392 -3254 -14328
rect -3190 -14392 -3174 -14328
rect -3301 -14408 -3174 -14392
rect -3301 -14472 -3254 -14408
rect -3190 -14472 -3174 -14408
rect -3301 -14488 -3174 -14472
rect -3301 -14552 -3254 -14488
rect -3190 -14552 -3174 -14488
rect -3301 -14568 -3174 -14552
rect -3301 -14632 -3254 -14568
rect -3190 -14632 -3174 -14568
rect -3301 -14648 -3174 -14632
rect -3301 -14712 -3254 -14648
rect -3190 -14712 -3174 -14648
rect -3301 -14728 -3174 -14712
rect -3301 -14792 -3254 -14728
rect -3190 -14792 -3174 -14728
rect -3301 -14808 -3174 -14792
rect -3301 -14872 -3254 -14808
rect -3190 -14872 -3174 -14808
rect -3301 -14888 -3174 -14872
rect -3301 -14952 -3254 -14888
rect -3190 -14952 -3174 -14888
rect -3301 -14968 -3174 -14952
rect -3301 -15032 -3254 -14968
rect -3190 -15032 -3174 -14968
rect -3301 -15048 -3174 -15032
rect -3301 -15112 -3254 -15048
rect -3190 -15112 -3174 -15048
rect -3301 -15128 -3174 -15112
rect -3301 -15192 -3254 -15128
rect -3190 -15192 -3174 -15128
rect -3301 -15208 -3174 -15192
rect -3301 -15272 -3254 -15208
rect -3190 -15272 -3174 -15208
rect -3301 -15288 -3174 -15272
rect -3301 -15352 -3254 -15288
rect -3190 -15352 -3174 -15288
rect -3301 -15368 -3174 -15352
rect -3301 -15432 -3254 -15368
rect -3190 -15432 -3174 -15368
rect -3301 -15448 -3174 -15432
rect -3301 -15512 -3254 -15448
rect -3190 -15512 -3174 -15448
rect -3301 -15528 -3174 -15512
rect -9620 -15608 -9493 -15592
rect -9620 -15672 -9573 -15608
rect -9509 -15672 -9493 -15608
rect -9620 -15688 -9493 -15672
rect -9620 -15812 -9516 -15688
rect -9620 -15828 -9493 -15812
rect -9620 -15892 -9573 -15828
rect -9509 -15892 -9493 -15828
rect -9620 -15908 -9493 -15892
rect -15939 -15988 -15812 -15972
rect -15939 -16052 -15892 -15988
rect -15828 -16052 -15812 -15988
rect -15939 -16068 -15812 -16052
rect -15939 -16132 -15892 -16068
rect -15828 -16132 -15812 -16068
rect -15939 -16148 -15812 -16132
rect -15939 -16212 -15892 -16148
rect -15828 -16212 -15812 -16148
rect -15939 -16228 -15812 -16212
rect -15939 -16292 -15892 -16228
rect -15828 -16292 -15812 -16228
rect -15939 -16308 -15812 -16292
rect -15939 -16372 -15892 -16308
rect -15828 -16372 -15812 -16308
rect -15939 -16388 -15812 -16372
rect -15939 -16452 -15892 -16388
rect -15828 -16452 -15812 -16388
rect -15939 -16468 -15812 -16452
rect -15939 -16532 -15892 -16468
rect -15828 -16532 -15812 -16468
rect -15939 -16548 -15812 -16532
rect -15939 -16612 -15892 -16548
rect -15828 -16612 -15812 -16548
rect -15939 -16628 -15812 -16612
rect -15939 -16692 -15892 -16628
rect -15828 -16692 -15812 -16628
rect -15939 -16708 -15812 -16692
rect -15939 -16772 -15892 -16708
rect -15828 -16772 -15812 -16708
rect -15939 -16788 -15812 -16772
rect -15939 -16852 -15892 -16788
rect -15828 -16852 -15812 -16788
rect -15939 -16868 -15812 -16852
rect -15939 -16932 -15892 -16868
rect -15828 -16932 -15812 -16868
rect -15939 -16948 -15812 -16932
rect -15939 -17012 -15892 -16948
rect -15828 -17012 -15812 -16948
rect -15939 -17028 -15812 -17012
rect -15939 -17092 -15892 -17028
rect -15828 -17092 -15812 -17028
rect -15939 -17108 -15812 -17092
rect -15939 -17172 -15892 -17108
rect -15828 -17172 -15812 -17108
rect -15939 -17188 -15812 -17172
rect -15939 -17252 -15892 -17188
rect -15828 -17252 -15812 -17188
rect -15939 -17268 -15812 -17252
rect -15939 -17332 -15892 -17268
rect -15828 -17332 -15812 -17268
rect -15939 -17348 -15812 -17332
rect -15939 -17412 -15892 -17348
rect -15828 -17412 -15812 -17348
rect -15939 -17428 -15812 -17412
rect -15939 -17492 -15892 -17428
rect -15828 -17492 -15812 -17428
rect -15939 -17508 -15812 -17492
rect -15939 -17572 -15892 -17508
rect -15828 -17572 -15812 -17508
rect -15939 -17588 -15812 -17572
rect -15939 -17652 -15892 -17588
rect -15828 -17652 -15812 -17588
rect -15939 -17668 -15812 -17652
rect -15939 -17732 -15892 -17668
rect -15828 -17732 -15812 -17668
rect -15939 -17748 -15812 -17732
rect -15939 -17812 -15892 -17748
rect -15828 -17812 -15812 -17748
rect -15939 -17828 -15812 -17812
rect -15939 -17892 -15892 -17828
rect -15828 -17892 -15812 -17828
rect -15939 -17908 -15812 -17892
rect -15939 -17972 -15892 -17908
rect -15828 -17972 -15812 -17908
rect -15939 -17988 -15812 -17972
rect -15939 -18052 -15892 -17988
rect -15828 -18052 -15812 -17988
rect -15939 -18068 -15812 -18052
rect -15939 -18132 -15892 -18068
rect -15828 -18132 -15812 -18068
rect -15939 -18148 -15812 -18132
rect -15939 -18212 -15892 -18148
rect -15828 -18212 -15812 -18148
rect -15939 -18228 -15812 -18212
rect -15939 -18292 -15892 -18228
rect -15828 -18292 -15812 -18228
rect -15939 -18308 -15812 -18292
rect -15939 -18372 -15892 -18308
rect -15828 -18372 -15812 -18308
rect -15939 -18388 -15812 -18372
rect -15939 -18452 -15892 -18388
rect -15828 -18452 -15812 -18388
rect -15939 -18468 -15812 -18452
rect -15939 -18532 -15892 -18468
rect -15828 -18532 -15812 -18468
rect -15939 -18548 -15812 -18532
rect -15939 -18612 -15892 -18548
rect -15828 -18612 -15812 -18548
rect -15939 -18628 -15812 -18612
rect -15939 -18692 -15892 -18628
rect -15828 -18692 -15812 -18628
rect -15939 -18708 -15812 -18692
rect -15939 -18772 -15892 -18708
rect -15828 -18772 -15812 -18708
rect -15939 -18788 -15812 -18772
rect -15939 -18852 -15892 -18788
rect -15828 -18852 -15812 -18788
rect -15939 -18868 -15812 -18852
rect -15939 -18932 -15892 -18868
rect -15828 -18932 -15812 -18868
rect -15939 -18948 -15812 -18932
rect -15939 -19012 -15892 -18948
rect -15828 -19012 -15812 -18948
rect -15939 -19028 -15812 -19012
rect -15939 -19092 -15892 -19028
rect -15828 -19092 -15812 -19028
rect -15939 -19108 -15812 -19092
rect -15939 -19172 -15892 -19108
rect -15828 -19172 -15812 -19108
rect -15939 -19188 -15812 -19172
rect -15939 -19252 -15892 -19188
rect -15828 -19252 -15812 -19188
rect -15939 -19268 -15812 -19252
rect -15939 -19332 -15892 -19268
rect -15828 -19332 -15812 -19268
rect -15939 -19348 -15812 -19332
rect -15939 -19412 -15892 -19348
rect -15828 -19412 -15812 -19348
rect -15939 -19428 -15812 -19412
rect -15939 -19492 -15892 -19428
rect -15828 -19492 -15812 -19428
rect -15939 -19508 -15812 -19492
rect -15939 -19572 -15892 -19508
rect -15828 -19572 -15812 -19508
rect -15939 -19588 -15812 -19572
rect -15939 -19652 -15892 -19588
rect -15828 -19652 -15812 -19588
rect -15939 -19668 -15812 -19652
rect -15939 -19732 -15892 -19668
rect -15828 -19732 -15812 -19668
rect -15939 -19748 -15812 -19732
rect -15939 -19812 -15892 -19748
rect -15828 -19812 -15812 -19748
rect -15939 -19828 -15812 -19812
rect -15939 -19892 -15892 -19828
rect -15828 -19892 -15812 -19828
rect -15939 -19908 -15812 -19892
rect -15939 -19972 -15892 -19908
rect -15828 -19972 -15812 -19908
rect -15939 -19988 -15812 -19972
rect -15939 -20052 -15892 -19988
rect -15828 -20052 -15812 -19988
rect -15939 -20068 -15812 -20052
rect -15939 -20132 -15892 -20068
rect -15828 -20132 -15812 -20068
rect -15939 -20148 -15812 -20132
rect -15939 -20212 -15892 -20148
rect -15828 -20212 -15812 -20148
rect -15939 -20228 -15812 -20212
rect -15939 -20292 -15892 -20228
rect -15828 -20292 -15812 -20228
rect -15939 -20308 -15812 -20292
rect -15939 -20372 -15892 -20308
rect -15828 -20372 -15812 -20308
rect -15939 -20388 -15812 -20372
rect -15939 -20452 -15892 -20388
rect -15828 -20452 -15812 -20388
rect -15939 -20468 -15812 -20452
rect -15939 -20532 -15892 -20468
rect -15828 -20532 -15812 -20468
rect -15939 -20548 -15812 -20532
rect -15939 -20612 -15892 -20548
rect -15828 -20612 -15812 -20548
rect -15939 -20628 -15812 -20612
rect -15939 -20692 -15892 -20628
rect -15828 -20692 -15812 -20628
rect -15939 -20708 -15812 -20692
rect -15939 -20772 -15892 -20708
rect -15828 -20772 -15812 -20708
rect -15939 -20788 -15812 -20772
rect -15939 -20852 -15892 -20788
rect -15828 -20852 -15812 -20788
rect -15939 -20868 -15812 -20852
rect -15939 -20932 -15892 -20868
rect -15828 -20932 -15812 -20868
rect -15939 -20948 -15812 -20932
rect -15939 -21012 -15892 -20948
rect -15828 -21012 -15812 -20948
rect -15939 -21028 -15812 -21012
rect -15939 -21092 -15892 -21028
rect -15828 -21092 -15812 -21028
rect -15939 -21108 -15812 -21092
rect -15939 -21172 -15892 -21108
rect -15828 -21172 -15812 -21108
rect -15939 -21188 -15812 -21172
rect -15939 -21252 -15892 -21188
rect -15828 -21252 -15812 -21188
rect -15939 -21268 -15812 -21252
rect -15939 -21332 -15892 -21268
rect -15828 -21332 -15812 -21268
rect -15939 -21348 -15812 -21332
rect -15939 -21412 -15892 -21348
rect -15828 -21412 -15812 -21348
rect -15939 -21428 -15812 -21412
rect -15939 -21492 -15892 -21428
rect -15828 -21492 -15812 -21428
rect -15939 -21508 -15812 -21492
rect -15939 -21572 -15892 -21508
rect -15828 -21572 -15812 -21508
rect -15939 -21588 -15812 -21572
rect -15939 -21652 -15892 -21588
rect -15828 -21652 -15812 -21588
rect -15939 -21668 -15812 -21652
rect -15939 -21732 -15892 -21668
rect -15828 -21732 -15812 -21668
rect -15939 -21748 -15812 -21732
rect -15939 -21812 -15892 -21748
rect -15828 -21812 -15812 -21748
rect -15939 -21828 -15812 -21812
rect -22258 -21908 -22131 -21892
rect -22258 -21972 -22211 -21908
rect -22147 -21972 -22131 -21908
rect -22258 -21988 -22131 -21972
rect -22258 -22112 -22154 -21988
rect -22258 -22128 -22131 -22112
rect -22258 -22192 -22211 -22128
rect -22147 -22192 -22131 -22128
rect -22258 -22208 -22131 -22192
rect -28577 -22288 -28450 -22272
rect -28577 -22352 -28530 -22288
rect -28466 -22352 -28450 -22288
rect -28577 -22368 -28450 -22352
rect -28577 -22432 -28530 -22368
rect -28466 -22432 -28450 -22368
rect -28577 -22448 -28450 -22432
rect -28577 -22512 -28530 -22448
rect -28466 -22512 -28450 -22448
rect -28577 -22528 -28450 -22512
rect -28577 -22592 -28530 -22528
rect -28466 -22592 -28450 -22528
rect -28577 -22608 -28450 -22592
rect -28577 -22672 -28530 -22608
rect -28466 -22672 -28450 -22608
rect -28577 -22688 -28450 -22672
rect -28577 -22752 -28530 -22688
rect -28466 -22752 -28450 -22688
rect -28577 -22768 -28450 -22752
rect -28577 -22832 -28530 -22768
rect -28466 -22832 -28450 -22768
rect -28577 -22848 -28450 -22832
rect -28577 -22912 -28530 -22848
rect -28466 -22912 -28450 -22848
rect -28577 -22928 -28450 -22912
rect -28577 -22992 -28530 -22928
rect -28466 -22992 -28450 -22928
rect -28577 -23008 -28450 -22992
rect -28577 -23072 -28530 -23008
rect -28466 -23072 -28450 -23008
rect -28577 -23088 -28450 -23072
rect -28577 -23152 -28530 -23088
rect -28466 -23152 -28450 -23088
rect -28577 -23168 -28450 -23152
rect -28577 -23232 -28530 -23168
rect -28466 -23232 -28450 -23168
rect -28577 -23248 -28450 -23232
rect -28577 -23312 -28530 -23248
rect -28466 -23312 -28450 -23248
rect -28577 -23328 -28450 -23312
rect -28577 -23392 -28530 -23328
rect -28466 -23392 -28450 -23328
rect -28577 -23408 -28450 -23392
rect -28577 -23472 -28530 -23408
rect -28466 -23472 -28450 -23408
rect -28577 -23488 -28450 -23472
rect -28577 -23552 -28530 -23488
rect -28466 -23552 -28450 -23488
rect -28577 -23568 -28450 -23552
rect -28577 -23632 -28530 -23568
rect -28466 -23632 -28450 -23568
rect -28577 -23648 -28450 -23632
rect -28577 -23712 -28530 -23648
rect -28466 -23712 -28450 -23648
rect -28577 -23728 -28450 -23712
rect -28577 -23792 -28530 -23728
rect -28466 -23792 -28450 -23728
rect -28577 -23808 -28450 -23792
rect -28577 -23872 -28530 -23808
rect -28466 -23872 -28450 -23808
rect -28577 -23888 -28450 -23872
rect -28577 -23952 -28530 -23888
rect -28466 -23952 -28450 -23888
rect -28577 -23968 -28450 -23952
rect -28577 -24032 -28530 -23968
rect -28466 -24032 -28450 -23968
rect -28577 -24048 -28450 -24032
rect -28577 -24112 -28530 -24048
rect -28466 -24112 -28450 -24048
rect -28577 -24128 -28450 -24112
rect -28577 -24192 -28530 -24128
rect -28466 -24192 -28450 -24128
rect -28577 -24208 -28450 -24192
rect -28577 -24272 -28530 -24208
rect -28466 -24272 -28450 -24208
rect -28577 -24288 -28450 -24272
rect -28577 -24352 -28530 -24288
rect -28466 -24352 -28450 -24288
rect -28577 -24368 -28450 -24352
rect -28577 -24432 -28530 -24368
rect -28466 -24432 -28450 -24368
rect -28577 -24448 -28450 -24432
rect -28577 -24512 -28530 -24448
rect -28466 -24512 -28450 -24448
rect -28577 -24528 -28450 -24512
rect -28577 -24592 -28530 -24528
rect -28466 -24592 -28450 -24528
rect -28577 -24608 -28450 -24592
rect -28577 -24672 -28530 -24608
rect -28466 -24672 -28450 -24608
rect -28577 -24688 -28450 -24672
rect -28577 -24752 -28530 -24688
rect -28466 -24752 -28450 -24688
rect -28577 -24768 -28450 -24752
rect -28577 -24832 -28530 -24768
rect -28466 -24832 -28450 -24768
rect -28577 -24848 -28450 -24832
rect -28577 -24912 -28530 -24848
rect -28466 -24912 -28450 -24848
rect -28577 -24928 -28450 -24912
rect -28577 -24992 -28530 -24928
rect -28466 -24992 -28450 -24928
rect -28577 -25008 -28450 -24992
rect -28577 -25072 -28530 -25008
rect -28466 -25072 -28450 -25008
rect -28577 -25088 -28450 -25072
rect -28577 -25152 -28530 -25088
rect -28466 -25152 -28450 -25088
rect -28577 -25168 -28450 -25152
rect -28577 -25232 -28530 -25168
rect -28466 -25232 -28450 -25168
rect -28577 -25248 -28450 -25232
rect -28577 -25312 -28530 -25248
rect -28466 -25312 -28450 -25248
rect -28577 -25328 -28450 -25312
rect -28577 -25392 -28530 -25328
rect -28466 -25392 -28450 -25328
rect -28577 -25408 -28450 -25392
rect -28577 -25472 -28530 -25408
rect -28466 -25472 -28450 -25408
rect -28577 -25488 -28450 -25472
rect -28577 -25552 -28530 -25488
rect -28466 -25552 -28450 -25488
rect -28577 -25568 -28450 -25552
rect -28577 -25632 -28530 -25568
rect -28466 -25632 -28450 -25568
rect -28577 -25648 -28450 -25632
rect -28577 -25712 -28530 -25648
rect -28466 -25712 -28450 -25648
rect -28577 -25728 -28450 -25712
rect -28577 -25792 -28530 -25728
rect -28466 -25792 -28450 -25728
rect -28577 -25808 -28450 -25792
rect -28577 -25872 -28530 -25808
rect -28466 -25872 -28450 -25808
rect -28577 -25888 -28450 -25872
rect -28577 -25952 -28530 -25888
rect -28466 -25952 -28450 -25888
rect -28577 -25968 -28450 -25952
rect -28577 -26032 -28530 -25968
rect -28466 -26032 -28450 -25968
rect -28577 -26048 -28450 -26032
rect -28577 -26112 -28530 -26048
rect -28466 -26112 -28450 -26048
rect -28577 -26128 -28450 -26112
rect -28577 -26192 -28530 -26128
rect -28466 -26192 -28450 -26128
rect -28577 -26208 -28450 -26192
rect -28577 -26272 -28530 -26208
rect -28466 -26272 -28450 -26208
rect -28577 -26288 -28450 -26272
rect -28577 -26352 -28530 -26288
rect -28466 -26352 -28450 -26288
rect -28577 -26368 -28450 -26352
rect -28577 -26432 -28530 -26368
rect -28466 -26432 -28450 -26368
rect -28577 -26448 -28450 -26432
rect -28577 -26512 -28530 -26448
rect -28466 -26512 -28450 -26448
rect -28577 -26528 -28450 -26512
rect -28577 -26592 -28530 -26528
rect -28466 -26592 -28450 -26528
rect -28577 -26608 -28450 -26592
rect -28577 -26672 -28530 -26608
rect -28466 -26672 -28450 -26608
rect -28577 -26688 -28450 -26672
rect -28577 -26752 -28530 -26688
rect -28466 -26752 -28450 -26688
rect -28577 -26768 -28450 -26752
rect -28577 -26832 -28530 -26768
rect -28466 -26832 -28450 -26768
rect -28577 -26848 -28450 -26832
rect -28577 -26912 -28530 -26848
rect -28466 -26912 -28450 -26848
rect -28577 -26928 -28450 -26912
rect -28577 -26992 -28530 -26928
rect -28466 -26992 -28450 -26928
rect -28577 -27008 -28450 -26992
rect -28577 -27072 -28530 -27008
rect -28466 -27072 -28450 -27008
rect -28577 -27088 -28450 -27072
rect -28577 -27152 -28530 -27088
rect -28466 -27152 -28450 -27088
rect -28577 -27168 -28450 -27152
rect -28577 -27232 -28530 -27168
rect -28466 -27232 -28450 -27168
rect -28577 -27248 -28450 -27232
rect -28577 -27312 -28530 -27248
rect -28466 -27312 -28450 -27248
rect -28577 -27328 -28450 -27312
rect -28577 -27392 -28530 -27328
rect -28466 -27392 -28450 -27328
rect -28577 -27408 -28450 -27392
rect -28577 -27472 -28530 -27408
rect -28466 -27472 -28450 -27408
rect -28577 -27488 -28450 -27472
rect -28577 -27552 -28530 -27488
rect -28466 -27552 -28450 -27488
rect -28577 -27568 -28450 -27552
rect -28577 -27632 -28530 -27568
rect -28466 -27632 -28450 -27568
rect -28577 -27648 -28450 -27632
rect -28577 -27712 -28530 -27648
rect -28466 -27712 -28450 -27648
rect -28577 -27728 -28450 -27712
rect -28577 -27792 -28530 -27728
rect -28466 -27792 -28450 -27728
rect -28577 -27808 -28450 -27792
rect -28577 -27872 -28530 -27808
rect -28466 -27872 -28450 -27808
rect -28577 -27888 -28450 -27872
rect -28577 -27952 -28530 -27888
rect -28466 -27952 -28450 -27888
rect -28577 -27968 -28450 -27952
rect -28577 -28032 -28530 -27968
rect -28466 -28032 -28450 -27968
rect -28577 -28048 -28450 -28032
rect -28577 -28112 -28530 -28048
rect -28466 -28112 -28450 -28048
rect -28577 -28128 -28450 -28112
rect -34896 -28208 -34769 -28192
rect -34896 -28272 -34849 -28208
rect -34785 -28272 -34769 -28208
rect -34896 -28288 -34769 -28272
rect -34896 -28412 -34792 -28288
rect -34896 -28428 -34769 -28412
rect -34896 -28492 -34849 -28428
rect -34785 -28492 -34769 -28428
rect -34896 -28508 -34769 -28492
rect -41215 -28588 -41088 -28572
rect -41215 -28652 -41168 -28588
rect -41104 -28652 -41088 -28588
rect -41215 -28668 -41088 -28652
rect -41215 -28732 -41168 -28668
rect -41104 -28732 -41088 -28668
rect -41215 -28748 -41088 -28732
rect -41215 -28812 -41168 -28748
rect -41104 -28812 -41088 -28748
rect -41215 -28828 -41088 -28812
rect -41215 -28892 -41168 -28828
rect -41104 -28892 -41088 -28828
rect -41215 -28908 -41088 -28892
rect -41215 -28972 -41168 -28908
rect -41104 -28972 -41088 -28908
rect -41215 -28988 -41088 -28972
rect -41215 -29052 -41168 -28988
rect -41104 -29052 -41088 -28988
rect -41215 -29068 -41088 -29052
rect -41215 -29132 -41168 -29068
rect -41104 -29132 -41088 -29068
rect -41215 -29148 -41088 -29132
rect -41215 -29212 -41168 -29148
rect -41104 -29212 -41088 -29148
rect -41215 -29228 -41088 -29212
rect -41215 -29292 -41168 -29228
rect -41104 -29292 -41088 -29228
rect -41215 -29308 -41088 -29292
rect -41215 -29372 -41168 -29308
rect -41104 -29372 -41088 -29308
rect -41215 -29388 -41088 -29372
rect -41215 -29452 -41168 -29388
rect -41104 -29452 -41088 -29388
rect -41215 -29468 -41088 -29452
rect -41215 -29532 -41168 -29468
rect -41104 -29532 -41088 -29468
rect -41215 -29548 -41088 -29532
rect -41215 -29612 -41168 -29548
rect -41104 -29612 -41088 -29548
rect -41215 -29628 -41088 -29612
rect -41215 -29692 -41168 -29628
rect -41104 -29692 -41088 -29628
rect -41215 -29708 -41088 -29692
rect -41215 -29772 -41168 -29708
rect -41104 -29772 -41088 -29708
rect -41215 -29788 -41088 -29772
rect -41215 -29852 -41168 -29788
rect -41104 -29852 -41088 -29788
rect -41215 -29868 -41088 -29852
rect -41215 -29932 -41168 -29868
rect -41104 -29932 -41088 -29868
rect -41215 -29948 -41088 -29932
rect -41215 -30012 -41168 -29948
rect -41104 -30012 -41088 -29948
rect -41215 -30028 -41088 -30012
rect -41215 -30092 -41168 -30028
rect -41104 -30092 -41088 -30028
rect -41215 -30108 -41088 -30092
rect -41215 -30172 -41168 -30108
rect -41104 -30172 -41088 -30108
rect -41215 -30188 -41088 -30172
rect -41215 -30252 -41168 -30188
rect -41104 -30252 -41088 -30188
rect -41215 -30268 -41088 -30252
rect -41215 -30332 -41168 -30268
rect -41104 -30332 -41088 -30268
rect -41215 -30348 -41088 -30332
rect -41215 -30412 -41168 -30348
rect -41104 -30412 -41088 -30348
rect -41215 -30428 -41088 -30412
rect -41215 -30492 -41168 -30428
rect -41104 -30492 -41088 -30428
rect -41215 -30508 -41088 -30492
rect -41215 -30572 -41168 -30508
rect -41104 -30572 -41088 -30508
rect -41215 -30588 -41088 -30572
rect -41215 -30652 -41168 -30588
rect -41104 -30652 -41088 -30588
rect -41215 -30668 -41088 -30652
rect -41215 -30732 -41168 -30668
rect -41104 -30732 -41088 -30668
rect -41215 -30748 -41088 -30732
rect -41215 -30812 -41168 -30748
rect -41104 -30812 -41088 -30748
rect -41215 -30828 -41088 -30812
rect -41215 -30892 -41168 -30828
rect -41104 -30892 -41088 -30828
rect -41215 -30908 -41088 -30892
rect -41215 -30972 -41168 -30908
rect -41104 -30972 -41088 -30908
rect -41215 -30988 -41088 -30972
rect -41215 -31052 -41168 -30988
rect -41104 -31052 -41088 -30988
rect -41215 -31068 -41088 -31052
rect -41215 -31132 -41168 -31068
rect -41104 -31132 -41088 -31068
rect -41215 -31148 -41088 -31132
rect -41215 -31212 -41168 -31148
rect -41104 -31212 -41088 -31148
rect -41215 -31228 -41088 -31212
rect -41215 -31292 -41168 -31228
rect -41104 -31292 -41088 -31228
rect -41215 -31308 -41088 -31292
rect -41215 -31372 -41168 -31308
rect -41104 -31372 -41088 -31308
rect -41215 -31388 -41088 -31372
rect -41215 -31452 -41168 -31388
rect -41104 -31452 -41088 -31388
rect -41215 -31468 -41088 -31452
rect -41215 -31532 -41168 -31468
rect -41104 -31532 -41088 -31468
rect -41215 -31548 -41088 -31532
rect -41215 -31612 -41168 -31548
rect -41104 -31612 -41088 -31548
rect -41215 -31628 -41088 -31612
rect -41215 -31692 -41168 -31628
rect -41104 -31692 -41088 -31628
rect -41215 -31708 -41088 -31692
rect -41215 -31772 -41168 -31708
rect -41104 -31772 -41088 -31708
rect -41215 -31788 -41088 -31772
rect -41215 -31852 -41168 -31788
rect -41104 -31852 -41088 -31788
rect -41215 -31868 -41088 -31852
rect -41215 -31932 -41168 -31868
rect -41104 -31932 -41088 -31868
rect -41215 -31948 -41088 -31932
rect -41215 -32012 -41168 -31948
rect -41104 -32012 -41088 -31948
rect -41215 -32028 -41088 -32012
rect -41215 -32092 -41168 -32028
rect -41104 -32092 -41088 -32028
rect -41215 -32108 -41088 -32092
rect -41215 -32172 -41168 -32108
rect -41104 -32172 -41088 -32108
rect -41215 -32188 -41088 -32172
rect -41215 -32252 -41168 -32188
rect -41104 -32252 -41088 -32188
rect -41215 -32268 -41088 -32252
rect -41215 -32332 -41168 -32268
rect -41104 -32332 -41088 -32268
rect -41215 -32348 -41088 -32332
rect -41215 -32412 -41168 -32348
rect -41104 -32412 -41088 -32348
rect -41215 -32428 -41088 -32412
rect -41215 -32492 -41168 -32428
rect -41104 -32492 -41088 -32428
rect -41215 -32508 -41088 -32492
rect -41215 -32572 -41168 -32508
rect -41104 -32572 -41088 -32508
rect -41215 -32588 -41088 -32572
rect -41215 -32652 -41168 -32588
rect -41104 -32652 -41088 -32588
rect -41215 -32668 -41088 -32652
rect -41215 -32732 -41168 -32668
rect -41104 -32732 -41088 -32668
rect -41215 -32748 -41088 -32732
rect -41215 -32812 -41168 -32748
rect -41104 -32812 -41088 -32748
rect -41215 -32828 -41088 -32812
rect -41215 -32892 -41168 -32828
rect -41104 -32892 -41088 -32828
rect -41215 -32908 -41088 -32892
rect -41215 -32972 -41168 -32908
rect -41104 -32972 -41088 -32908
rect -41215 -32988 -41088 -32972
rect -41215 -33052 -41168 -32988
rect -41104 -33052 -41088 -32988
rect -41215 -33068 -41088 -33052
rect -41215 -33132 -41168 -33068
rect -41104 -33132 -41088 -33068
rect -41215 -33148 -41088 -33132
rect -41215 -33212 -41168 -33148
rect -41104 -33212 -41088 -33148
rect -41215 -33228 -41088 -33212
rect -41215 -33292 -41168 -33228
rect -41104 -33292 -41088 -33228
rect -41215 -33308 -41088 -33292
rect -41215 -33372 -41168 -33308
rect -41104 -33372 -41088 -33308
rect -41215 -33388 -41088 -33372
rect -41215 -33452 -41168 -33388
rect -41104 -33452 -41088 -33388
rect -41215 -33468 -41088 -33452
rect -41215 -33532 -41168 -33468
rect -41104 -33532 -41088 -33468
rect -41215 -33548 -41088 -33532
rect -41215 -33612 -41168 -33548
rect -41104 -33612 -41088 -33548
rect -41215 -33628 -41088 -33612
rect -41215 -33692 -41168 -33628
rect -41104 -33692 -41088 -33628
rect -41215 -33708 -41088 -33692
rect -41215 -33772 -41168 -33708
rect -41104 -33772 -41088 -33708
rect -41215 -33788 -41088 -33772
rect -41215 -33852 -41168 -33788
rect -41104 -33852 -41088 -33788
rect -41215 -33868 -41088 -33852
rect -41215 -33932 -41168 -33868
rect -41104 -33932 -41088 -33868
rect -41215 -33948 -41088 -33932
rect -41215 -34012 -41168 -33948
rect -41104 -34012 -41088 -33948
rect -41215 -34028 -41088 -34012
rect -41215 -34092 -41168 -34028
rect -41104 -34092 -41088 -34028
rect -41215 -34108 -41088 -34092
rect -41215 -34172 -41168 -34108
rect -41104 -34172 -41088 -34108
rect -41215 -34188 -41088 -34172
rect -41215 -34252 -41168 -34188
rect -41104 -34252 -41088 -34188
rect -41215 -34268 -41088 -34252
rect -41215 -34332 -41168 -34268
rect -41104 -34332 -41088 -34268
rect -41215 -34348 -41088 -34332
rect -41215 -34412 -41168 -34348
rect -41104 -34412 -41088 -34348
rect -41215 -34428 -41088 -34412
rect -44335 -34839 -44231 -34461
rect -41215 -34492 -41168 -34428
rect -41104 -34492 -41088 -34428
rect -40925 -28548 -35003 -28539
rect -40925 -34452 -40916 -28548
rect -35012 -34452 -35003 -28548
rect -40925 -34461 -35003 -34452
rect -34896 -28572 -34849 -28508
rect -34785 -28572 -34769 -28508
rect -31697 -28539 -31593 -28161
rect -28577 -28192 -28530 -28128
rect -28466 -28192 -28450 -28128
rect -28287 -22248 -22365 -22239
rect -28287 -28152 -28278 -22248
rect -22374 -28152 -22365 -22248
rect -28287 -28161 -22365 -28152
rect -22258 -22272 -22211 -22208
rect -22147 -22272 -22131 -22208
rect -19059 -22239 -18955 -21861
rect -15939 -21892 -15892 -21828
rect -15828 -21892 -15812 -21828
rect -15649 -15948 -9727 -15939
rect -15649 -21852 -15640 -15948
rect -9736 -21852 -9727 -15948
rect -15649 -21861 -9727 -21852
rect -9620 -15972 -9573 -15908
rect -9509 -15972 -9493 -15908
rect -6421 -15939 -6317 -15561
rect -3301 -15592 -3254 -15528
rect -3190 -15592 -3174 -15528
rect -3011 -9648 2911 -9639
rect -3011 -15552 -3002 -9648
rect 2902 -15552 2911 -9648
rect -3011 -15561 2911 -15552
rect 3018 -9672 3065 -9608
rect 3129 -9672 3145 -9608
rect 6217 -9639 6321 -9261
rect 9337 -9292 9384 -9228
rect 9448 -9292 9464 -9228
rect 9627 -3348 15549 -3339
rect 9627 -9252 9636 -3348
rect 15540 -9252 15549 -3348
rect 9627 -9261 15549 -9252
rect 15656 -3372 15703 -3308
rect 15767 -3372 15783 -3308
rect 18855 -3339 18959 -2961
rect 21975 -2992 22022 -2928
rect 22086 -2992 22102 -2928
rect 22265 2952 28187 2961
rect 22265 -2952 22274 2952
rect 28178 -2952 28187 2952
rect 22265 -2961 28187 -2952
rect 28294 2928 28341 2992
rect 28405 2928 28421 2992
rect 31493 2961 31597 3339
rect 34613 3308 34660 3372
rect 34724 3308 34740 3372
rect 34903 9252 40825 9261
rect 34903 3348 34912 9252
rect 40816 3348 40825 9252
rect 34903 3339 40825 3348
rect 40932 9228 40979 9292
rect 41043 9228 41059 9292
rect 44131 9261 44235 9639
rect 47251 9608 47298 9672
rect 47362 9608 47378 9672
rect 47251 9592 47378 9608
rect 47251 9528 47298 9592
rect 47362 9528 47378 9592
rect 47251 9512 47378 9528
rect 47251 9388 47355 9512
rect 47251 9372 47378 9388
rect 47251 9308 47298 9372
rect 47362 9308 47378 9372
rect 47251 9292 47378 9308
rect 40932 9212 41059 9228
rect 40932 9148 40979 9212
rect 41043 9148 41059 9212
rect 40932 9132 41059 9148
rect 40932 9068 40979 9132
rect 41043 9068 41059 9132
rect 40932 9052 41059 9068
rect 40932 8988 40979 9052
rect 41043 8988 41059 9052
rect 40932 8972 41059 8988
rect 40932 8908 40979 8972
rect 41043 8908 41059 8972
rect 40932 8892 41059 8908
rect 40932 8828 40979 8892
rect 41043 8828 41059 8892
rect 40932 8812 41059 8828
rect 40932 8748 40979 8812
rect 41043 8748 41059 8812
rect 40932 8732 41059 8748
rect 40932 8668 40979 8732
rect 41043 8668 41059 8732
rect 40932 8652 41059 8668
rect 40932 8588 40979 8652
rect 41043 8588 41059 8652
rect 40932 8572 41059 8588
rect 40932 8508 40979 8572
rect 41043 8508 41059 8572
rect 40932 8492 41059 8508
rect 40932 8428 40979 8492
rect 41043 8428 41059 8492
rect 40932 8412 41059 8428
rect 40932 8348 40979 8412
rect 41043 8348 41059 8412
rect 40932 8332 41059 8348
rect 40932 8268 40979 8332
rect 41043 8268 41059 8332
rect 40932 8252 41059 8268
rect 40932 8188 40979 8252
rect 41043 8188 41059 8252
rect 40932 8172 41059 8188
rect 40932 8108 40979 8172
rect 41043 8108 41059 8172
rect 40932 8092 41059 8108
rect 40932 8028 40979 8092
rect 41043 8028 41059 8092
rect 40932 8012 41059 8028
rect 40932 7948 40979 8012
rect 41043 7948 41059 8012
rect 40932 7932 41059 7948
rect 40932 7868 40979 7932
rect 41043 7868 41059 7932
rect 40932 7852 41059 7868
rect 40932 7788 40979 7852
rect 41043 7788 41059 7852
rect 40932 7772 41059 7788
rect 40932 7708 40979 7772
rect 41043 7708 41059 7772
rect 40932 7692 41059 7708
rect 40932 7628 40979 7692
rect 41043 7628 41059 7692
rect 40932 7612 41059 7628
rect 40932 7548 40979 7612
rect 41043 7548 41059 7612
rect 40932 7532 41059 7548
rect 40932 7468 40979 7532
rect 41043 7468 41059 7532
rect 40932 7452 41059 7468
rect 40932 7388 40979 7452
rect 41043 7388 41059 7452
rect 40932 7372 41059 7388
rect 40932 7308 40979 7372
rect 41043 7308 41059 7372
rect 40932 7292 41059 7308
rect 40932 7228 40979 7292
rect 41043 7228 41059 7292
rect 40932 7212 41059 7228
rect 40932 7148 40979 7212
rect 41043 7148 41059 7212
rect 40932 7132 41059 7148
rect 40932 7068 40979 7132
rect 41043 7068 41059 7132
rect 40932 7052 41059 7068
rect 40932 6988 40979 7052
rect 41043 6988 41059 7052
rect 40932 6972 41059 6988
rect 40932 6908 40979 6972
rect 41043 6908 41059 6972
rect 40932 6892 41059 6908
rect 40932 6828 40979 6892
rect 41043 6828 41059 6892
rect 40932 6812 41059 6828
rect 40932 6748 40979 6812
rect 41043 6748 41059 6812
rect 40932 6732 41059 6748
rect 40932 6668 40979 6732
rect 41043 6668 41059 6732
rect 40932 6652 41059 6668
rect 40932 6588 40979 6652
rect 41043 6588 41059 6652
rect 40932 6572 41059 6588
rect 40932 6508 40979 6572
rect 41043 6508 41059 6572
rect 40932 6492 41059 6508
rect 40932 6428 40979 6492
rect 41043 6428 41059 6492
rect 40932 6412 41059 6428
rect 40932 6348 40979 6412
rect 41043 6348 41059 6412
rect 40932 6332 41059 6348
rect 40932 6268 40979 6332
rect 41043 6268 41059 6332
rect 40932 6252 41059 6268
rect 40932 6188 40979 6252
rect 41043 6188 41059 6252
rect 40932 6172 41059 6188
rect 40932 6108 40979 6172
rect 41043 6108 41059 6172
rect 40932 6092 41059 6108
rect 40932 6028 40979 6092
rect 41043 6028 41059 6092
rect 40932 6012 41059 6028
rect 40932 5948 40979 6012
rect 41043 5948 41059 6012
rect 40932 5932 41059 5948
rect 40932 5868 40979 5932
rect 41043 5868 41059 5932
rect 40932 5852 41059 5868
rect 40932 5788 40979 5852
rect 41043 5788 41059 5852
rect 40932 5772 41059 5788
rect 40932 5708 40979 5772
rect 41043 5708 41059 5772
rect 40932 5692 41059 5708
rect 40932 5628 40979 5692
rect 41043 5628 41059 5692
rect 40932 5612 41059 5628
rect 40932 5548 40979 5612
rect 41043 5548 41059 5612
rect 40932 5532 41059 5548
rect 40932 5468 40979 5532
rect 41043 5468 41059 5532
rect 40932 5452 41059 5468
rect 40932 5388 40979 5452
rect 41043 5388 41059 5452
rect 40932 5372 41059 5388
rect 40932 5308 40979 5372
rect 41043 5308 41059 5372
rect 40932 5292 41059 5308
rect 40932 5228 40979 5292
rect 41043 5228 41059 5292
rect 40932 5212 41059 5228
rect 40932 5148 40979 5212
rect 41043 5148 41059 5212
rect 40932 5132 41059 5148
rect 40932 5068 40979 5132
rect 41043 5068 41059 5132
rect 40932 5052 41059 5068
rect 40932 4988 40979 5052
rect 41043 4988 41059 5052
rect 40932 4972 41059 4988
rect 40932 4908 40979 4972
rect 41043 4908 41059 4972
rect 40932 4892 41059 4908
rect 40932 4828 40979 4892
rect 41043 4828 41059 4892
rect 40932 4812 41059 4828
rect 40932 4748 40979 4812
rect 41043 4748 41059 4812
rect 40932 4732 41059 4748
rect 40932 4668 40979 4732
rect 41043 4668 41059 4732
rect 40932 4652 41059 4668
rect 40932 4588 40979 4652
rect 41043 4588 41059 4652
rect 40932 4572 41059 4588
rect 40932 4508 40979 4572
rect 41043 4508 41059 4572
rect 40932 4492 41059 4508
rect 40932 4428 40979 4492
rect 41043 4428 41059 4492
rect 40932 4412 41059 4428
rect 40932 4348 40979 4412
rect 41043 4348 41059 4412
rect 40932 4332 41059 4348
rect 40932 4268 40979 4332
rect 41043 4268 41059 4332
rect 40932 4252 41059 4268
rect 40932 4188 40979 4252
rect 41043 4188 41059 4252
rect 40932 4172 41059 4188
rect 40932 4108 40979 4172
rect 41043 4108 41059 4172
rect 40932 4092 41059 4108
rect 40932 4028 40979 4092
rect 41043 4028 41059 4092
rect 40932 4012 41059 4028
rect 40932 3948 40979 4012
rect 41043 3948 41059 4012
rect 40932 3932 41059 3948
rect 40932 3868 40979 3932
rect 41043 3868 41059 3932
rect 40932 3852 41059 3868
rect 40932 3788 40979 3852
rect 41043 3788 41059 3852
rect 40932 3772 41059 3788
rect 40932 3708 40979 3772
rect 41043 3708 41059 3772
rect 40932 3692 41059 3708
rect 40932 3628 40979 3692
rect 41043 3628 41059 3692
rect 40932 3612 41059 3628
rect 40932 3548 40979 3612
rect 41043 3548 41059 3612
rect 40932 3532 41059 3548
rect 40932 3468 40979 3532
rect 41043 3468 41059 3532
rect 40932 3452 41059 3468
rect 40932 3388 40979 3452
rect 41043 3388 41059 3452
rect 40932 3372 41059 3388
rect 34613 3292 34740 3308
rect 34613 3228 34660 3292
rect 34724 3228 34740 3292
rect 34613 3212 34740 3228
rect 34613 3088 34717 3212
rect 34613 3072 34740 3088
rect 34613 3008 34660 3072
rect 34724 3008 34740 3072
rect 34613 2992 34740 3008
rect 28294 2912 28421 2928
rect 28294 2848 28341 2912
rect 28405 2848 28421 2912
rect 28294 2832 28421 2848
rect 28294 2768 28341 2832
rect 28405 2768 28421 2832
rect 28294 2752 28421 2768
rect 28294 2688 28341 2752
rect 28405 2688 28421 2752
rect 28294 2672 28421 2688
rect 28294 2608 28341 2672
rect 28405 2608 28421 2672
rect 28294 2592 28421 2608
rect 28294 2528 28341 2592
rect 28405 2528 28421 2592
rect 28294 2512 28421 2528
rect 28294 2448 28341 2512
rect 28405 2448 28421 2512
rect 28294 2432 28421 2448
rect 28294 2368 28341 2432
rect 28405 2368 28421 2432
rect 28294 2352 28421 2368
rect 28294 2288 28341 2352
rect 28405 2288 28421 2352
rect 28294 2272 28421 2288
rect 28294 2208 28341 2272
rect 28405 2208 28421 2272
rect 28294 2192 28421 2208
rect 28294 2128 28341 2192
rect 28405 2128 28421 2192
rect 28294 2112 28421 2128
rect 28294 2048 28341 2112
rect 28405 2048 28421 2112
rect 28294 2032 28421 2048
rect 28294 1968 28341 2032
rect 28405 1968 28421 2032
rect 28294 1952 28421 1968
rect 28294 1888 28341 1952
rect 28405 1888 28421 1952
rect 28294 1872 28421 1888
rect 28294 1808 28341 1872
rect 28405 1808 28421 1872
rect 28294 1792 28421 1808
rect 28294 1728 28341 1792
rect 28405 1728 28421 1792
rect 28294 1712 28421 1728
rect 28294 1648 28341 1712
rect 28405 1648 28421 1712
rect 28294 1632 28421 1648
rect 28294 1568 28341 1632
rect 28405 1568 28421 1632
rect 28294 1552 28421 1568
rect 28294 1488 28341 1552
rect 28405 1488 28421 1552
rect 28294 1472 28421 1488
rect 28294 1408 28341 1472
rect 28405 1408 28421 1472
rect 28294 1392 28421 1408
rect 28294 1328 28341 1392
rect 28405 1328 28421 1392
rect 28294 1312 28421 1328
rect 28294 1248 28341 1312
rect 28405 1248 28421 1312
rect 28294 1232 28421 1248
rect 28294 1168 28341 1232
rect 28405 1168 28421 1232
rect 28294 1152 28421 1168
rect 28294 1088 28341 1152
rect 28405 1088 28421 1152
rect 28294 1072 28421 1088
rect 28294 1008 28341 1072
rect 28405 1008 28421 1072
rect 28294 992 28421 1008
rect 28294 928 28341 992
rect 28405 928 28421 992
rect 28294 912 28421 928
rect 28294 848 28341 912
rect 28405 848 28421 912
rect 28294 832 28421 848
rect 28294 768 28341 832
rect 28405 768 28421 832
rect 28294 752 28421 768
rect 28294 688 28341 752
rect 28405 688 28421 752
rect 28294 672 28421 688
rect 28294 608 28341 672
rect 28405 608 28421 672
rect 28294 592 28421 608
rect 28294 528 28341 592
rect 28405 528 28421 592
rect 28294 512 28421 528
rect 28294 448 28341 512
rect 28405 448 28421 512
rect 28294 432 28421 448
rect 28294 368 28341 432
rect 28405 368 28421 432
rect 28294 352 28421 368
rect 28294 288 28341 352
rect 28405 288 28421 352
rect 28294 272 28421 288
rect 28294 208 28341 272
rect 28405 208 28421 272
rect 28294 192 28421 208
rect 28294 128 28341 192
rect 28405 128 28421 192
rect 28294 112 28421 128
rect 28294 48 28341 112
rect 28405 48 28421 112
rect 28294 32 28421 48
rect 28294 -32 28341 32
rect 28405 -32 28421 32
rect 28294 -48 28421 -32
rect 28294 -112 28341 -48
rect 28405 -112 28421 -48
rect 28294 -128 28421 -112
rect 28294 -192 28341 -128
rect 28405 -192 28421 -128
rect 28294 -208 28421 -192
rect 28294 -272 28341 -208
rect 28405 -272 28421 -208
rect 28294 -288 28421 -272
rect 28294 -352 28341 -288
rect 28405 -352 28421 -288
rect 28294 -368 28421 -352
rect 28294 -432 28341 -368
rect 28405 -432 28421 -368
rect 28294 -448 28421 -432
rect 28294 -512 28341 -448
rect 28405 -512 28421 -448
rect 28294 -528 28421 -512
rect 28294 -592 28341 -528
rect 28405 -592 28421 -528
rect 28294 -608 28421 -592
rect 28294 -672 28341 -608
rect 28405 -672 28421 -608
rect 28294 -688 28421 -672
rect 28294 -752 28341 -688
rect 28405 -752 28421 -688
rect 28294 -768 28421 -752
rect 28294 -832 28341 -768
rect 28405 -832 28421 -768
rect 28294 -848 28421 -832
rect 28294 -912 28341 -848
rect 28405 -912 28421 -848
rect 28294 -928 28421 -912
rect 28294 -992 28341 -928
rect 28405 -992 28421 -928
rect 28294 -1008 28421 -992
rect 28294 -1072 28341 -1008
rect 28405 -1072 28421 -1008
rect 28294 -1088 28421 -1072
rect 28294 -1152 28341 -1088
rect 28405 -1152 28421 -1088
rect 28294 -1168 28421 -1152
rect 28294 -1232 28341 -1168
rect 28405 -1232 28421 -1168
rect 28294 -1248 28421 -1232
rect 28294 -1312 28341 -1248
rect 28405 -1312 28421 -1248
rect 28294 -1328 28421 -1312
rect 28294 -1392 28341 -1328
rect 28405 -1392 28421 -1328
rect 28294 -1408 28421 -1392
rect 28294 -1472 28341 -1408
rect 28405 -1472 28421 -1408
rect 28294 -1488 28421 -1472
rect 28294 -1552 28341 -1488
rect 28405 -1552 28421 -1488
rect 28294 -1568 28421 -1552
rect 28294 -1632 28341 -1568
rect 28405 -1632 28421 -1568
rect 28294 -1648 28421 -1632
rect 28294 -1712 28341 -1648
rect 28405 -1712 28421 -1648
rect 28294 -1728 28421 -1712
rect 28294 -1792 28341 -1728
rect 28405 -1792 28421 -1728
rect 28294 -1808 28421 -1792
rect 28294 -1872 28341 -1808
rect 28405 -1872 28421 -1808
rect 28294 -1888 28421 -1872
rect 28294 -1952 28341 -1888
rect 28405 -1952 28421 -1888
rect 28294 -1968 28421 -1952
rect 28294 -2032 28341 -1968
rect 28405 -2032 28421 -1968
rect 28294 -2048 28421 -2032
rect 28294 -2112 28341 -2048
rect 28405 -2112 28421 -2048
rect 28294 -2128 28421 -2112
rect 28294 -2192 28341 -2128
rect 28405 -2192 28421 -2128
rect 28294 -2208 28421 -2192
rect 28294 -2272 28341 -2208
rect 28405 -2272 28421 -2208
rect 28294 -2288 28421 -2272
rect 28294 -2352 28341 -2288
rect 28405 -2352 28421 -2288
rect 28294 -2368 28421 -2352
rect 28294 -2432 28341 -2368
rect 28405 -2432 28421 -2368
rect 28294 -2448 28421 -2432
rect 28294 -2512 28341 -2448
rect 28405 -2512 28421 -2448
rect 28294 -2528 28421 -2512
rect 28294 -2592 28341 -2528
rect 28405 -2592 28421 -2528
rect 28294 -2608 28421 -2592
rect 28294 -2672 28341 -2608
rect 28405 -2672 28421 -2608
rect 28294 -2688 28421 -2672
rect 28294 -2752 28341 -2688
rect 28405 -2752 28421 -2688
rect 28294 -2768 28421 -2752
rect 28294 -2832 28341 -2768
rect 28405 -2832 28421 -2768
rect 28294 -2848 28421 -2832
rect 28294 -2912 28341 -2848
rect 28405 -2912 28421 -2848
rect 28294 -2928 28421 -2912
rect 21975 -3008 22102 -2992
rect 21975 -3072 22022 -3008
rect 22086 -3072 22102 -3008
rect 21975 -3088 22102 -3072
rect 21975 -3212 22079 -3088
rect 21975 -3228 22102 -3212
rect 21975 -3292 22022 -3228
rect 22086 -3292 22102 -3228
rect 21975 -3308 22102 -3292
rect 15656 -3388 15783 -3372
rect 15656 -3452 15703 -3388
rect 15767 -3452 15783 -3388
rect 15656 -3468 15783 -3452
rect 15656 -3532 15703 -3468
rect 15767 -3532 15783 -3468
rect 15656 -3548 15783 -3532
rect 15656 -3612 15703 -3548
rect 15767 -3612 15783 -3548
rect 15656 -3628 15783 -3612
rect 15656 -3692 15703 -3628
rect 15767 -3692 15783 -3628
rect 15656 -3708 15783 -3692
rect 15656 -3772 15703 -3708
rect 15767 -3772 15783 -3708
rect 15656 -3788 15783 -3772
rect 15656 -3852 15703 -3788
rect 15767 -3852 15783 -3788
rect 15656 -3868 15783 -3852
rect 15656 -3932 15703 -3868
rect 15767 -3932 15783 -3868
rect 15656 -3948 15783 -3932
rect 15656 -4012 15703 -3948
rect 15767 -4012 15783 -3948
rect 15656 -4028 15783 -4012
rect 15656 -4092 15703 -4028
rect 15767 -4092 15783 -4028
rect 15656 -4108 15783 -4092
rect 15656 -4172 15703 -4108
rect 15767 -4172 15783 -4108
rect 15656 -4188 15783 -4172
rect 15656 -4252 15703 -4188
rect 15767 -4252 15783 -4188
rect 15656 -4268 15783 -4252
rect 15656 -4332 15703 -4268
rect 15767 -4332 15783 -4268
rect 15656 -4348 15783 -4332
rect 15656 -4412 15703 -4348
rect 15767 -4412 15783 -4348
rect 15656 -4428 15783 -4412
rect 15656 -4492 15703 -4428
rect 15767 -4492 15783 -4428
rect 15656 -4508 15783 -4492
rect 15656 -4572 15703 -4508
rect 15767 -4572 15783 -4508
rect 15656 -4588 15783 -4572
rect 15656 -4652 15703 -4588
rect 15767 -4652 15783 -4588
rect 15656 -4668 15783 -4652
rect 15656 -4732 15703 -4668
rect 15767 -4732 15783 -4668
rect 15656 -4748 15783 -4732
rect 15656 -4812 15703 -4748
rect 15767 -4812 15783 -4748
rect 15656 -4828 15783 -4812
rect 15656 -4892 15703 -4828
rect 15767 -4892 15783 -4828
rect 15656 -4908 15783 -4892
rect 15656 -4972 15703 -4908
rect 15767 -4972 15783 -4908
rect 15656 -4988 15783 -4972
rect 15656 -5052 15703 -4988
rect 15767 -5052 15783 -4988
rect 15656 -5068 15783 -5052
rect 15656 -5132 15703 -5068
rect 15767 -5132 15783 -5068
rect 15656 -5148 15783 -5132
rect 15656 -5212 15703 -5148
rect 15767 -5212 15783 -5148
rect 15656 -5228 15783 -5212
rect 15656 -5292 15703 -5228
rect 15767 -5292 15783 -5228
rect 15656 -5308 15783 -5292
rect 15656 -5372 15703 -5308
rect 15767 -5372 15783 -5308
rect 15656 -5388 15783 -5372
rect 15656 -5452 15703 -5388
rect 15767 -5452 15783 -5388
rect 15656 -5468 15783 -5452
rect 15656 -5532 15703 -5468
rect 15767 -5532 15783 -5468
rect 15656 -5548 15783 -5532
rect 15656 -5612 15703 -5548
rect 15767 -5612 15783 -5548
rect 15656 -5628 15783 -5612
rect 15656 -5692 15703 -5628
rect 15767 -5692 15783 -5628
rect 15656 -5708 15783 -5692
rect 15656 -5772 15703 -5708
rect 15767 -5772 15783 -5708
rect 15656 -5788 15783 -5772
rect 15656 -5852 15703 -5788
rect 15767 -5852 15783 -5788
rect 15656 -5868 15783 -5852
rect 15656 -5932 15703 -5868
rect 15767 -5932 15783 -5868
rect 15656 -5948 15783 -5932
rect 15656 -6012 15703 -5948
rect 15767 -6012 15783 -5948
rect 15656 -6028 15783 -6012
rect 15656 -6092 15703 -6028
rect 15767 -6092 15783 -6028
rect 15656 -6108 15783 -6092
rect 15656 -6172 15703 -6108
rect 15767 -6172 15783 -6108
rect 15656 -6188 15783 -6172
rect 15656 -6252 15703 -6188
rect 15767 -6252 15783 -6188
rect 15656 -6268 15783 -6252
rect 15656 -6332 15703 -6268
rect 15767 -6332 15783 -6268
rect 15656 -6348 15783 -6332
rect 15656 -6412 15703 -6348
rect 15767 -6412 15783 -6348
rect 15656 -6428 15783 -6412
rect 15656 -6492 15703 -6428
rect 15767 -6492 15783 -6428
rect 15656 -6508 15783 -6492
rect 15656 -6572 15703 -6508
rect 15767 -6572 15783 -6508
rect 15656 -6588 15783 -6572
rect 15656 -6652 15703 -6588
rect 15767 -6652 15783 -6588
rect 15656 -6668 15783 -6652
rect 15656 -6732 15703 -6668
rect 15767 -6732 15783 -6668
rect 15656 -6748 15783 -6732
rect 15656 -6812 15703 -6748
rect 15767 -6812 15783 -6748
rect 15656 -6828 15783 -6812
rect 15656 -6892 15703 -6828
rect 15767 -6892 15783 -6828
rect 15656 -6908 15783 -6892
rect 15656 -6972 15703 -6908
rect 15767 -6972 15783 -6908
rect 15656 -6988 15783 -6972
rect 15656 -7052 15703 -6988
rect 15767 -7052 15783 -6988
rect 15656 -7068 15783 -7052
rect 15656 -7132 15703 -7068
rect 15767 -7132 15783 -7068
rect 15656 -7148 15783 -7132
rect 15656 -7212 15703 -7148
rect 15767 -7212 15783 -7148
rect 15656 -7228 15783 -7212
rect 15656 -7292 15703 -7228
rect 15767 -7292 15783 -7228
rect 15656 -7308 15783 -7292
rect 15656 -7372 15703 -7308
rect 15767 -7372 15783 -7308
rect 15656 -7388 15783 -7372
rect 15656 -7452 15703 -7388
rect 15767 -7452 15783 -7388
rect 15656 -7468 15783 -7452
rect 15656 -7532 15703 -7468
rect 15767 -7532 15783 -7468
rect 15656 -7548 15783 -7532
rect 15656 -7612 15703 -7548
rect 15767 -7612 15783 -7548
rect 15656 -7628 15783 -7612
rect 15656 -7692 15703 -7628
rect 15767 -7692 15783 -7628
rect 15656 -7708 15783 -7692
rect 15656 -7772 15703 -7708
rect 15767 -7772 15783 -7708
rect 15656 -7788 15783 -7772
rect 15656 -7852 15703 -7788
rect 15767 -7852 15783 -7788
rect 15656 -7868 15783 -7852
rect 15656 -7932 15703 -7868
rect 15767 -7932 15783 -7868
rect 15656 -7948 15783 -7932
rect 15656 -8012 15703 -7948
rect 15767 -8012 15783 -7948
rect 15656 -8028 15783 -8012
rect 15656 -8092 15703 -8028
rect 15767 -8092 15783 -8028
rect 15656 -8108 15783 -8092
rect 15656 -8172 15703 -8108
rect 15767 -8172 15783 -8108
rect 15656 -8188 15783 -8172
rect 15656 -8252 15703 -8188
rect 15767 -8252 15783 -8188
rect 15656 -8268 15783 -8252
rect 15656 -8332 15703 -8268
rect 15767 -8332 15783 -8268
rect 15656 -8348 15783 -8332
rect 15656 -8412 15703 -8348
rect 15767 -8412 15783 -8348
rect 15656 -8428 15783 -8412
rect 15656 -8492 15703 -8428
rect 15767 -8492 15783 -8428
rect 15656 -8508 15783 -8492
rect 15656 -8572 15703 -8508
rect 15767 -8572 15783 -8508
rect 15656 -8588 15783 -8572
rect 15656 -8652 15703 -8588
rect 15767 -8652 15783 -8588
rect 15656 -8668 15783 -8652
rect 15656 -8732 15703 -8668
rect 15767 -8732 15783 -8668
rect 15656 -8748 15783 -8732
rect 15656 -8812 15703 -8748
rect 15767 -8812 15783 -8748
rect 15656 -8828 15783 -8812
rect 15656 -8892 15703 -8828
rect 15767 -8892 15783 -8828
rect 15656 -8908 15783 -8892
rect 15656 -8972 15703 -8908
rect 15767 -8972 15783 -8908
rect 15656 -8988 15783 -8972
rect 15656 -9052 15703 -8988
rect 15767 -9052 15783 -8988
rect 15656 -9068 15783 -9052
rect 15656 -9132 15703 -9068
rect 15767 -9132 15783 -9068
rect 15656 -9148 15783 -9132
rect 15656 -9212 15703 -9148
rect 15767 -9212 15783 -9148
rect 15656 -9228 15783 -9212
rect 9337 -9308 9464 -9292
rect 9337 -9372 9384 -9308
rect 9448 -9372 9464 -9308
rect 9337 -9388 9464 -9372
rect 9337 -9512 9441 -9388
rect 9337 -9528 9464 -9512
rect 9337 -9592 9384 -9528
rect 9448 -9592 9464 -9528
rect 9337 -9608 9464 -9592
rect 3018 -9688 3145 -9672
rect 3018 -9752 3065 -9688
rect 3129 -9752 3145 -9688
rect 3018 -9768 3145 -9752
rect 3018 -9832 3065 -9768
rect 3129 -9832 3145 -9768
rect 3018 -9848 3145 -9832
rect 3018 -9912 3065 -9848
rect 3129 -9912 3145 -9848
rect 3018 -9928 3145 -9912
rect 3018 -9992 3065 -9928
rect 3129 -9992 3145 -9928
rect 3018 -10008 3145 -9992
rect 3018 -10072 3065 -10008
rect 3129 -10072 3145 -10008
rect 3018 -10088 3145 -10072
rect 3018 -10152 3065 -10088
rect 3129 -10152 3145 -10088
rect 3018 -10168 3145 -10152
rect 3018 -10232 3065 -10168
rect 3129 -10232 3145 -10168
rect 3018 -10248 3145 -10232
rect 3018 -10312 3065 -10248
rect 3129 -10312 3145 -10248
rect 3018 -10328 3145 -10312
rect 3018 -10392 3065 -10328
rect 3129 -10392 3145 -10328
rect 3018 -10408 3145 -10392
rect 3018 -10472 3065 -10408
rect 3129 -10472 3145 -10408
rect 3018 -10488 3145 -10472
rect 3018 -10552 3065 -10488
rect 3129 -10552 3145 -10488
rect 3018 -10568 3145 -10552
rect 3018 -10632 3065 -10568
rect 3129 -10632 3145 -10568
rect 3018 -10648 3145 -10632
rect 3018 -10712 3065 -10648
rect 3129 -10712 3145 -10648
rect 3018 -10728 3145 -10712
rect 3018 -10792 3065 -10728
rect 3129 -10792 3145 -10728
rect 3018 -10808 3145 -10792
rect 3018 -10872 3065 -10808
rect 3129 -10872 3145 -10808
rect 3018 -10888 3145 -10872
rect 3018 -10952 3065 -10888
rect 3129 -10952 3145 -10888
rect 3018 -10968 3145 -10952
rect 3018 -11032 3065 -10968
rect 3129 -11032 3145 -10968
rect 3018 -11048 3145 -11032
rect 3018 -11112 3065 -11048
rect 3129 -11112 3145 -11048
rect 3018 -11128 3145 -11112
rect 3018 -11192 3065 -11128
rect 3129 -11192 3145 -11128
rect 3018 -11208 3145 -11192
rect 3018 -11272 3065 -11208
rect 3129 -11272 3145 -11208
rect 3018 -11288 3145 -11272
rect 3018 -11352 3065 -11288
rect 3129 -11352 3145 -11288
rect 3018 -11368 3145 -11352
rect 3018 -11432 3065 -11368
rect 3129 -11432 3145 -11368
rect 3018 -11448 3145 -11432
rect 3018 -11512 3065 -11448
rect 3129 -11512 3145 -11448
rect 3018 -11528 3145 -11512
rect 3018 -11592 3065 -11528
rect 3129 -11592 3145 -11528
rect 3018 -11608 3145 -11592
rect 3018 -11672 3065 -11608
rect 3129 -11672 3145 -11608
rect 3018 -11688 3145 -11672
rect 3018 -11752 3065 -11688
rect 3129 -11752 3145 -11688
rect 3018 -11768 3145 -11752
rect 3018 -11832 3065 -11768
rect 3129 -11832 3145 -11768
rect 3018 -11848 3145 -11832
rect 3018 -11912 3065 -11848
rect 3129 -11912 3145 -11848
rect 3018 -11928 3145 -11912
rect 3018 -11992 3065 -11928
rect 3129 -11992 3145 -11928
rect 3018 -12008 3145 -11992
rect 3018 -12072 3065 -12008
rect 3129 -12072 3145 -12008
rect 3018 -12088 3145 -12072
rect 3018 -12152 3065 -12088
rect 3129 -12152 3145 -12088
rect 3018 -12168 3145 -12152
rect 3018 -12232 3065 -12168
rect 3129 -12232 3145 -12168
rect 3018 -12248 3145 -12232
rect 3018 -12312 3065 -12248
rect 3129 -12312 3145 -12248
rect 3018 -12328 3145 -12312
rect 3018 -12392 3065 -12328
rect 3129 -12392 3145 -12328
rect 3018 -12408 3145 -12392
rect 3018 -12472 3065 -12408
rect 3129 -12472 3145 -12408
rect 3018 -12488 3145 -12472
rect 3018 -12552 3065 -12488
rect 3129 -12552 3145 -12488
rect 3018 -12568 3145 -12552
rect 3018 -12632 3065 -12568
rect 3129 -12632 3145 -12568
rect 3018 -12648 3145 -12632
rect 3018 -12712 3065 -12648
rect 3129 -12712 3145 -12648
rect 3018 -12728 3145 -12712
rect 3018 -12792 3065 -12728
rect 3129 -12792 3145 -12728
rect 3018 -12808 3145 -12792
rect 3018 -12872 3065 -12808
rect 3129 -12872 3145 -12808
rect 3018 -12888 3145 -12872
rect 3018 -12952 3065 -12888
rect 3129 -12952 3145 -12888
rect 3018 -12968 3145 -12952
rect 3018 -13032 3065 -12968
rect 3129 -13032 3145 -12968
rect 3018 -13048 3145 -13032
rect 3018 -13112 3065 -13048
rect 3129 -13112 3145 -13048
rect 3018 -13128 3145 -13112
rect 3018 -13192 3065 -13128
rect 3129 -13192 3145 -13128
rect 3018 -13208 3145 -13192
rect 3018 -13272 3065 -13208
rect 3129 -13272 3145 -13208
rect 3018 -13288 3145 -13272
rect 3018 -13352 3065 -13288
rect 3129 -13352 3145 -13288
rect 3018 -13368 3145 -13352
rect 3018 -13432 3065 -13368
rect 3129 -13432 3145 -13368
rect 3018 -13448 3145 -13432
rect 3018 -13512 3065 -13448
rect 3129 -13512 3145 -13448
rect 3018 -13528 3145 -13512
rect 3018 -13592 3065 -13528
rect 3129 -13592 3145 -13528
rect 3018 -13608 3145 -13592
rect 3018 -13672 3065 -13608
rect 3129 -13672 3145 -13608
rect 3018 -13688 3145 -13672
rect 3018 -13752 3065 -13688
rect 3129 -13752 3145 -13688
rect 3018 -13768 3145 -13752
rect 3018 -13832 3065 -13768
rect 3129 -13832 3145 -13768
rect 3018 -13848 3145 -13832
rect 3018 -13912 3065 -13848
rect 3129 -13912 3145 -13848
rect 3018 -13928 3145 -13912
rect 3018 -13992 3065 -13928
rect 3129 -13992 3145 -13928
rect 3018 -14008 3145 -13992
rect 3018 -14072 3065 -14008
rect 3129 -14072 3145 -14008
rect 3018 -14088 3145 -14072
rect 3018 -14152 3065 -14088
rect 3129 -14152 3145 -14088
rect 3018 -14168 3145 -14152
rect 3018 -14232 3065 -14168
rect 3129 -14232 3145 -14168
rect 3018 -14248 3145 -14232
rect 3018 -14312 3065 -14248
rect 3129 -14312 3145 -14248
rect 3018 -14328 3145 -14312
rect 3018 -14392 3065 -14328
rect 3129 -14392 3145 -14328
rect 3018 -14408 3145 -14392
rect 3018 -14472 3065 -14408
rect 3129 -14472 3145 -14408
rect 3018 -14488 3145 -14472
rect 3018 -14552 3065 -14488
rect 3129 -14552 3145 -14488
rect 3018 -14568 3145 -14552
rect 3018 -14632 3065 -14568
rect 3129 -14632 3145 -14568
rect 3018 -14648 3145 -14632
rect 3018 -14712 3065 -14648
rect 3129 -14712 3145 -14648
rect 3018 -14728 3145 -14712
rect 3018 -14792 3065 -14728
rect 3129 -14792 3145 -14728
rect 3018 -14808 3145 -14792
rect 3018 -14872 3065 -14808
rect 3129 -14872 3145 -14808
rect 3018 -14888 3145 -14872
rect 3018 -14952 3065 -14888
rect 3129 -14952 3145 -14888
rect 3018 -14968 3145 -14952
rect 3018 -15032 3065 -14968
rect 3129 -15032 3145 -14968
rect 3018 -15048 3145 -15032
rect 3018 -15112 3065 -15048
rect 3129 -15112 3145 -15048
rect 3018 -15128 3145 -15112
rect 3018 -15192 3065 -15128
rect 3129 -15192 3145 -15128
rect 3018 -15208 3145 -15192
rect 3018 -15272 3065 -15208
rect 3129 -15272 3145 -15208
rect 3018 -15288 3145 -15272
rect 3018 -15352 3065 -15288
rect 3129 -15352 3145 -15288
rect 3018 -15368 3145 -15352
rect 3018 -15432 3065 -15368
rect 3129 -15432 3145 -15368
rect 3018 -15448 3145 -15432
rect 3018 -15512 3065 -15448
rect 3129 -15512 3145 -15448
rect 3018 -15528 3145 -15512
rect -3301 -15608 -3174 -15592
rect -3301 -15672 -3254 -15608
rect -3190 -15672 -3174 -15608
rect -3301 -15688 -3174 -15672
rect -3301 -15812 -3197 -15688
rect -3301 -15828 -3174 -15812
rect -3301 -15892 -3254 -15828
rect -3190 -15892 -3174 -15828
rect -3301 -15908 -3174 -15892
rect -9620 -15988 -9493 -15972
rect -9620 -16052 -9573 -15988
rect -9509 -16052 -9493 -15988
rect -9620 -16068 -9493 -16052
rect -9620 -16132 -9573 -16068
rect -9509 -16132 -9493 -16068
rect -9620 -16148 -9493 -16132
rect -9620 -16212 -9573 -16148
rect -9509 -16212 -9493 -16148
rect -9620 -16228 -9493 -16212
rect -9620 -16292 -9573 -16228
rect -9509 -16292 -9493 -16228
rect -9620 -16308 -9493 -16292
rect -9620 -16372 -9573 -16308
rect -9509 -16372 -9493 -16308
rect -9620 -16388 -9493 -16372
rect -9620 -16452 -9573 -16388
rect -9509 -16452 -9493 -16388
rect -9620 -16468 -9493 -16452
rect -9620 -16532 -9573 -16468
rect -9509 -16532 -9493 -16468
rect -9620 -16548 -9493 -16532
rect -9620 -16612 -9573 -16548
rect -9509 -16612 -9493 -16548
rect -9620 -16628 -9493 -16612
rect -9620 -16692 -9573 -16628
rect -9509 -16692 -9493 -16628
rect -9620 -16708 -9493 -16692
rect -9620 -16772 -9573 -16708
rect -9509 -16772 -9493 -16708
rect -9620 -16788 -9493 -16772
rect -9620 -16852 -9573 -16788
rect -9509 -16852 -9493 -16788
rect -9620 -16868 -9493 -16852
rect -9620 -16932 -9573 -16868
rect -9509 -16932 -9493 -16868
rect -9620 -16948 -9493 -16932
rect -9620 -17012 -9573 -16948
rect -9509 -17012 -9493 -16948
rect -9620 -17028 -9493 -17012
rect -9620 -17092 -9573 -17028
rect -9509 -17092 -9493 -17028
rect -9620 -17108 -9493 -17092
rect -9620 -17172 -9573 -17108
rect -9509 -17172 -9493 -17108
rect -9620 -17188 -9493 -17172
rect -9620 -17252 -9573 -17188
rect -9509 -17252 -9493 -17188
rect -9620 -17268 -9493 -17252
rect -9620 -17332 -9573 -17268
rect -9509 -17332 -9493 -17268
rect -9620 -17348 -9493 -17332
rect -9620 -17412 -9573 -17348
rect -9509 -17412 -9493 -17348
rect -9620 -17428 -9493 -17412
rect -9620 -17492 -9573 -17428
rect -9509 -17492 -9493 -17428
rect -9620 -17508 -9493 -17492
rect -9620 -17572 -9573 -17508
rect -9509 -17572 -9493 -17508
rect -9620 -17588 -9493 -17572
rect -9620 -17652 -9573 -17588
rect -9509 -17652 -9493 -17588
rect -9620 -17668 -9493 -17652
rect -9620 -17732 -9573 -17668
rect -9509 -17732 -9493 -17668
rect -9620 -17748 -9493 -17732
rect -9620 -17812 -9573 -17748
rect -9509 -17812 -9493 -17748
rect -9620 -17828 -9493 -17812
rect -9620 -17892 -9573 -17828
rect -9509 -17892 -9493 -17828
rect -9620 -17908 -9493 -17892
rect -9620 -17972 -9573 -17908
rect -9509 -17972 -9493 -17908
rect -9620 -17988 -9493 -17972
rect -9620 -18052 -9573 -17988
rect -9509 -18052 -9493 -17988
rect -9620 -18068 -9493 -18052
rect -9620 -18132 -9573 -18068
rect -9509 -18132 -9493 -18068
rect -9620 -18148 -9493 -18132
rect -9620 -18212 -9573 -18148
rect -9509 -18212 -9493 -18148
rect -9620 -18228 -9493 -18212
rect -9620 -18292 -9573 -18228
rect -9509 -18292 -9493 -18228
rect -9620 -18308 -9493 -18292
rect -9620 -18372 -9573 -18308
rect -9509 -18372 -9493 -18308
rect -9620 -18388 -9493 -18372
rect -9620 -18452 -9573 -18388
rect -9509 -18452 -9493 -18388
rect -9620 -18468 -9493 -18452
rect -9620 -18532 -9573 -18468
rect -9509 -18532 -9493 -18468
rect -9620 -18548 -9493 -18532
rect -9620 -18612 -9573 -18548
rect -9509 -18612 -9493 -18548
rect -9620 -18628 -9493 -18612
rect -9620 -18692 -9573 -18628
rect -9509 -18692 -9493 -18628
rect -9620 -18708 -9493 -18692
rect -9620 -18772 -9573 -18708
rect -9509 -18772 -9493 -18708
rect -9620 -18788 -9493 -18772
rect -9620 -18852 -9573 -18788
rect -9509 -18852 -9493 -18788
rect -9620 -18868 -9493 -18852
rect -9620 -18932 -9573 -18868
rect -9509 -18932 -9493 -18868
rect -9620 -18948 -9493 -18932
rect -9620 -19012 -9573 -18948
rect -9509 -19012 -9493 -18948
rect -9620 -19028 -9493 -19012
rect -9620 -19092 -9573 -19028
rect -9509 -19092 -9493 -19028
rect -9620 -19108 -9493 -19092
rect -9620 -19172 -9573 -19108
rect -9509 -19172 -9493 -19108
rect -9620 -19188 -9493 -19172
rect -9620 -19252 -9573 -19188
rect -9509 -19252 -9493 -19188
rect -9620 -19268 -9493 -19252
rect -9620 -19332 -9573 -19268
rect -9509 -19332 -9493 -19268
rect -9620 -19348 -9493 -19332
rect -9620 -19412 -9573 -19348
rect -9509 -19412 -9493 -19348
rect -9620 -19428 -9493 -19412
rect -9620 -19492 -9573 -19428
rect -9509 -19492 -9493 -19428
rect -9620 -19508 -9493 -19492
rect -9620 -19572 -9573 -19508
rect -9509 -19572 -9493 -19508
rect -9620 -19588 -9493 -19572
rect -9620 -19652 -9573 -19588
rect -9509 -19652 -9493 -19588
rect -9620 -19668 -9493 -19652
rect -9620 -19732 -9573 -19668
rect -9509 -19732 -9493 -19668
rect -9620 -19748 -9493 -19732
rect -9620 -19812 -9573 -19748
rect -9509 -19812 -9493 -19748
rect -9620 -19828 -9493 -19812
rect -9620 -19892 -9573 -19828
rect -9509 -19892 -9493 -19828
rect -9620 -19908 -9493 -19892
rect -9620 -19972 -9573 -19908
rect -9509 -19972 -9493 -19908
rect -9620 -19988 -9493 -19972
rect -9620 -20052 -9573 -19988
rect -9509 -20052 -9493 -19988
rect -9620 -20068 -9493 -20052
rect -9620 -20132 -9573 -20068
rect -9509 -20132 -9493 -20068
rect -9620 -20148 -9493 -20132
rect -9620 -20212 -9573 -20148
rect -9509 -20212 -9493 -20148
rect -9620 -20228 -9493 -20212
rect -9620 -20292 -9573 -20228
rect -9509 -20292 -9493 -20228
rect -9620 -20308 -9493 -20292
rect -9620 -20372 -9573 -20308
rect -9509 -20372 -9493 -20308
rect -9620 -20388 -9493 -20372
rect -9620 -20452 -9573 -20388
rect -9509 -20452 -9493 -20388
rect -9620 -20468 -9493 -20452
rect -9620 -20532 -9573 -20468
rect -9509 -20532 -9493 -20468
rect -9620 -20548 -9493 -20532
rect -9620 -20612 -9573 -20548
rect -9509 -20612 -9493 -20548
rect -9620 -20628 -9493 -20612
rect -9620 -20692 -9573 -20628
rect -9509 -20692 -9493 -20628
rect -9620 -20708 -9493 -20692
rect -9620 -20772 -9573 -20708
rect -9509 -20772 -9493 -20708
rect -9620 -20788 -9493 -20772
rect -9620 -20852 -9573 -20788
rect -9509 -20852 -9493 -20788
rect -9620 -20868 -9493 -20852
rect -9620 -20932 -9573 -20868
rect -9509 -20932 -9493 -20868
rect -9620 -20948 -9493 -20932
rect -9620 -21012 -9573 -20948
rect -9509 -21012 -9493 -20948
rect -9620 -21028 -9493 -21012
rect -9620 -21092 -9573 -21028
rect -9509 -21092 -9493 -21028
rect -9620 -21108 -9493 -21092
rect -9620 -21172 -9573 -21108
rect -9509 -21172 -9493 -21108
rect -9620 -21188 -9493 -21172
rect -9620 -21252 -9573 -21188
rect -9509 -21252 -9493 -21188
rect -9620 -21268 -9493 -21252
rect -9620 -21332 -9573 -21268
rect -9509 -21332 -9493 -21268
rect -9620 -21348 -9493 -21332
rect -9620 -21412 -9573 -21348
rect -9509 -21412 -9493 -21348
rect -9620 -21428 -9493 -21412
rect -9620 -21492 -9573 -21428
rect -9509 -21492 -9493 -21428
rect -9620 -21508 -9493 -21492
rect -9620 -21572 -9573 -21508
rect -9509 -21572 -9493 -21508
rect -9620 -21588 -9493 -21572
rect -9620 -21652 -9573 -21588
rect -9509 -21652 -9493 -21588
rect -9620 -21668 -9493 -21652
rect -9620 -21732 -9573 -21668
rect -9509 -21732 -9493 -21668
rect -9620 -21748 -9493 -21732
rect -9620 -21812 -9573 -21748
rect -9509 -21812 -9493 -21748
rect -9620 -21828 -9493 -21812
rect -15939 -21908 -15812 -21892
rect -15939 -21972 -15892 -21908
rect -15828 -21972 -15812 -21908
rect -15939 -21988 -15812 -21972
rect -15939 -22112 -15835 -21988
rect -15939 -22128 -15812 -22112
rect -15939 -22192 -15892 -22128
rect -15828 -22192 -15812 -22128
rect -15939 -22208 -15812 -22192
rect -22258 -22288 -22131 -22272
rect -22258 -22352 -22211 -22288
rect -22147 -22352 -22131 -22288
rect -22258 -22368 -22131 -22352
rect -22258 -22432 -22211 -22368
rect -22147 -22432 -22131 -22368
rect -22258 -22448 -22131 -22432
rect -22258 -22512 -22211 -22448
rect -22147 -22512 -22131 -22448
rect -22258 -22528 -22131 -22512
rect -22258 -22592 -22211 -22528
rect -22147 -22592 -22131 -22528
rect -22258 -22608 -22131 -22592
rect -22258 -22672 -22211 -22608
rect -22147 -22672 -22131 -22608
rect -22258 -22688 -22131 -22672
rect -22258 -22752 -22211 -22688
rect -22147 -22752 -22131 -22688
rect -22258 -22768 -22131 -22752
rect -22258 -22832 -22211 -22768
rect -22147 -22832 -22131 -22768
rect -22258 -22848 -22131 -22832
rect -22258 -22912 -22211 -22848
rect -22147 -22912 -22131 -22848
rect -22258 -22928 -22131 -22912
rect -22258 -22992 -22211 -22928
rect -22147 -22992 -22131 -22928
rect -22258 -23008 -22131 -22992
rect -22258 -23072 -22211 -23008
rect -22147 -23072 -22131 -23008
rect -22258 -23088 -22131 -23072
rect -22258 -23152 -22211 -23088
rect -22147 -23152 -22131 -23088
rect -22258 -23168 -22131 -23152
rect -22258 -23232 -22211 -23168
rect -22147 -23232 -22131 -23168
rect -22258 -23248 -22131 -23232
rect -22258 -23312 -22211 -23248
rect -22147 -23312 -22131 -23248
rect -22258 -23328 -22131 -23312
rect -22258 -23392 -22211 -23328
rect -22147 -23392 -22131 -23328
rect -22258 -23408 -22131 -23392
rect -22258 -23472 -22211 -23408
rect -22147 -23472 -22131 -23408
rect -22258 -23488 -22131 -23472
rect -22258 -23552 -22211 -23488
rect -22147 -23552 -22131 -23488
rect -22258 -23568 -22131 -23552
rect -22258 -23632 -22211 -23568
rect -22147 -23632 -22131 -23568
rect -22258 -23648 -22131 -23632
rect -22258 -23712 -22211 -23648
rect -22147 -23712 -22131 -23648
rect -22258 -23728 -22131 -23712
rect -22258 -23792 -22211 -23728
rect -22147 -23792 -22131 -23728
rect -22258 -23808 -22131 -23792
rect -22258 -23872 -22211 -23808
rect -22147 -23872 -22131 -23808
rect -22258 -23888 -22131 -23872
rect -22258 -23952 -22211 -23888
rect -22147 -23952 -22131 -23888
rect -22258 -23968 -22131 -23952
rect -22258 -24032 -22211 -23968
rect -22147 -24032 -22131 -23968
rect -22258 -24048 -22131 -24032
rect -22258 -24112 -22211 -24048
rect -22147 -24112 -22131 -24048
rect -22258 -24128 -22131 -24112
rect -22258 -24192 -22211 -24128
rect -22147 -24192 -22131 -24128
rect -22258 -24208 -22131 -24192
rect -22258 -24272 -22211 -24208
rect -22147 -24272 -22131 -24208
rect -22258 -24288 -22131 -24272
rect -22258 -24352 -22211 -24288
rect -22147 -24352 -22131 -24288
rect -22258 -24368 -22131 -24352
rect -22258 -24432 -22211 -24368
rect -22147 -24432 -22131 -24368
rect -22258 -24448 -22131 -24432
rect -22258 -24512 -22211 -24448
rect -22147 -24512 -22131 -24448
rect -22258 -24528 -22131 -24512
rect -22258 -24592 -22211 -24528
rect -22147 -24592 -22131 -24528
rect -22258 -24608 -22131 -24592
rect -22258 -24672 -22211 -24608
rect -22147 -24672 -22131 -24608
rect -22258 -24688 -22131 -24672
rect -22258 -24752 -22211 -24688
rect -22147 -24752 -22131 -24688
rect -22258 -24768 -22131 -24752
rect -22258 -24832 -22211 -24768
rect -22147 -24832 -22131 -24768
rect -22258 -24848 -22131 -24832
rect -22258 -24912 -22211 -24848
rect -22147 -24912 -22131 -24848
rect -22258 -24928 -22131 -24912
rect -22258 -24992 -22211 -24928
rect -22147 -24992 -22131 -24928
rect -22258 -25008 -22131 -24992
rect -22258 -25072 -22211 -25008
rect -22147 -25072 -22131 -25008
rect -22258 -25088 -22131 -25072
rect -22258 -25152 -22211 -25088
rect -22147 -25152 -22131 -25088
rect -22258 -25168 -22131 -25152
rect -22258 -25232 -22211 -25168
rect -22147 -25232 -22131 -25168
rect -22258 -25248 -22131 -25232
rect -22258 -25312 -22211 -25248
rect -22147 -25312 -22131 -25248
rect -22258 -25328 -22131 -25312
rect -22258 -25392 -22211 -25328
rect -22147 -25392 -22131 -25328
rect -22258 -25408 -22131 -25392
rect -22258 -25472 -22211 -25408
rect -22147 -25472 -22131 -25408
rect -22258 -25488 -22131 -25472
rect -22258 -25552 -22211 -25488
rect -22147 -25552 -22131 -25488
rect -22258 -25568 -22131 -25552
rect -22258 -25632 -22211 -25568
rect -22147 -25632 -22131 -25568
rect -22258 -25648 -22131 -25632
rect -22258 -25712 -22211 -25648
rect -22147 -25712 -22131 -25648
rect -22258 -25728 -22131 -25712
rect -22258 -25792 -22211 -25728
rect -22147 -25792 -22131 -25728
rect -22258 -25808 -22131 -25792
rect -22258 -25872 -22211 -25808
rect -22147 -25872 -22131 -25808
rect -22258 -25888 -22131 -25872
rect -22258 -25952 -22211 -25888
rect -22147 -25952 -22131 -25888
rect -22258 -25968 -22131 -25952
rect -22258 -26032 -22211 -25968
rect -22147 -26032 -22131 -25968
rect -22258 -26048 -22131 -26032
rect -22258 -26112 -22211 -26048
rect -22147 -26112 -22131 -26048
rect -22258 -26128 -22131 -26112
rect -22258 -26192 -22211 -26128
rect -22147 -26192 -22131 -26128
rect -22258 -26208 -22131 -26192
rect -22258 -26272 -22211 -26208
rect -22147 -26272 -22131 -26208
rect -22258 -26288 -22131 -26272
rect -22258 -26352 -22211 -26288
rect -22147 -26352 -22131 -26288
rect -22258 -26368 -22131 -26352
rect -22258 -26432 -22211 -26368
rect -22147 -26432 -22131 -26368
rect -22258 -26448 -22131 -26432
rect -22258 -26512 -22211 -26448
rect -22147 -26512 -22131 -26448
rect -22258 -26528 -22131 -26512
rect -22258 -26592 -22211 -26528
rect -22147 -26592 -22131 -26528
rect -22258 -26608 -22131 -26592
rect -22258 -26672 -22211 -26608
rect -22147 -26672 -22131 -26608
rect -22258 -26688 -22131 -26672
rect -22258 -26752 -22211 -26688
rect -22147 -26752 -22131 -26688
rect -22258 -26768 -22131 -26752
rect -22258 -26832 -22211 -26768
rect -22147 -26832 -22131 -26768
rect -22258 -26848 -22131 -26832
rect -22258 -26912 -22211 -26848
rect -22147 -26912 -22131 -26848
rect -22258 -26928 -22131 -26912
rect -22258 -26992 -22211 -26928
rect -22147 -26992 -22131 -26928
rect -22258 -27008 -22131 -26992
rect -22258 -27072 -22211 -27008
rect -22147 -27072 -22131 -27008
rect -22258 -27088 -22131 -27072
rect -22258 -27152 -22211 -27088
rect -22147 -27152 -22131 -27088
rect -22258 -27168 -22131 -27152
rect -22258 -27232 -22211 -27168
rect -22147 -27232 -22131 -27168
rect -22258 -27248 -22131 -27232
rect -22258 -27312 -22211 -27248
rect -22147 -27312 -22131 -27248
rect -22258 -27328 -22131 -27312
rect -22258 -27392 -22211 -27328
rect -22147 -27392 -22131 -27328
rect -22258 -27408 -22131 -27392
rect -22258 -27472 -22211 -27408
rect -22147 -27472 -22131 -27408
rect -22258 -27488 -22131 -27472
rect -22258 -27552 -22211 -27488
rect -22147 -27552 -22131 -27488
rect -22258 -27568 -22131 -27552
rect -22258 -27632 -22211 -27568
rect -22147 -27632 -22131 -27568
rect -22258 -27648 -22131 -27632
rect -22258 -27712 -22211 -27648
rect -22147 -27712 -22131 -27648
rect -22258 -27728 -22131 -27712
rect -22258 -27792 -22211 -27728
rect -22147 -27792 -22131 -27728
rect -22258 -27808 -22131 -27792
rect -22258 -27872 -22211 -27808
rect -22147 -27872 -22131 -27808
rect -22258 -27888 -22131 -27872
rect -22258 -27952 -22211 -27888
rect -22147 -27952 -22131 -27888
rect -22258 -27968 -22131 -27952
rect -22258 -28032 -22211 -27968
rect -22147 -28032 -22131 -27968
rect -22258 -28048 -22131 -28032
rect -22258 -28112 -22211 -28048
rect -22147 -28112 -22131 -28048
rect -22258 -28128 -22131 -28112
rect -28577 -28208 -28450 -28192
rect -28577 -28272 -28530 -28208
rect -28466 -28272 -28450 -28208
rect -28577 -28288 -28450 -28272
rect -28577 -28412 -28473 -28288
rect -28577 -28428 -28450 -28412
rect -28577 -28492 -28530 -28428
rect -28466 -28492 -28450 -28428
rect -28577 -28508 -28450 -28492
rect -34896 -28588 -34769 -28572
rect -34896 -28652 -34849 -28588
rect -34785 -28652 -34769 -28588
rect -34896 -28668 -34769 -28652
rect -34896 -28732 -34849 -28668
rect -34785 -28732 -34769 -28668
rect -34896 -28748 -34769 -28732
rect -34896 -28812 -34849 -28748
rect -34785 -28812 -34769 -28748
rect -34896 -28828 -34769 -28812
rect -34896 -28892 -34849 -28828
rect -34785 -28892 -34769 -28828
rect -34896 -28908 -34769 -28892
rect -34896 -28972 -34849 -28908
rect -34785 -28972 -34769 -28908
rect -34896 -28988 -34769 -28972
rect -34896 -29052 -34849 -28988
rect -34785 -29052 -34769 -28988
rect -34896 -29068 -34769 -29052
rect -34896 -29132 -34849 -29068
rect -34785 -29132 -34769 -29068
rect -34896 -29148 -34769 -29132
rect -34896 -29212 -34849 -29148
rect -34785 -29212 -34769 -29148
rect -34896 -29228 -34769 -29212
rect -34896 -29292 -34849 -29228
rect -34785 -29292 -34769 -29228
rect -34896 -29308 -34769 -29292
rect -34896 -29372 -34849 -29308
rect -34785 -29372 -34769 -29308
rect -34896 -29388 -34769 -29372
rect -34896 -29452 -34849 -29388
rect -34785 -29452 -34769 -29388
rect -34896 -29468 -34769 -29452
rect -34896 -29532 -34849 -29468
rect -34785 -29532 -34769 -29468
rect -34896 -29548 -34769 -29532
rect -34896 -29612 -34849 -29548
rect -34785 -29612 -34769 -29548
rect -34896 -29628 -34769 -29612
rect -34896 -29692 -34849 -29628
rect -34785 -29692 -34769 -29628
rect -34896 -29708 -34769 -29692
rect -34896 -29772 -34849 -29708
rect -34785 -29772 -34769 -29708
rect -34896 -29788 -34769 -29772
rect -34896 -29852 -34849 -29788
rect -34785 -29852 -34769 -29788
rect -34896 -29868 -34769 -29852
rect -34896 -29932 -34849 -29868
rect -34785 -29932 -34769 -29868
rect -34896 -29948 -34769 -29932
rect -34896 -30012 -34849 -29948
rect -34785 -30012 -34769 -29948
rect -34896 -30028 -34769 -30012
rect -34896 -30092 -34849 -30028
rect -34785 -30092 -34769 -30028
rect -34896 -30108 -34769 -30092
rect -34896 -30172 -34849 -30108
rect -34785 -30172 -34769 -30108
rect -34896 -30188 -34769 -30172
rect -34896 -30252 -34849 -30188
rect -34785 -30252 -34769 -30188
rect -34896 -30268 -34769 -30252
rect -34896 -30332 -34849 -30268
rect -34785 -30332 -34769 -30268
rect -34896 -30348 -34769 -30332
rect -34896 -30412 -34849 -30348
rect -34785 -30412 -34769 -30348
rect -34896 -30428 -34769 -30412
rect -34896 -30492 -34849 -30428
rect -34785 -30492 -34769 -30428
rect -34896 -30508 -34769 -30492
rect -34896 -30572 -34849 -30508
rect -34785 -30572 -34769 -30508
rect -34896 -30588 -34769 -30572
rect -34896 -30652 -34849 -30588
rect -34785 -30652 -34769 -30588
rect -34896 -30668 -34769 -30652
rect -34896 -30732 -34849 -30668
rect -34785 -30732 -34769 -30668
rect -34896 -30748 -34769 -30732
rect -34896 -30812 -34849 -30748
rect -34785 -30812 -34769 -30748
rect -34896 -30828 -34769 -30812
rect -34896 -30892 -34849 -30828
rect -34785 -30892 -34769 -30828
rect -34896 -30908 -34769 -30892
rect -34896 -30972 -34849 -30908
rect -34785 -30972 -34769 -30908
rect -34896 -30988 -34769 -30972
rect -34896 -31052 -34849 -30988
rect -34785 -31052 -34769 -30988
rect -34896 -31068 -34769 -31052
rect -34896 -31132 -34849 -31068
rect -34785 -31132 -34769 -31068
rect -34896 -31148 -34769 -31132
rect -34896 -31212 -34849 -31148
rect -34785 -31212 -34769 -31148
rect -34896 -31228 -34769 -31212
rect -34896 -31292 -34849 -31228
rect -34785 -31292 -34769 -31228
rect -34896 -31308 -34769 -31292
rect -34896 -31372 -34849 -31308
rect -34785 -31372 -34769 -31308
rect -34896 -31388 -34769 -31372
rect -34896 -31452 -34849 -31388
rect -34785 -31452 -34769 -31388
rect -34896 -31468 -34769 -31452
rect -34896 -31532 -34849 -31468
rect -34785 -31532 -34769 -31468
rect -34896 -31548 -34769 -31532
rect -34896 -31612 -34849 -31548
rect -34785 -31612 -34769 -31548
rect -34896 -31628 -34769 -31612
rect -34896 -31692 -34849 -31628
rect -34785 -31692 -34769 -31628
rect -34896 -31708 -34769 -31692
rect -34896 -31772 -34849 -31708
rect -34785 -31772 -34769 -31708
rect -34896 -31788 -34769 -31772
rect -34896 -31852 -34849 -31788
rect -34785 -31852 -34769 -31788
rect -34896 -31868 -34769 -31852
rect -34896 -31932 -34849 -31868
rect -34785 -31932 -34769 -31868
rect -34896 -31948 -34769 -31932
rect -34896 -32012 -34849 -31948
rect -34785 -32012 -34769 -31948
rect -34896 -32028 -34769 -32012
rect -34896 -32092 -34849 -32028
rect -34785 -32092 -34769 -32028
rect -34896 -32108 -34769 -32092
rect -34896 -32172 -34849 -32108
rect -34785 -32172 -34769 -32108
rect -34896 -32188 -34769 -32172
rect -34896 -32252 -34849 -32188
rect -34785 -32252 -34769 -32188
rect -34896 -32268 -34769 -32252
rect -34896 -32332 -34849 -32268
rect -34785 -32332 -34769 -32268
rect -34896 -32348 -34769 -32332
rect -34896 -32412 -34849 -32348
rect -34785 -32412 -34769 -32348
rect -34896 -32428 -34769 -32412
rect -34896 -32492 -34849 -32428
rect -34785 -32492 -34769 -32428
rect -34896 -32508 -34769 -32492
rect -34896 -32572 -34849 -32508
rect -34785 -32572 -34769 -32508
rect -34896 -32588 -34769 -32572
rect -34896 -32652 -34849 -32588
rect -34785 -32652 -34769 -32588
rect -34896 -32668 -34769 -32652
rect -34896 -32732 -34849 -32668
rect -34785 -32732 -34769 -32668
rect -34896 -32748 -34769 -32732
rect -34896 -32812 -34849 -32748
rect -34785 -32812 -34769 -32748
rect -34896 -32828 -34769 -32812
rect -34896 -32892 -34849 -32828
rect -34785 -32892 -34769 -32828
rect -34896 -32908 -34769 -32892
rect -34896 -32972 -34849 -32908
rect -34785 -32972 -34769 -32908
rect -34896 -32988 -34769 -32972
rect -34896 -33052 -34849 -32988
rect -34785 -33052 -34769 -32988
rect -34896 -33068 -34769 -33052
rect -34896 -33132 -34849 -33068
rect -34785 -33132 -34769 -33068
rect -34896 -33148 -34769 -33132
rect -34896 -33212 -34849 -33148
rect -34785 -33212 -34769 -33148
rect -34896 -33228 -34769 -33212
rect -34896 -33292 -34849 -33228
rect -34785 -33292 -34769 -33228
rect -34896 -33308 -34769 -33292
rect -34896 -33372 -34849 -33308
rect -34785 -33372 -34769 -33308
rect -34896 -33388 -34769 -33372
rect -34896 -33452 -34849 -33388
rect -34785 -33452 -34769 -33388
rect -34896 -33468 -34769 -33452
rect -34896 -33532 -34849 -33468
rect -34785 -33532 -34769 -33468
rect -34896 -33548 -34769 -33532
rect -34896 -33612 -34849 -33548
rect -34785 -33612 -34769 -33548
rect -34896 -33628 -34769 -33612
rect -34896 -33692 -34849 -33628
rect -34785 -33692 -34769 -33628
rect -34896 -33708 -34769 -33692
rect -34896 -33772 -34849 -33708
rect -34785 -33772 -34769 -33708
rect -34896 -33788 -34769 -33772
rect -34896 -33852 -34849 -33788
rect -34785 -33852 -34769 -33788
rect -34896 -33868 -34769 -33852
rect -34896 -33932 -34849 -33868
rect -34785 -33932 -34769 -33868
rect -34896 -33948 -34769 -33932
rect -34896 -34012 -34849 -33948
rect -34785 -34012 -34769 -33948
rect -34896 -34028 -34769 -34012
rect -34896 -34092 -34849 -34028
rect -34785 -34092 -34769 -34028
rect -34896 -34108 -34769 -34092
rect -34896 -34172 -34849 -34108
rect -34785 -34172 -34769 -34108
rect -34896 -34188 -34769 -34172
rect -34896 -34252 -34849 -34188
rect -34785 -34252 -34769 -34188
rect -34896 -34268 -34769 -34252
rect -34896 -34332 -34849 -34268
rect -34785 -34332 -34769 -34268
rect -34896 -34348 -34769 -34332
rect -34896 -34412 -34849 -34348
rect -34785 -34412 -34769 -34348
rect -34896 -34428 -34769 -34412
rect -41215 -34508 -41088 -34492
rect -41215 -34572 -41168 -34508
rect -41104 -34572 -41088 -34508
rect -41215 -34588 -41088 -34572
rect -41215 -34712 -41111 -34588
rect -41215 -34728 -41088 -34712
rect -41215 -34792 -41168 -34728
rect -41104 -34792 -41088 -34728
rect -41215 -34808 -41088 -34792
rect -47244 -34848 -41322 -34839
rect -47244 -40752 -47235 -34848
rect -41331 -40752 -41322 -34848
rect -47244 -40761 -41322 -40752
rect -41215 -34872 -41168 -34808
rect -41104 -34872 -41088 -34808
rect -38016 -34839 -37912 -34461
rect -34896 -34492 -34849 -34428
rect -34785 -34492 -34769 -34428
rect -34606 -28548 -28684 -28539
rect -34606 -34452 -34597 -28548
rect -28693 -34452 -28684 -28548
rect -34606 -34461 -28684 -34452
rect -28577 -28572 -28530 -28508
rect -28466 -28572 -28450 -28508
rect -25378 -28539 -25274 -28161
rect -22258 -28192 -22211 -28128
rect -22147 -28192 -22131 -28128
rect -21968 -22248 -16046 -22239
rect -21968 -28152 -21959 -22248
rect -16055 -28152 -16046 -22248
rect -21968 -28161 -16046 -28152
rect -15939 -22272 -15892 -22208
rect -15828 -22272 -15812 -22208
rect -12740 -22239 -12636 -21861
rect -9620 -21892 -9573 -21828
rect -9509 -21892 -9493 -21828
rect -9330 -15948 -3408 -15939
rect -9330 -21852 -9321 -15948
rect -3417 -21852 -3408 -15948
rect -9330 -21861 -3408 -21852
rect -3301 -15972 -3254 -15908
rect -3190 -15972 -3174 -15908
rect -102 -15939 2 -15561
rect 3018 -15592 3065 -15528
rect 3129 -15592 3145 -15528
rect 3308 -9648 9230 -9639
rect 3308 -15552 3317 -9648
rect 9221 -15552 9230 -9648
rect 3308 -15561 9230 -15552
rect 9337 -9672 9384 -9608
rect 9448 -9672 9464 -9608
rect 12536 -9639 12640 -9261
rect 15656 -9292 15703 -9228
rect 15767 -9292 15783 -9228
rect 15946 -3348 21868 -3339
rect 15946 -9252 15955 -3348
rect 21859 -9252 21868 -3348
rect 15946 -9261 21868 -9252
rect 21975 -3372 22022 -3308
rect 22086 -3372 22102 -3308
rect 25174 -3339 25278 -2961
rect 28294 -2992 28341 -2928
rect 28405 -2992 28421 -2928
rect 28584 2952 34506 2961
rect 28584 -2952 28593 2952
rect 34497 -2952 34506 2952
rect 28584 -2961 34506 -2952
rect 34613 2928 34660 2992
rect 34724 2928 34740 2992
rect 37812 2961 37916 3339
rect 40932 3308 40979 3372
rect 41043 3308 41059 3372
rect 41222 9252 47144 9261
rect 41222 3348 41231 9252
rect 47135 3348 47144 9252
rect 41222 3339 47144 3348
rect 47251 9228 47298 9292
rect 47362 9228 47378 9292
rect 47251 9212 47378 9228
rect 47251 9148 47298 9212
rect 47362 9148 47378 9212
rect 47251 9132 47378 9148
rect 47251 9068 47298 9132
rect 47362 9068 47378 9132
rect 47251 9052 47378 9068
rect 47251 8988 47298 9052
rect 47362 8988 47378 9052
rect 47251 8972 47378 8988
rect 47251 8908 47298 8972
rect 47362 8908 47378 8972
rect 47251 8892 47378 8908
rect 47251 8828 47298 8892
rect 47362 8828 47378 8892
rect 47251 8812 47378 8828
rect 47251 8748 47298 8812
rect 47362 8748 47378 8812
rect 47251 8732 47378 8748
rect 47251 8668 47298 8732
rect 47362 8668 47378 8732
rect 47251 8652 47378 8668
rect 47251 8588 47298 8652
rect 47362 8588 47378 8652
rect 47251 8572 47378 8588
rect 47251 8508 47298 8572
rect 47362 8508 47378 8572
rect 47251 8492 47378 8508
rect 47251 8428 47298 8492
rect 47362 8428 47378 8492
rect 47251 8412 47378 8428
rect 47251 8348 47298 8412
rect 47362 8348 47378 8412
rect 47251 8332 47378 8348
rect 47251 8268 47298 8332
rect 47362 8268 47378 8332
rect 47251 8252 47378 8268
rect 47251 8188 47298 8252
rect 47362 8188 47378 8252
rect 47251 8172 47378 8188
rect 47251 8108 47298 8172
rect 47362 8108 47378 8172
rect 47251 8092 47378 8108
rect 47251 8028 47298 8092
rect 47362 8028 47378 8092
rect 47251 8012 47378 8028
rect 47251 7948 47298 8012
rect 47362 7948 47378 8012
rect 47251 7932 47378 7948
rect 47251 7868 47298 7932
rect 47362 7868 47378 7932
rect 47251 7852 47378 7868
rect 47251 7788 47298 7852
rect 47362 7788 47378 7852
rect 47251 7772 47378 7788
rect 47251 7708 47298 7772
rect 47362 7708 47378 7772
rect 47251 7692 47378 7708
rect 47251 7628 47298 7692
rect 47362 7628 47378 7692
rect 47251 7612 47378 7628
rect 47251 7548 47298 7612
rect 47362 7548 47378 7612
rect 47251 7532 47378 7548
rect 47251 7468 47298 7532
rect 47362 7468 47378 7532
rect 47251 7452 47378 7468
rect 47251 7388 47298 7452
rect 47362 7388 47378 7452
rect 47251 7372 47378 7388
rect 47251 7308 47298 7372
rect 47362 7308 47378 7372
rect 47251 7292 47378 7308
rect 47251 7228 47298 7292
rect 47362 7228 47378 7292
rect 47251 7212 47378 7228
rect 47251 7148 47298 7212
rect 47362 7148 47378 7212
rect 47251 7132 47378 7148
rect 47251 7068 47298 7132
rect 47362 7068 47378 7132
rect 47251 7052 47378 7068
rect 47251 6988 47298 7052
rect 47362 6988 47378 7052
rect 47251 6972 47378 6988
rect 47251 6908 47298 6972
rect 47362 6908 47378 6972
rect 47251 6892 47378 6908
rect 47251 6828 47298 6892
rect 47362 6828 47378 6892
rect 47251 6812 47378 6828
rect 47251 6748 47298 6812
rect 47362 6748 47378 6812
rect 47251 6732 47378 6748
rect 47251 6668 47298 6732
rect 47362 6668 47378 6732
rect 47251 6652 47378 6668
rect 47251 6588 47298 6652
rect 47362 6588 47378 6652
rect 47251 6572 47378 6588
rect 47251 6508 47298 6572
rect 47362 6508 47378 6572
rect 47251 6492 47378 6508
rect 47251 6428 47298 6492
rect 47362 6428 47378 6492
rect 47251 6412 47378 6428
rect 47251 6348 47298 6412
rect 47362 6348 47378 6412
rect 47251 6332 47378 6348
rect 47251 6268 47298 6332
rect 47362 6268 47378 6332
rect 47251 6252 47378 6268
rect 47251 6188 47298 6252
rect 47362 6188 47378 6252
rect 47251 6172 47378 6188
rect 47251 6108 47298 6172
rect 47362 6108 47378 6172
rect 47251 6092 47378 6108
rect 47251 6028 47298 6092
rect 47362 6028 47378 6092
rect 47251 6012 47378 6028
rect 47251 5948 47298 6012
rect 47362 5948 47378 6012
rect 47251 5932 47378 5948
rect 47251 5868 47298 5932
rect 47362 5868 47378 5932
rect 47251 5852 47378 5868
rect 47251 5788 47298 5852
rect 47362 5788 47378 5852
rect 47251 5772 47378 5788
rect 47251 5708 47298 5772
rect 47362 5708 47378 5772
rect 47251 5692 47378 5708
rect 47251 5628 47298 5692
rect 47362 5628 47378 5692
rect 47251 5612 47378 5628
rect 47251 5548 47298 5612
rect 47362 5548 47378 5612
rect 47251 5532 47378 5548
rect 47251 5468 47298 5532
rect 47362 5468 47378 5532
rect 47251 5452 47378 5468
rect 47251 5388 47298 5452
rect 47362 5388 47378 5452
rect 47251 5372 47378 5388
rect 47251 5308 47298 5372
rect 47362 5308 47378 5372
rect 47251 5292 47378 5308
rect 47251 5228 47298 5292
rect 47362 5228 47378 5292
rect 47251 5212 47378 5228
rect 47251 5148 47298 5212
rect 47362 5148 47378 5212
rect 47251 5132 47378 5148
rect 47251 5068 47298 5132
rect 47362 5068 47378 5132
rect 47251 5052 47378 5068
rect 47251 4988 47298 5052
rect 47362 4988 47378 5052
rect 47251 4972 47378 4988
rect 47251 4908 47298 4972
rect 47362 4908 47378 4972
rect 47251 4892 47378 4908
rect 47251 4828 47298 4892
rect 47362 4828 47378 4892
rect 47251 4812 47378 4828
rect 47251 4748 47298 4812
rect 47362 4748 47378 4812
rect 47251 4732 47378 4748
rect 47251 4668 47298 4732
rect 47362 4668 47378 4732
rect 47251 4652 47378 4668
rect 47251 4588 47298 4652
rect 47362 4588 47378 4652
rect 47251 4572 47378 4588
rect 47251 4508 47298 4572
rect 47362 4508 47378 4572
rect 47251 4492 47378 4508
rect 47251 4428 47298 4492
rect 47362 4428 47378 4492
rect 47251 4412 47378 4428
rect 47251 4348 47298 4412
rect 47362 4348 47378 4412
rect 47251 4332 47378 4348
rect 47251 4268 47298 4332
rect 47362 4268 47378 4332
rect 47251 4252 47378 4268
rect 47251 4188 47298 4252
rect 47362 4188 47378 4252
rect 47251 4172 47378 4188
rect 47251 4108 47298 4172
rect 47362 4108 47378 4172
rect 47251 4092 47378 4108
rect 47251 4028 47298 4092
rect 47362 4028 47378 4092
rect 47251 4012 47378 4028
rect 47251 3948 47298 4012
rect 47362 3948 47378 4012
rect 47251 3932 47378 3948
rect 47251 3868 47298 3932
rect 47362 3868 47378 3932
rect 47251 3852 47378 3868
rect 47251 3788 47298 3852
rect 47362 3788 47378 3852
rect 47251 3772 47378 3788
rect 47251 3708 47298 3772
rect 47362 3708 47378 3772
rect 47251 3692 47378 3708
rect 47251 3628 47298 3692
rect 47362 3628 47378 3692
rect 47251 3612 47378 3628
rect 47251 3548 47298 3612
rect 47362 3548 47378 3612
rect 47251 3532 47378 3548
rect 47251 3468 47298 3532
rect 47362 3468 47378 3532
rect 47251 3452 47378 3468
rect 47251 3388 47298 3452
rect 47362 3388 47378 3452
rect 47251 3372 47378 3388
rect 40932 3292 41059 3308
rect 40932 3228 40979 3292
rect 41043 3228 41059 3292
rect 40932 3212 41059 3228
rect 40932 3088 41036 3212
rect 40932 3072 41059 3088
rect 40932 3008 40979 3072
rect 41043 3008 41059 3072
rect 40932 2992 41059 3008
rect 34613 2912 34740 2928
rect 34613 2848 34660 2912
rect 34724 2848 34740 2912
rect 34613 2832 34740 2848
rect 34613 2768 34660 2832
rect 34724 2768 34740 2832
rect 34613 2752 34740 2768
rect 34613 2688 34660 2752
rect 34724 2688 34740 2752
rect 34613 2672 34740 2688
rect 34613 2608 34660 2672
rect 34724 2608 34740 2672
rect 34613 2592 34740 2608
rect 34613 2528 34660 2592
rect 34724 2528 34740 2592
rect 34613 2512 34740 2528
rect 34613 2448 34660 2512
rect 34724 2448 34740 2512
rect 34613 2432 34740 2448
rect 34613 2368 34660 2432
rect 34724 2368 34740 2432
rect 34613 2352 34740 2368
rect 34613 2288 34660 2352
rect 34724 2288 34740 2352
rect 34613 2272 34740 2288
rect 34613 2208 34660 2272
rect 34724 2208 34740 2272
rect 34613 2192 34740 2208
rect 34613 2128 34660 2192
rect 34724 2128 34740 2192
rect 34613 2112 34740 2128
rect 34613 2048 34660 2112
rect 34724 2048 34740 2112
rect 34613 2032 34740 2048
rect 34613 1968 34660 2032
rect 34724 1968 34740 2032
rect 34613 1952 34740 1968
rect 34613 1888 34660 1952
rect 34724 1888 34740 1952
rect 34613 1872 34740 1888
rect 34613 1808 34660 1872
rect 34724 1808 34740 1872
rect 34613 1792 34740 1808
rect 34613 1728 34660 1792
rect 34724 1728 34740 1792
rect 34613 1712 34740 1728
rect 34613 1648 34660 1712
rect 34724 1648 34740 1712
rect 34613 1632 34740 1648
rect 34613 1568 34660 1632
rect 34724 1568 34740 1632
rect 34613 1552 34740 1568
rect 34613 1488 34660 1552
rect 34724 1488 34740 1552
rect 34613 1472 34740 1488
rect 34613 1408 34660 1472
rect 34724 1408 34740 1472
rect 34613 1392 34740 1408
rect 34613 1328 34660 1392
rect 34724 1328 34740 1392
rect 34613 1312 34740 1328
rect 34613 1248 34660 1312
rect 34724 1248 34740 1312
rect 34613 1232 34740 1248
rect 34613 1168 34660 1232
rect 34724 1168 34740 1232
rect 34613 1152 34740 1168
rect 34613 1088 34660 1152
rect 34724 1088 34740 1152
rect 34613 1072 34740 1088
rect 34613 1008 34660 1072
rect 34724 1008 34740 1072
rect 34613 992 34740 1008
rect 34613 928 34660 992
rect 34724 928 34740 992
rect 34613 912 34740 928
rect 34613 848 34660 912
rect 34724 848 34740 912
rect 34613 832 34740 848
rect 34613 768 34660 832
rect 34724 768 34740 832
rect 34613 752 34740 768
rect 34613 688 34660 752
rect 34724 688 34740 752
rect 34613 672 34740 688
rect 34613 608 34660 672
rect 34724 608 34740 672
rect 34613 592 34740 608
rect 34613 528 34660 592
rect 34724 528 34740 592
rect 34613 512 34740 528
rect 34613 448 34660 512
rect 34724 448 34740 512
rect 34613 432 34740 448
rect 34613 368 34660 432
rect 34724 368 34740 432
rect 34613 352 34740 368
rect 34613 288 34660 352
rect 34724 288 34740 352
rect 34613 272 34740 288
rect 34613 208 34660 272
rect 34724 208 34740 272
rect 34613 192 34740 208
rect 34613 128 34660 192
rect 34724 128 34740 192
rect 34613 112 34740 128
rect 34613 48 34660 112
rect 34724 48 34740 112
rect 34613 32 34740 48
rect 34613 -32 34660 32
rect 34724 -32 34740 32
rect 34613 -48 34740 -32
rect 34613 -112 34660 -48
rect 34724 -112 34740 -48
rect 34613 -128 34740 -112
rect 34613 -192 34660 -128
rect 34724 -192 34740 -128
rect 34613 -208 34740 -192
rect 34613 -272 34660 -208
rect 34724 -272 34740 -208
rect 34613 -288 34740 -272
rect 34613 -352 34660 -288
rect 34724 -352 34740 -288
rect 34613 -368 34740 -352
rect 34613 -432 34660 -368
rect 34724 -432 34740 -368
rect 34613 -448 34740 -432
rect 34613 -512 34660 -448
rect 34724 -512 34740 -448
rect 34613 -528 34740 -512
rect 34613 -592 34660 -528
rect 34724 -592 34740 -528
rect 34613 -608 34740 -592
rect 34613 -672 34660 -608
rect 34724 -672 34740 -608
rect 34613 -688 34740 -672
rect 34613 -752 34660 -688
rect 34724 -752 34740 -688
rect 34613 -768 34740 -752
rect 34613 -832 34660 -768
rect 34724 -832 34740 -768
rect 34613 -848 34740 -832
rect 34613 -912 34660 -848
rect 34724 -912 34740 -848
rect 34613 -928 34740 -912
rect 34613 -992 34660 -928
rect 34724 -992 34740 -928
rect 34613 -1008 34740 -992
rect 34613 -1072 34660 -1008
rect 34724 -1072 34740 -1008
rect 34613 -1088 34740 -1072
rect 34613 -1152 34660 -1088
rect 34724 -1152 34740 -1088
rect 34613 -1168 34740 -1152
rect 34613 -1232 34660 -1168
rect 34724 -1232 34740 -1168
rect 34613 -1248 34740 -1232
rect 34613 -1312 34660 -1248
rect 34724 -1312 34740 -1248
rect 34613 -1328 34740 -1312
rect 34613 -1392 34660 -1328
rect 34724 -1392 34740 -1328
rect 34613 -1408 34740 -1392
rect 34613 -1472 34660 -1408
rect 34724 -1472 34740 -1408
rect 34613 -1488 34740 -1472
rect 34613 -1552 34660 -1488
rect 34724 -1552 34740 -1488
rect 34613 -1568 34740 -1552
rect 34613 -1632 34660 -1568
rect 34724 -1632 34740 -1568
rect 34613 -1648 34740 -1632
rect 34613 -1712 34660 -1648
rect 34724 -1712 34740 -1648
rect 34613 -1728 34740 -1712
rect 34613 -1792 34660 -1728
rect 34724 -1792 34740 -1728
rect 34613 -1808 34740 -1792
rect 34613 -1872 34660 -1808
rect 34724 -1872 34740 -1808
rect 34613 -1888 34740 -1872
rect 34613 -1952 34660 -1888
rect 34724 -1952 34740 -1888
rect 34613 -1968 34740 -1952
rect 34613 -2032 34660 -1968
rect 34724 -2032 34740 -1968
rect 34613 -2048 34740 -2032
rect 34613 -2112 34660 -2048
rect 34724 -2112 34740 -2048
rect 34613 -2128 34740 -2112
rect 34613 -2192 34660 -2128
rect 34724 -2192 34740 -2128
rect 34613 -2208 34740 -2192
rect 34613 -2272 34660 -2208
rect 34724 -2272 34740 -2208
rect 34613 -2288 34740 -2272
rect 34613 -2352 34660 -2288
rect 34724 -2352 34740 -2288
rect 34613 -2368 34740 -2352
rect 34613 -2432 34660 -2368
rect 34724 -2432 34740 -2368
rect 34613 -2448 34740 -2432
rect 34613 -2512 34660 -2448
rect 34724 -2512 34740 -2448
rect 34613 -2528 34740 -2512
rect 34613 -2592 34660 -2528
rect 34724 -2592 34740 -2528
rect 34613 -2608 34740 -2592
rect 34613 -2672 34660 -2608
rect 34724 -2672 34740 -2608
rect 34613 -2688 34740 -2672
rect 34613 -2752 34660 -2688
rect 34724 -2752 34740 -2688
rect 34613 -2768 34740 -2752
rect 34613 -2832 34660 -2768
rect 34724 -2832 34740 -2768
rect 34613 -2848 34740 -2832
rect 34613 -2912 34660 -2848
rect 34724 -2912 34740 -2848
rect 34613 -2928 34740 -2912
rect 28294 -3008 28421 -2992
rect 28294 -3072 28341 -3008
rect 28405 -3072 28421 -3008
rect 28294 -3088 28421 -3072
rect 28294 -3212 28398 -3088
rect 28294 -3228 28421 -3212
rect 28294 -3292 28341 -3228
rect 28405 -3292 28421 -3228
rect 28294 -3308 28421 -3292
rect 21975 -3388 22102 -3372
rect 21975 -3452 22022 -3388
rect 22086 -3452 22102 -3388
rect 21975 -3468 22102 -3452
rect 21975 -3532 22022 -3468
rect 22086 -3532 22102 -3468
rect 21975 -3548 22102 -3532
rect 21975 -3612 22022 -3548
rect 22086 -3612 22102 -3548
rect 21975 -3628 22102 -3612
rect 21975 -3692 22022 -3628
rect 22086 -3692 22102 -3628
rect 21975 -3708 22102 -3692
rect 21975 -3772 22022 -3708
rect 22086 -3772 22102 -3708
rect 21975 -3788 22102 -3772
rect 21975 -3852 22022 -3788
rect 22086 -3852 22102 -3788
rect 21975 -3868 22102 -3852
rect 21975 -3932 22022 -3868
rect 22086 -3932 22102 -3868
rect 21975 -3948 22102 -3932
rect 21975 -4012 22022 -3948
rect 22086 -4012 22102 -3948
rect 21975 -4028 22102 -4012
rect 21975 -4092 22022 -4028
rect 22086 -4092 22102 -4028
rect 21975 -4108 22102 -4092
rect 21975 -4172 22022 -4108
rect 22086 -4172 22102 -4108
rect 21975 -4188 22102 -4172
rect 21975 -4252 22022 -4188
rect 22086 -4252 22102 -4188
rect 21975 -4268 22102 -4252
rect 21975 -4332 22022 -4268
rect 22086 -4332 22102 -4268
rect 21975 -4348 22102 -4332
rect 21975 -4412 22022 -4348
rect 22086 -4412 22102 -4348
rect 21975 -4428 22102 -4412
rect 21975 -4492 22022 -4428
rect 22086 -4492 22102 -4428
rect 21975 -4508 22102 -4492
rect 21975 -4572 22022 -4508
rect 22086 -4572 22102 -4508
rect 21975 -4588 22102 -4572
rect 21975 -4652 22022 -4588
rect 22086 -4652 22102 -4588
rect 21975 -4668 22102 -4652
rect 21975 -4732 22022 -4668
rect 22086 -4732 22102 -4668
rect 21975 -4748 22102 -4732
rect 21975 -4812 22022 -4748
rect 22086 -4812 22102 -4748
rect 21975 -4828 22102 -4812
rect 21975 -4892 22022 -4828
rect 22086 -4892 22102 -4828
rect 21975 -4908 22102 -4892
rect 21975 -4972 22022 -4908
rect 22086 -4972 22102 -4908
rect 21975 -4988 22102 -4972
rect 21975 -5052 22022 -4988
rect 22086 -5052 22102 -4988
rect 21975 -5068 22102 -5052
rect 21975 -5132 22022 -5068
rect 22086 -5132 22102 -5068
rect 21975 -5148 22102 -5132
rect 21975 -5212 22022 -5148
rect 22086 -5212 22102 -5148
rect 21975 -5228 22102 -5212
rect 21975 -5292 22022 -5228
rect 22086 -5292 22102 -5228
rect 21975 -5308 22102 -5292
rect 21975 -5372 22022 -5308
rect 22086 -5372 22102 -5308
rect 21975 -5388 22102 -5372
rect 21975 -5452 22022 -5388
rect 22086 -5452 22102 -5388
rect 21975 -5468 22102 -5452
rect 21975 -5532 22022 -5468
rect 22086 -5532 22102 -5468
rect 21975 -5548 22102 -5532
rect 21975 -5612 22022 -5548
rect 22086 -5612 22102 -5548
rect 21975 -5628 22102 -5612
rect 21975 -5692 22022 -5628
rect 22086 -5692 22102 -5628
rect 21975 -5708 22102 -5692
rect 21975 -5772 22022 -5708
rect 22086 -5772 22102 -5708
rect 21975 -5788 22102 -5772
rect 21975 -5852 22022 -5788
rect 22086 -5852 22102 -5788
rect 21975 -5868 22102 -5852
rect 21975 -5932 22022 -5868
rect 22086 -5932 22102 -5868
rect 21975 -5948 22102 -5932
rect 21975 -6012 22022 -5948
rect 22086 -6012 22102 -5948
rect 21975 -6028 22102 -6012
rect 21975 -6092 22022 -6028
rect 22086 -6092 22102 -6028
rect 21975 -6108 22102 -6092
rect 21975 -6172 22022 -6108
rect 22086 -6172 22102 -6108
rect 21975 -6188 22102 -6172
rect 21975 -6252 22022 -6188
rect 22086 -6252 22102 -6188
rect 21975 -6268 22102 -6252
rect 21975 -6332 22022 -6268
rect 22086 -6332 22102 -6268
rect 21975 -6348 22102 -6332
rect 21975 -6412 22022 -6348
rect 22086 -6412 22102 -6348
rect 21975 -6428 22102 -6412
rect 21975 -6492 22022 -6428
rect 22086 -6492 22102 -6428
rect 21975 -6508 22102 -6492
rect 21975 -6572 22022 -6508
rect 22086 -6572 22102 -6508
rect 21975 -6588 22102 -6572
rect 21975 -6652 22022 -6588
rect 22086 -6652 22102 -6588
rect 21975 -6668 22102 -6652
rect 21975 -6732 22022 -6668
rect 22086 -6732 22102 -6668
rect 21975 -6748 22102 -6732
rect 21975 -6812 22022 -6748
rect 22086 -6812 22102 -6748
rect 21975 -6828 22102 -6812
rect 21975 -6892 22022 -6828
rect 22086 -6892 22102 -6828
rect 21975 -6908 22102 -6892
rect 21975 -6972 22022 -6908
rect 22086 -6972 22102 -6908
rect 21975 -6988 22102 -6972
rect 21975 -7052 22022 -6988
rect 22086 -7052 22102 -6988
rect 21975 -7068 22102 -7052
rect 21975 -7132 22022 -7068
rect 22086 -7132 22102 -7068
rect 21975 -7148 22102 -7132
rect 21975 -7212 22022 -7148
rect 22086 -7212 22102 -7148
rect 21975 -7228 22102 -7212
rect 21975 -7292 22022 -7228
rect 22086 -7292 22102 -7228
rect 21975 -7308 22102 -7292
rect 21975 -7372 22022 -7308
rect 22086 -7372 22102 -7308
rect 21975 -7388 22102 -7372
rect 21975 -7452 22022 -7388
rect 22086 -7452 22102 -7388
rect 21975 -7468 22102 -7452
rect 21975 -7532 22022 -7468
rect 22086 -7532 22102 -7468
rect 21975 -7548 22102 -7532
rect 21975 -7612 22022 -7548
rect 22086 -7612 22102 -7548
rect 21975 -7628 22102 -7612
rect 21975 -7692 22022 -7628
rect 22086 -7692 22102 -7628
rect 21975 -7708 22102 -7692
rect 21975 -7772 22022 -7708
rect 22086 -7772 22102 -7708
rect 21975 -7788 22102 -7772
rect 21975 -7852 22022 -7788
rect 22086 -7852 22102 -7788
rect 21975 -7868 22102 -7852
rect 21975 -7932 22022 -7868
rect 22086 -7932 22102 -7868
rect 21975 -7948 22102 -7932
rect 21975 -8012 22022 -7948
rect 22086 -8012 22102 -7948
rect 21975 -8028 22102 -8012
rect 21975 -8092 22022 -8028
rect 22086 -8092 22102 -8028
rect 21975 -8108 22102 -8092
rect 21975 -8172 22022 -8108
rect 22086 -8172 22102 -8108
rect 21975 -8188 22102 -8172
rect 21975 -8252 22022 -8188
rect 22086 -8252 22102 -8188
rect 21975 -8268 22102 -8252
rect 21975 -8332 22022 -8268
rect 22086 -8332 22102 -8268
rect 21975 -8348 22102 -8332
rect 21975 -8412 22022 -8348
rect 22086 -8412 22102 -8348
rect 21975 -8428 22102 -8412
rect 21975 -8492 22022 -8428
rect 22086 -8492 22102 -8428
rect 21975 -8508 22102 -8492
rect 21975 -8572 22022 -8508
rect 22086 -8572 22102 -8508
rect 21975 -8588 22102 -8572
rect 21975 -8652 22022 -8588
rect 22086 -8652 22102 -8588
rect 21975 -8668 22102 -8652
rect 21975 -8732 22022 -8668
rect 22086 -8732 22102 -8668
rect 21975 -8748 22102 -8732
rect 21975 -8812 22022 -8748
rect 22086 -8812 22102 -8748
rect 21975 -8828 22102 -8812
rect 21975 -8892 22022 -8828
rect 22086 -8892 22102 -8828
rect 21975 -8908 22102 -8892
rect 21975 -8972 22022 -8908
rect 22086 -8972 22102 -8908
rect 21975 -8988 22102 -8972
rect 21975 -9052 22022 -8988
rect 22086 -9052 22102 -8988
rect 21975 -9068 22102 -9052
rect 21975 -9132 22022 -9068
rect 22086 -9132 22102 -9068
rect 21975 -9148 22102 -9132
rect 21975 -9212 22022 -9148
rect 22086 -9212 22102 -9148
rect 21975 -9228 22102 -9212
rect 15656 -9308 15783 -9292
rect 15656 -9372 15703 -9308
rect 15767 -9372 15783 -9308
rect 15656 -9388 15783 -9372
rect 15656 -9512 15760 -9388
rect 15656 -9528 15783 -9512
rect 15656 -9592 15703 -9528
rect 15767 -9592 15783 -9528
rect 15656 -9608 15783 -9592
rect 9337 -9688 9464 -9672
rect 9337 -9752 9384 -9688
rect 9448 -9752 9464 -9688
rect 9337 -9768 9464 -9752
rect 9337 -9832 9384 -9768
rect 9448 -9832 9464 -9768
rect 9337 -9848 9464 -9832
rect 9337 -9912 9384 -9848
rect 9448 -9912 9464 -9848
rect 9337 -9928 9464 -9912
rect 9337 -9992 9384 -9928
rect 9448 -9992 9464 -9928
rect 9337 -10008 9464 -9992
rect 9337 -10072 9384 -10008
rect 9448 -10072 9464 -10008
rect 9337 -10088 9464 -10072
rect 9337 -10152 9384 -10088
rect 9448 -10152 9464 -10088
rect 9337 -10168 9464 -10152
rect 9337 -10232 9384 -10168
rect 9448 -10232 9464 -10168
rect 9337 -10248 9464 -10232
rect 9337 -10312 9384 -10248
rect 9448 -10312 9464 -10248
rect 9337 -10328 9464 -10312
rect 9337 -10392 9384 -10328
rect 9448 -10392 9464 -10328
rect 9337 -10408 9464 -10392
rect 9337 -10472 9384 -10408
rect 9448 -10472 9464 -10408
rect 9337 -10488 9464 -10472
rect 9337 -10552 9384 -10488
rect 9448 -10552 9464 -10488
rect 9337 -10568 9464 -10552
rect 9337 -10632 9384 -10568
rect 9448 -10632 9464 -10568
rect 9337 -10648 9464 -10632
rect 9337 -10712 9384 -10648
rect 9448 -10712 9464 -10648
rect 9337 -10728 9464 -10712
rect 9337 -10792 9384 -10728
rect 9448 -10792 9464 -10728
rect 9337 -10808 9464 -10792
rect 9337 -10872 9384 -10808
rect 9448 -10872 9464 -10808
rect 9337 -10888 9464 -10872
rect 9337 -10952 9384 -10888
rect 9448 -10952 9464 -10888
rect 9337 -10968 9464 -10952
rect 9337 -11032 9384 -10968
rect 9448 -11032 9464 -10968
rect 9337 -11048 9464 -11032
rect 9337 -11112 9384 -11048
rect 9448 -11112 9464 -11048
rect 9337 -11128 9464 -11112
rect 9337 -11192 9384 -11128
rect 9448 -11192 9464 -11128
rect 9337 -11208 9464 -11192
rect 9337 -11272 9384 -11208
rect 9448 -11272 9464 -11208
rect 9337 -11288 9464 -11272
rect 9337 -11352 9384 -11288
rect 9448 -11352 9464 -11288
rect 9337 -11368 9464 -11352
rect 9337 -11432 9384 -11368
rect 9448 -11432 9464 -11368
rect 9337 -11448 9464 -11432
rect 9337 -11512 9384 -11448
rect 9448 -11512 9464 -11448
rect 9337 -11528 9464 -11512
rect 9337 -11592 9384 -11528
rect 9448 -11592 9464 -11528
rect 9337 -11608 9464 -11592
rect 9337 -11672 9384 -11608
rect 9448 -11672 9464 -11608
rect 9337 -11688 9464 -11672
rect 9337 -11752 9384 -11688
rect 9448 -11752 9464 -11688
rect 9337 -11768 9464 -11752
rect 9337 -11832 9384 -11768
rect 9448 -11832 9464 -11768
rect 9337 -11848 9464 -11832
rect 9337 -11912 9384 -11848
rect 9448 -11912 9464 -11848
rect 9337 -11928 9464 -11912
rect 9337 -11992 9384 -11928
rect 9448 -11992 9464 -11928
rect 9337 -12008 9464 -11992
rect 9337 -12072 9384 -12008
rect 9448 -12072 9464 -12008
rect 9337 -12088 9464 -12072
rect 9337 -12152 9384 -12088
rect 9448 -12152 9464 -12088
rect 9337 -12168 9464 -12152
rect 9337 -12232 9384 -12168
rect 9448 -12232 9464 -12168
rect 9337 -12248 9464 -12232
rect 9337 -12312 9384 -12248
rect 9448 -12312 9464 -12248
rect 9337 -12328 9464 -12312
rect 9337 -12392 9384 -12328
rect 9448 -12392 9464 -12328
rect 9337 -12408 9464 -12392
rect 9337 -12472 9384 -12408
rect 9448 -12472 9464 -12408
rect 9337 -12488 9464 -12472
rect 9337 -12552 9384 -12488
rect 9448 -12552 9464 -12488
rect 9337 -12568 9464 -12552
rect 9337 -12632 9384 -12568
rect 9448 -12632 9464 -12568
rect 9337 -12648 9464 -12632
rect 9337 -12712 9384 -12648
rect 9448 -12712 9464 -12648
rect 9337 -12728 9464 -12712
rect 9337 -12792 9384 -12728
rect 9448 -12792 9464 -12728
rect 9337 -12808 9464 -12792
rect 9337 -12872 9384 -12808
rect 9448 -12872 9464 -12808
rect 9337 -12888 9464 -12872
rect 9337 -12952 9384 -12888
rect 9448 -12952 9464 -12888
rect 9337 -12968 9464 -12952
rect 9337 -13032 9384 -12968
rect 9448 -13032 9464 -12968
rect 9337 -13048 9464 -13032
rect 9337 -13112 9384 -13048
rect 9448 -13112 9464 -13048
rect 9337 -13128 9464 -13112
rect 9337 -13192 9384 -13128
rect 9448 -13192 9464 -13128
rect 9337 -13208 9464 -13192
rect 9337 -13272 9384 -13208
rect 9448 -13272 9464 -13208
rect 9337 -13288 9464 -13272
rect 9337 -13352 9384 -13288
rect 9448 -13352 9464 -13288
rect 9337 -13368 9464 -13352
rect 9337 -13432 9384 -13368
rect 9448 -13432 9464 -13368
rect 9337 -13448 9464 -13432
rect 9337 -13512 9384 -13448
rect 9448 -13512 9464 -13448
rect 9337 -13528 9464 -13512
rect 9337 -13592 9384 -13528
rect 9448 -13592 9464 -13528
rect 9337 -13608 9464 -13592
rect 9337 -13672 9384 -13608
rect 9448 -13672 9464 -13608
rect 9337 -13688 9464 -13672
rect 9337 -13752 9384 -13688
rect 9448 -13752 9464 -13688
rect 9337 -13768 9464 -13752
rect 9337 -13832 9384 -13768
rect 9448 -13832 9464 -13768
rect 9337 -13848 9464 -13832
rect 9337 -13912 9384 -13848
rect 9448 -13912 9464 -13848
rect 9337 -13928 9464 -13912
rect 9337 -13992 9384 -13928
rect 9448 -13992 9464 -13928
rect 9337 -14008 9464 -13992
rect 9337 -14072 9384 -14008
rect 9448 -14072 9464 -14008
rect 9337 -14088 9464 -14072
rect 9337 -14152 9384 -14088
rect 9448 -14152 9464 -14088
rect 9337 -14168 9464 -14152
rect 9337 -14232 9384 -14168
rect 9448 -14232 9464 -14168
rect 9337 -14248 9464 -14232
rect 9337 -14312 9384 -14248
rect 9448 -14312 9464 -14248
rect 9337 -14328 9464 -14312
rect 9337 -14392 9384 -14328
rect 9448 -14392 9464 -14328
rect 9337 -14408 9464 -14392
rect 9337 -14472 9384 -14408
rect 9448 -14472 9464 -14408
rect 9337 -14488 9464 -14472
rect 9337 -14552 9384 -14488
rect 9448 -14552 9464 -14488
rect 9337 -14568 9464 -14552
rect 9337 -14632 9384 -14568
rect 9448 -14632 9464 -14568
rect 9337 -14648 9464 -14632
rect 9337 -14712 9384 -14648
rect 9448 -14712 9464 -14648
rect 9337 -14728 9464 -14712
rect 9337 -14792 9384 -14728
rect 9448 -14792 9464 -14728
rect 9337 -14808 9464 -14792
rect 9337 -14872 9384 -14808
rect 9448 -14872 9464 -14808
rect 9337 -14888 9464 -14872
rect 9337 -14952 9384 -14888
rect 9448 -14952 9464 -14888
rect 9337 -14968 9464 -14952
rect 9337 -15032 9384 -14968
rect 9448 -15032 9464 -14968
rect 9337 -15048 9464 -15032
rect 9337 -15112 9384 -15048
rect 9448 -15112 9464 -15048
rect 9337 -15128 9464 -15112
rect 9337 -15192 9384 -15128
rect 9448 -15192 9464 -15128
rect 9337 -15208 9464 -15192
rect 9337 -15272 9384 -15208
rect 9448 -15272 9464 -15208
rect 9337 -15288 9464 -15272
rect 9337 -15352 9384 -15288
rect 9448 -15352 9464 -15288
rect 9337 -15368 9464 -15352
rect 9337 -15432 9384 -15368
rect 9448 -15432 9464 -15368
rect 9337 -15448 9464 -15432
rect 9337 -15512 9384 -15448
rect 9448 -15512 9464 -15448
rect 9337 -15528 9464 -15512
rect 3018 -15608 3145 -15592
rect 3018 -15672 3065 -15608
rect 3129 -15672 3145 -15608
rect 3018 -15688 3145 -15672
rect 3018 -15812 3122 -15688
rect 3018 -15828 3145 -15812
rect 3018 -15892 3065 -15828
rect 3129 -15892 3145 -15828
rect 3018 -15908 3145 -15892
rect -3301 -15988 -3174 -15972
rect -3301 -16052 -3254 -15988
rect -3190 -16052 -3174 -15988
rect -3301 -16068 -3174 -16052
rect -3301 -16132 -3254 -16068
rect -3190 -16132 -3174 -16068
rect -3301 -16148 -3174 -16132
rect -3301 -16212 -3254 -16148
rect -3190 -16212 -3174 -16148
rect -3301 -16228 -3174 -16212
rect -3301 -16292 -3254 -16228
rect -3190 -16292 -3174 -16228
rect -3301 -16308 -3174 -16292
rect -3301 -16372 -3254 -16308
rect -3190 -16372 -3174 -16308
rect -3301 -16388 -3174 -16372
rect -3301 -16452 -3254 -16388
rect -3190 -16452 -3174 -16388
rect -3301 -16468 -3174 -16452
rect -3301 -16532 -3254 -16468
rect -3190 -16532 -3174 -16468
rect -3301 -16548 -3174 -16532
rect -3301 -16612 -3254 -16548
rect -3190 -16612 -3174 -16548
rect -3301 -16628 -3174 -16612
rect -3301 -16692 -3254 -16628
rect -3190 -16692 -3174 -16628
rect -3301 -16708 -3174 -16692
rect -3301 -16772 -3254 -16708
rect -3190 -16772 -3174 -16708
rect -3301 -16788 -3174 -16772
rect -3301 -16852 -3254 -16788
rect -3190 -16852 -3174 -16788
rect -3301 -16868 -3174 -16852
rect -3301 -16932 -3254 -16868
rect -3190 -16932 -3174 -16868
rect -3301 -16948 -3174 -16932
rect -3301 -17012 -3254 -16948
rect -3190 -17012 -3174 -16948
rect -3301 -17028 -3174 -17012
rect -3301 -17092 -3254 -17028
rect -3190 -17092 -3174 -17028
rect -3301 -17108 -3174 -17092
rect -3301 -17172 -3254 -17108
rect -3190 -17172 -3174 -17108
rect -3301 -17188 -3174 -17172
rect -3301 -17252 -3254 -17188
rect -3190 -17252 -3174 -17188
rect -3301 -17268 -3174 -17252
rect -3301 -17332 -3254 -17268
rect -3190 -17332 -3174 -17268
rect -3301 -17348 -3174 -17332
rect -3301 -17412 -3254 -17348
rect -3190 -17412 -3174 -17348
rect -3301 -17428 -3174 -17412
rect -3301 -17492 -3254 -17428
rect -3190 -17492 -3174 -17428
rect -3301 -17508 -3174 -17492
rect -3301 -17572 -3254 -17508
rect -3190 -17572 -3174 -17508
rect -3301 -17588 -3174 -17572
rect -3301 -17652 -3254 -17588
rect -3190 -17652 -3174 -17588
rect -3301 -17668 -3174 -17652
rect -3301 -17732 -3254 -17668
rect -3190 -17732 -3174 -17668
rect -3301 -17748 -3174 -17732
rect -3301 -17812 -3254 -17748
rect -3190 -17812 -3174 -17748
rect -3301 -17828 -3174 -17812
rect -3301 -17892 -3254 -17828
rect -3190 -17892 -3174 -17828
rect -3301 -17908 -3174 -17892
rect -3301 -17972 -3254 -17908
rect -3190 -17972 -3174 -17908
rect -3301 -17988 -3174 -17972
rect -3301 -18052 -3254 -17988
rect -3190 -18052 -3174 -17988
rect -3301 -18068 -3174 -18052
rect -3301 -18132 -3254 -18068
rect -3190 -18132 -3174 -18068
rect -3301 -18148 -3174 -18132
rect -3301 -18212 -3254 -18148
rect -3190 -18212 -3174 -18148
rect -3301 -18228 -3174 -18212
rect -3301 -18292 -3254 -18228
rect -3190 -18292 -3174 -18228
rect -3301 -18308 -3174 -18292
rect -3301 -18372 -3254 -18308
rect -3190 -18372 -3174 -18308
rect -3301 -18388 -3174 -18372
rect -3301 -18452 -3254 -18388
rect -3190 -18452 -3174 -18388
rect -3301 -18468 -3174 -18452
rect -3301 -18532 -3254 -18468
rect -3190 -18532 -3174 -18468
rect -3301 -18548 -3174 -18532
rect -3301 -18612 -3254 -18548
rect -3190 -18612 -3174 -18548
rect -3301 -18628 -3174 -18612
rect -3301 -18692 -3254 -18628
rect -3190 -18692 -3174 -18628
rect -3301 -18708 -3174 -18692
rect -3301 -18772 -3254 -18708
rect -3190 -18772 -3174 -18708
rect -3301 -18788 -3174 -18772
rect -3301 -18852 -3254 -18788
rect -3190 -18852 -3174 -18788
rect -3301 -18868 -3174 -18852
rect -3301 -18932 -3254 -18868
rect -3190 -18932 -3174 -18868
rect -3301 -18948 -3174 -18932
rect -3301 -19012 -3254 -18948
rect -3190 -19012 -3174 -18948
rect -3301 -19028 -3174 -19012
rect -3301 -19092 -3254 -19028
rect -3190 -19092 -3174 -19028
rect -3301 -19108 -3174 -19092
rect -3301 -19172 -3254 -19108
rect -3190 -19172 -3174 -19108
rect -3301 -19188 -3174 -19172
rect -3301 -19252 -3254 -19188
rect -3190 -19252 -3174 -19188
rect -3301 -19268 -3174 -19252
rect -3301 -19332 -3254 -19268
rect -3190 -19332 -3174 -19268
rect -3301 -19348 -3174 -19332
rect -3301 -19412 -3254 -19348
rect -3190 -19412 -3174 -19348
rect -3301 -19428 -3174 -19412
rect -3301 -19492 -3254 -19428
rect -3190 -19492 -3174 -19428
rect -3301 -19508 -3174 -19492
rect -3301 -19572 -3254 -19508
rect -3190 -19572 -3174 -19508
rect -3301 -19588 -3174 -19572
rect -3301 -19652 -3254 -19588
rect -3190 -19652 -3174 -19588
rect -3301 -19668 -3174 -19652
rect -3301 -19732 -3254 -19668
rect -3190 -19732 -3174 -19668
rect -3301 -19748 -3174 -19732
rect -3301 -19812 -3254 -19748
rect -3190 -19812 -3174 -19748
rect -3301 -19828 -3174 -19812
rect -3301 -19892 -3254 -19828
rect -3190 -19892 -3174 -19828
rect -3301 -19908 -3174 -19892
rect -3301 -19972 -3254 -19908
rect -3190 -19972 -3174 -19908
rect -3301 -19988 -3174 -19972
rect -3301 -20052 -3254 -19988
rect -3190 -20052 -3174 -19988
rect -3301 -20068 -3174 -20052
rect -3301 -20132 -3254 -20068
rect -3190 -20132 -3174 -20068
rect -3301 -20148 -3174 -20132
rect -3301 -20212 -3254 -20148
rect -3190 -20212 -3174 -20148
rect -3301 -20228 -3174 -20212
rect -3301 -20292 -3254 -20228
rect -3190 -20292 -3174 -20228
rect -3301 -20308 -3174 -20292
rect -3301 -20372 -3254 -20308
rect -3190 -20372 -3174 -20308
rect -3301 -20388 -3174 -20372
rect -3301 -20452 -3254 -20388
rect -3190 -20452 -3174 -20388
rect -3301 -20468 -3174 -20452
rect -3301 -20532 -3254 -20468
rect -3190 -20532 -3174 -20468
rect -3301 -20548 -3174 -20532
rect -3301 -20612 -3254 -20548
rect -3190 -20612 -3174 -20548
rect -3301 -20628 -3174 -20612
rect -3301 -20692 -3254 -20628
rect -3190 -20692 -3174 -20628
rect -3301 -20708 -3174 -20692
rect -3301 -20772 -3254 -20708
rect -3190 -20772 -3174 -20708
rect -3301 -20788 -3174 -20772
rect -3301 -20852 -3254 -20788
rect -3190 -20852 -3174 -20788
rect -3301 -20868 -3174 -20852
rect -3301 -20932 -3254 -20868
rect -3190 -20932 -3174 -20868
rect -3301 -20948 -3174 -20932
rect -3301 -21012 -3254 -20948
rect -3190 -21012 -3174 -20948
rect -3301 -21028 -3174 -21012
rect -3301 -21092 -3254 -21028
rect -3190 -21092 -3174 -21028
rect -3301 -21108 -3174 -21092
rect -3301 -21172 -3254 -21108
rect -3190 -21172 -3174 -21108
rect -3301 -21188 -3174 -21172
rect -3301 -21252 -3254 -21188
rect -3190 -21252 -3174 -21188
rect -3301 -21268 -3174 -21252
rect -3301 -21332 -3254 -21268
rect -3190 -21332 -3174 -21268
rect -3301 -21348 -3174 -21332
rect -3301 -21412 -3254 -21348
rect -3190 -21412 -3174 -21348
rect -3301 -21428 -3174 -21412
rect -3301 -21492 -3254 -21428
rect -3190 -21492 -3174 -21428
rect -3301 -21508 -3174 -21492
rect -3301 -21572 -3254 -21508
rect -3190 -21572 -3174 -21508
rect -3301 -21588 -3174 -21572
rect -3301 -21652 -3254 -21588
rect -3190 -21652 -3174 -21588
rect -3301 -21668 -3174 -21652
rect -3301 -21732 -3254 -21668
rect -3190 -21732 -3174 -21668
rect -3301 -21748 -3174 -21732
rect -3301 -21812 -3254 -21748
rect -3190 -21812 -3174 -21748
rect -3301 -21828 -3174 -21812
rect -9620 -21908 -9493 -21892
rect -9620 -21972 -9573 -21908
rect -9509 -21972 -9493 -21908
rect -9620 -21988 -9493 -21972
rect -9620 -22112 -9516 -21988
rect -9620 -22128 -9493 -22112
rect -9620 -22192 -9573 -22128
rect -9509 -22192 -9493 -22128
rect -9620 -22208 -9493 -22192
rect -15939 -22288 -15812 -22272
rect -15939 -22352 -15892 -22288
rect -15828 -22352 -15812 -22288
rect -15939 -22368 -15812 -22352
rect -15939 -22432 -15892 -22368
rect -15828 -22432 -15812 -22368
rect -15939 -22448 -15812 -22432
rect -15939 -22512 -15892 -22448
rect -15828 -22512 -15812 -22448
rect -15939 -22528 -15812 -22512
rect -15939 -22592 -15892 -22528
rect -15828 -22592 -15812 -22528
rect -15939 -22608 -15812 -22592
rect -15939 -22672 -15892 -22608
rect -15828 -22672 -15812 -22608
rect -15939 -22688 -15812 -22672
rect -15939 -22752 -15892 -22688
rect -15828 -22752 -15812 -22688
rect -15939 -22768 -15812 -22752
rect -15939 -22832 -15892 -22768
rect -15828 -22832 -15812 -22768
rect -15939 -22848 -15812 -22832
rect -15939 -22912 -15892 -22848
rect -15828 -22912 -15812 -22848
rect -15939 -22928 -15812 -22912
rect -15939 -22992 -15892 -22928
rect -15828 -22992 -15812 -22928
rect -15939 -23008 -15812 -22992
rect -15939 -23072 -15892 -23008
rect -15828 -23072 -15812 -23008
rect -15939 -23088 -15812 -23072
rect -15939 -23152 -15892 -23088
rect -15828 -23152 -15812 -23088
rect -15939 -23168 -15812 -23152
rect -15939 -23232 -15892 -23168
rect -15828 -23232 -15812 -23168
rect -15939 -23248 -15812 -23232
rect -15939 -23312 -15892 -23248
rect -15828 -23312 -15812 -23248
rect -15939 -23328 -15812 -23312
rect -15939 -23392 -15892 -23328
rect -15828 -23392 -15812 -23328
rect -15939 -23408 -15812 -23392
rect -15939 -23472 -15892 -23408
rect -15828 -23472 -15812 -23408
rect -15939 -23488 -15812 -23472
rect -15939 -23552 -15892 -23488
rect -15828 -23552 -15812 -23488
rect -15939 -23568 -15812 -23552
rect -15939 -23632 -15892 -23568
rect -15828 -23632 -15812 -23568
rect -15939 -23648 -15812 -23632
rect -15939 -23712 -15892 -23648
rect -15828 -23712 -15812 -23648
rect -15939 -23728 -15812 -23712
rect -15939 -23792 -15892 -23728
rect -15828 -23792 -15812 -23728
rect -15939 -23808 -15812 -23792
rect -15939 -23872 -15892 -23808
rect -15828 -23872 -15812 -23808
rect -15939 -23888 -15812 -23872
rect -15939 -23952 -15892 -23888
rect -15828 -23952 -15812 -23888
rect -15939 -23968 -15812 -23952
rect -15939 -24032 -15892 -23968
rect -15828 -24032 -15812 -23968
rect -15939 -24048 -15812 -24032
rect -15939 -24112 -15892 -24048
rect -15828 -24112 -15812 -24048
rect -15939 -24128 -15812 -24112
rect -15939 -24192 -15892 -24128
rect -15828 -24192 -15812 -24128
rect -15939 -24208 -15812 -24192
rect -15939 -24272 -15892 -24208
rect -15828 -24272 -15812 -24208
rect -15939 -24288 -15812 -24272
rect -15939 -24352 -15892 -24288
rect -15828 -24352 -15812 -24288
rect -15939 -24368 -15812 -24352
rect -15939 -24432 -15892 -24368
rect -15828 -24432 -15812 -24368
rect -15939 -24448 -15812 -24432
rect -15939 -24512 -15892 -24448
rect -15828 -24512 -15812 -24448
rect -15939 -24528 -15812 -24512
rect -15939 -24592 -15892 -24528
rect -15828 -24592 -15812 -24528
rect -15939 -24608 -15812 -24592
rect -15939 -24672 -15892 -24608
rect -15828 -24672 -15812 -24608
rect -15939 -24688 -15812 -24672
rect -15939 -24752 -15892 -24688
rect -15828 -24752 -15812 -24688
rect -15939 -24768 -15812 -24752
rect -15939 -24832 -15892 -24768
rect -15828 -24832 -15812 -24768
rect -15939 -24848 -15812 -24832
rect -15939 -24912 -15892 -24848
rect -15828 -24912 -15812 -24848
rect -15939 -24928 -15812 -24912
rect -15939 -24992 -15892 -24928
rect -15828 -24992 -15812 -24928
rect -15939 -25008 -15812 -24992
rect -15939 -25072 -15892 -25008
rect -15828 -25072 -15812 -25008
rect -15939 -25088 -15812 -25072
rect -15939 -25152 -15892 -25088
rect -15828 -25152 -15812 -25088
rect -15939 -25168 -15812 -25152
rect -15939 -25232 -15892 -25168
rect -15828 -25232 -15812 -25168
rect -15939 -25248 -15812 -25232
rect -15939 -25312 -15892 -25248
rect -15828 -25312 -15812 -25248
rect -15939 -25328 -15812 -25312
rect -15939 -25392 -15892 -25328
rect -15828 -25392 -15812 -25328
rect -15939 -25408 -15812 -25392
rect -15939 -25472 -15892 -25408
rect -15828 -25472 -15812 -25408
rect -15939 -25488 -15812 -25472
rect -15939 -25552 -15892 -25488
rect -15828 -25552 -15812 -25488
rect -15939 -25568 -15812 -25552
rect -15939 -25632 -15892 -25568
rect -15828 -25632 -15812 -25568
rect -15939 -25648 -15812 -25632
rect -15939 -25712 -15892 -25648
rect -15828 -25712 -15812 -25648
rect -15939 -25728 -15812 -25712
rect -15939 -25792 -15892 -25728
rect -15828 -25792 -15812 -25728
rect -15939 -25808 -15812 -25792
rect -15939 -25872 -15892 -25808
rect -15828 -25872 -15812 -25808
rect -15939 -25888 -15812 -25872
rect -15939 -25952 -15892 -25888
rect -15828 -25952 -15812 -25888
rect -15939 -25968 -15812 -25952
rect -15939 -26032 -15892 -25968
rect -15828 -26032 -15812 -25968
rect -15939 -26048 -15812 -26032
rect -15939 -26112 -15892 -26048
rect -15828 -26112 -15812 -26048
rect -15939 -26128 -15812 -26112
rect -15939 -26192 -15892 -26128
rect -15828 -26192 -15812 -26128
rect -15939 -26208 -15812 -26192
rect -15939 -26272 -15892 -26208
rect -15828 -26272 -15812 -26208
rect -15939 -26288 -15812 -26272
rect -15939 -26352 -15892 -26288
rect -15828 -26352 -15812 -26288
rect -15939 -26368 -15812 -26352
rect -15939 -26432 -15892 -26368
rect -15828 -26432 -15812 -26368
rect -15939 -26448 -15812 -26432
rect -15939 -26512 -15892 -26448
rect -15828 -26512 -15812 -26448
rect -15939 -26528 -15812 -26512
rect -15939 -26592 -15892 -26528
rect -15828 -26592 -15812 -26528
rect -15939 -26608 -15812 -26592
rect -15939 -26672 -15892 -26608
rect -15828 -26672 -15812 -26608
rect -15939 -26688 -15812 -26672
rect -15939 -26752 -15892 -26688
rect -15828 -26752 -15812 -26688
rect -15939 -26768 -15812 -26752
rect -15939 -26832 -15892 -26768
rect -15828 -26832 -15812 -26768
rect -15939 -26848 -15812 -26832
rect -15939 -26912 -15892 -26848
rect -15828 -26912 -15812 -26848
rect -15939 -26928 -15812 -26912
rect -15939 -26992 -15892 -26928
rect -15828 -26992 -15812 -26928
rect -15939 -27008 -15812 -26992
rect -15939 -27072 -15892 -27008
rect -15828 -27072 -15812 -27008
rect -15939 -27088 -15812 -27072
rect -15939 -27152 -15892 -27088
rect -15828 -27152 -15812 -27088
rect -15939 -27168 -15812 -27152
rect -15939 -27232 -15892 -27168
rect -15828 -27232 -15812 -27168
rect -15939 -27248 -15812 -27232
rect -15939 -27312 -15892 -27248
rect -15828 -27312 -15812 -27248
rect -15939 -27328 -15812 -27312
rect -15939 -27392 -15892 -27328
rect -15828 -27392 -15812 -27328
rect -15939 -27408 -15812 -27392
rect -15939 -27472 -15892 -27408
rect -15828 -27472 -15812 -27408
rect -15939 -27488 -15812 -27472
rect -15939 -27552 -15892 -27488
rect -15828 -27552 -15812 -27488
rect -15939 -27568 -15812 -27552
rect -15939 -27632 -15892 -27568
rect -15828 -27632 -15812 -27568
rect -15939 -27648 -15812 -27632
rect -15939 -27712 -15892 -27648
rect -15828 -27712 -15812 -27648
rect -15939 -27728 -15812 -27712
rect -15939 -27792 -15892 -27728
rect -15828 -27792 -15812 -27728
rect -15939 -27808 -15812 -27792
rect -15939 -27872 -15892 -27808
rect -15828 -27872 -15812 -27808
rect -15939 -27888 -15812 -27872
rect -15939 -27952 -15892 -27888
rect -15828 -27952 -15812 -27888
rect -15939 -27968 -15812 -27952
rect -15939 -28032 -15892 -27968
rect -15828 -28032 -15812 -27968
rect -15939 -28048 -15812 -28032
rect -15939 -28112 -15892 -28048
rect -15828 -28112 -15812 -28048
rect -15939 -28128 -15812 -28112
rect -22258 -28208 -22131 -28192
rect -22258 -28272 -22211 -28208
rect -22147 -28272 -22131 -28208
rect -22258 -28288 -22131 -28272
rect -22258 -28412 -22154 -28288
rect -22258 -28428 -22131 -28412
rect -22258 -28492 -22211 -28428
rect -22147 -28492 -22131 -28428
rect -22258 -28508 -22131 -28492
rect -28577 -28588 -28450 -28572
rect -28577 -28652 -28530 -28588
rect -28466 -28652 -28450 -28588
rect -28577 -28668 -28450 -28652
rect -28577 -28732 -28530 -28668
rect -28466 -28732 -28450 -28668
rect -28577 -28748 -28450 -28732
rect -28577 -28812 -28530 -28748
rect -28466 -28812 -28450 -28748
rect -28577 -28828 -28450 -28812
rect -28577 -28892 -28530 -28828
rect -28466 -28892 -28450 -28828
rect -28577 -28908 -28450 -28892
rect -28577 -28972 -28530 -28908
rect -28466 -28972 -28450 -28908
rect -28577 -28988 -28450 -28972
rect -28577 -29052 -28530 -28988
rect -28466 -29052 -28450 -28988
rect -28577 -29068 -28450 -29052
rect -28577 -29132 -28530 -29068
rect -28466 -29132 -28450 -29068
rect -28577 -29148 -28450 -29132
rect -28577 -29212 -28530 -29148
rect -28466 -29212 -28450 -29148
rect -28577 -29228 -28450 -29212
rect -28577 -29292 -28530 -29228
rect -28466 -29292 -28450 -29228
rect -28577 -29308 -28450 -29292
rect -28577 -29372 -28530 -29308
rect -28466 -29372 -28450 -29308
rect -28577 -29388 -28450 -29372
rect -28577 -29452 -28530 -29388
rect -28466 -29452 -28450 -29388
rect -28577 -29468 -28450 -29452
rect -28577 -29532 -28530 -29468
rect -28466 -29532 -28450 -29468
rect -28577 -29548 -28450 -29532
rect -28577 -29612 -28530 -29548
rect -28466 -29612 -28450 -29548
rect -28577 -29628 -28450 -29612
rect -28577 -29692 -28530 -29628
rect -28466 -29692 -28450 -29628
rect -28577 -29708 -28450 -29692
rect -28577 -29772 -28530 -29708
rect -28466 -29772 -28450 -29708
rect -28577 -29788 -28450 -29772
rect -28577 -29852 -28530 -29788
rect -28466 -29852 -28450 -29788
rect -28577 -29868 -28450 -29852
rect -28577 -29932 -28530 -29868
rect -28466 -29932 -28450 -29868
rect -28577 -29948 -28450 -29932
rect -28577 -30012 -28530 -29948
rect -28466 -30012 -28450 -29948
rect -28577 -30028 -28450 -30012
rect -28577 -30092 -28530 -30028
rect -28466 -30092 -28450 -30028
rect -28577 -30108 -28450 -30092
rect -28577 -30172 -28530 -30108
rect -28466 -30172 -28450 -30108
rect -28577 -30188 -28450 -30172
rect -28577 -30252 -28530 -30188
rect -28466 -30252 -28450 -30188
rect -28577 -30268 -28450 -30252
rect -28577 -30332 -28530 -30268
rect -28466 -30332 -28450 -30268
rect -28577 -30348 -28450 -30332
rect -28577 -30412 -28530 -30348
rect -28466 -30412 -28450 -30348
rect -28577 -30428 -28450 -30412
rect -28577 -30492 -28530 -30428
rect -28466 -30492 -28450 -30428
rect -28577 -30508 -28450 -30492
rect -28577 -30572 -28530 -30508
rect -28466 -30572 -28450 -30508
rect -28577 -30588 -28450 -30572
rect -28577 -30652 -28530 -30588
rect -28466 -30652 -28450 -30588
rect -28577 -30668 -28450 -30652
rect -28577 -30732 -28530 -30668
rect -28466 -30732 -28450 -30668
rect -28577 -30748 -28450 -30732
rect -28577 -30812 -28530 -30748
rect -28466 -30812 -28450 -30748
rect -28577 -30828 -28450 -30812
rect -28577 -30892 -28530 -30828
rect -28466 -30892 -28450 -30828
rect -28577 -30908 -28450 -30892
rect -28577 -30972 -28530 -30908
rect -28466 -30972 -28450 -30908
rect -28577 -30988 -28450 -30972
rect -28577 -31052 -28530 -30988
rect -28466 -31052 -28450 -30988
rect -28577 -31068 -28450 -31052
rect -28577 -31132 -28530 -31068
rect -28466 -31132 -28450 -31068
rect -28577 -31148 -28450 -31132
rect -28577 -31212 -28530 -31148
rect -28466 -31212 -28450 -31148
rect -28577 -31228 -28450 -31212
rect -28577 -31292 -28530 -31228
rect -28466 -31292 -28450 -31228
rect -28577 -31308 -28450 -31292
rect -28577 -31372 -28530 -31308
rect -28466 -31372 -28450 -31308
rect -28577 -31388 -28450 -31372
rect -28577 -31452 -28530 -31388
rect -28466 -31452 -28450 -31388
rect -28577 -31468 -28450 -31452
rect -28577 -31532 -28530 -31468
rect -28466 -31532 -28450 -31468
rect -28577 -31548 -28450 -31532
rect -28577 -31612 -28530 -31548
rect -28466 -31612 -28450 -31548
rect -28577 -31628 -28450 -31612
rect -28577 -31692 -28530 -31628
rect -28466 -31692 -28450 -31628
rect -28577 -31708 -28450 -31692
rect -28577 -31772 -28530 -31708
rect -28466 -31772 -28450 -31708
rect -28577 -31788 -28450 -31772
rect -28577 -31852 -28530 -31788
rect -28466 -31852 -28450 -31788
rect -28577 -31868 -28450 -31852
rect -28577 -31932 -28530 -31868
rect -28466 -31932 -28450 -31868
rect -28577 -31948 -28450 -31932
rect -28577 -32012 -28530 -31948
rect -28466 -32012 -28450 -31948
rect -28577 -32028 -28450 -32012
rect -28577 -32092 -28530 -32028
rect -28466 -32092 -28450 -32028
rect -28577 -32108 -28450 -32092
rect -28577 -32172 -28530 -32108
rect -28466 -32172 -28450 -32108
rect -28577 -32188 -28450 -32172
rect -28577 -32252 -28530 -32188
rect -28466 -32252 -28450 -32188
rect -28577 -32268 -28450 -32252
rect -28577 -32332 -28530 -32268
rect -28466 -32332 -28450 -32268
rect -28577 -32348 -28450 -32332
rect -28577 -32412 -28530 -32348
rect -28466 -32412 -28450 -32348
rect -28577 -32428 -28450 -32412
rect -28577 -32492 -28530 -32428
rect -28466 -32492 -28450 -32428
rect -28577 -32508 -28450 -32492
rect -28577 -32572 -28530 -32508
rect -28466 -32572 -28450 -32508
rect -28577 -32588 -28450 -32572
rect -28577 -32652 -28530 -32588
rect -28466 -32652 -28450 -32588
rect -28577 -32668 -28450 -32652
rect -28577 -32732 -28530 -32668
rect -28466 -32732 -28450 -32668
rect -28577 -32748 -28450 -32732
rect -28577 -32812 -28530 -32748
rect -28466 -32812 -28450 -32748
rect -28577 -32828 -28450 -32812
rect -28577 -32892 -28530 -32828
rect -28466 -32892 -28450 -32828
rect -28577 -32908 -28450 -32892
rect -28577 -32972 -28530 -32908
rect -28466 -32972 -28450 -32908
rect -28577 -32988 -28450 -32972
rect -28577 -33052 -28530 -32988
rect -28466 -33052 -28450 -32988
rect -28577 -33068 -28450 -33052
rect -28577 -33132 -28530 -33068
rect -28466 -33132 -28450 -33068
rect -28577 -33148 -28450 -33132
rect -28577 -33212 -28530 -33148
rect -28466 -33212 -28450 -33148
rect -28577 -33228 -28450 -33212
rect -28577 -33292 -28530 -33228
rect -28466 -33292 -28450 -33228
rect -28577 -33308 -28450 -33292
rect -28577 -33372 -28530 -33308
rect -28466 -33372 -28450 -33308
rect -28577 -33388 -28450 -33372
rect -28577 -33452 -28530 -33388
rect -28466 -33452 -28450 -33388
rect -28577 -33468 -28450 -33452
rect -28577 -33532 -28530 -33468
rect -28466 -33532 -28450 -33468
rect -28577 -33548 -28450 -33532
rect -28577 -33612 -28530 -33548
rect -28466 -33612 -28450 -33548
rect -28577 -33628 -28450 -33612
rect -28577 -33692 -28530 -33628
rect -28466 -33692 -28450 -33628
rect -28577 -33708 -28450 -33692
rect -28577 -33772 -28530 -33708
rect -28466 -33772 -28450 -33708
rect -28577 -33788 -28450 -33772
rect -28577 -33852 -28530 -33788
rect -28466 -33852 -28450 -33788
rect -28577 -33868 -28450 -33852
rect -28577 -33932 -28530 -33868
rect -28466 -33932 -28450 -33868
rect -28577 -33948 -28450 -33932
rect -28577 -34012 -28530 -33948
rect -28466 -34012 -28450 -33948
rect -28577 -34028 -28450 -34012
rect -28577 -34092 -28530 -34028
rect -28466 -34092 -28450 -34028
rect -28577 -34108 -28450 -34092
rect -28577 -34172 -28530 -34108
rect -28466 -34172 -28450 -34108
rect -28577 -34188 -28450 -34172
rect -28577 -34252 -28530 -34188
rect -28466 -34252 -28450 -34188
rect -28577 -34268 -28450 -34252
rect -28577 -34332 -28530 -34268
rect -28466 -34332 -28450 -34268
rect -28577 -34348 -28450 -34332
rect -28577 -34412 -28530 -34348
rect -28466 -34412 -28450 -34348
rect -28577 -34428 -28450 -34412
rect -34896 -34508 -34769 -34492
rect -34896 -34572 -34849 -34508
rect -34785 -34572 -34769 -34508
rect -34896 -34588 -34769 -34572
rect -34896 -34712 -34792 -34588
rect -34896 -34728 -34769 -34712
rect -34896 -34792 -34849 -34728
rect -34785 -34792 -34769 -34728
rect -34896 -34808 -34769 -34792
rect -41215 -34888 -41088 -34872
rect -41215 -34952 -41168 -34888
rect -41104 -34952 -41088 -34888
rect -41215 -34968 -41088 -34952
rect -41215 -35032 -41168 -34968
rect -41104 -35032 -41088 -34968
rect -41215 -35048 -41088 -35032
rect -41215 -35112 -41168 -35048
rect -41104 -35112 -41088 -35048
rect -41215 -35128 -41088 -35112
rect -41215 -35192 -41168 -35128
rect -41104 -35192 -41088 -35128
rect -41215 -35208 -41088 -35192
rect -41215 -35272 -41168 -35208
rect -41104 -35272 -41088 -35208
rect -41215 -35288 -41088 -35272
rect -41215 -35352 -41168 -35288
rect -41104 -35352 -41088 -35288
rect -41215 -35368 -41088 -35352
rect -41215 -35432 -41168 -35368
rect -41104 -35432 -41088 -35368
rect -41215 -35448 -41088 -35432
rect -41215 -35512 -41168 -35448
rect -41104 -35512 -41088 -35448
rect -41215 -35528 -41088 -35512
rect -41215 -35592 -41168 -35528
rect -41104 -35592 -41088 -35528
rect -41215 -35608 -41088 -35592
rect -41215 -35672 -41168 -35608
rect -41104 -35672 -41088 -35608
rect -41215 -35688 -41088 -35672
rect -41215 -35752 -41168 -35688
rect -41104 -35752 -41088 -35688
rect -41215 -35768 -41088 -35752
rect -41215 -35832 -41168 -35768
rect -41104 -35832 -41088 -35768
rect -41215 -35848 -41088 -35832
rect -41215 -35912 -41168 -35848
rect -41104 -35912 -41088 -35848
rect -41215 -35928 -41088 -35912
rect -41215 -35992 -41168 -35928
rect -41104 -35992 -41088 -35928
rect -41215 -36008 -41088 -35992
rect -41215 -36072 -41168 -36008
rect -41104 -36072 -41088 -36008
rect -41215 -36088 -41088 -36072
rect -41215 -36152 -41168 -36088
rect -41104 -36152 -41088 -36088
rect -41215 -36168 -41088 -36152
rect -41215 -36232 -41168 -36168
rect -41104 -36232 -41088 -36168
rect -41215 -36248 -41088 -36232
rect -41215 -36312 -41168 -36248
rect -41104 -36312 -41088 -36248
rect -41215 -36328 -41088 -36312
rect -41215 -36392 -41168 -36328
rect -41104 -36392 -41088 -36328
rect -41215 -36408 -41088 -36392
rect -41215 -36472 -41168 -36408
rect -41104 -36472 -41088 -36408
rect -41215 -36488 -41088 -36472
rect -41215 -36552 -41168 -36488
rect -41104 -36552 -41088 -36488
rect -41215 -36568 -41088 -36552
rect -41215 -36632 -41168 -36568
rect -41104 -36632 -41088 -36568
rect -41215 -36648 -41088 -36632
rect -41215 -36712 -41168 -36648
rect -41104 -36712 -41088 -36648
rect -41215 -36728 -41088 -36712
rect -41215 -36792 -41168 -36728
rect -41104 -36792 -41088 -36728
rect -41215 -36808 -41088 -36792
rect -41215 -36872 -41168 -36808
rect -41104 -36872 -41088 -36808
rect -41215 -36888 -41088 -36872
rect -41215 -36952 -41168 -36888
rect -41104 -36952 -41088 -36888
rect -41215 -36968 -41088 -36952
rect -41215 -37032 -41168 -36968
rect -41104 -37032 -41088 -36968
rect -41215 -37048 -41088 -37032
rect -41215 -37112 -41168 -37048
rect -41104 -37112 -41088 -37048
rect -41215 -37128 -41088 -37112
rect -41215 -37192 -41168 -37128
rect -41104 -37192 -41088 -37128
rect -41215 -37208 -41088 -37192
rect -41215 -37272 -41168 -37208
rect -41104 -37272 -41088 -37208
rect -41215 -37288 -41088 -37272
rect -41215 -37352 -41168 -37288
rect -41104 -37352 -41088 -37288
rect -41215 -37368 -41088 -37352
rect -41215 -37432 -41168 -37368
rect -41104 -37432 -41088 -37368
rect -41215 -37448 -41088 -37432
rect -41215 -37512 -41168 -37448
rect -41104 -37512 -41088 -37448
rect -41215 -37528 -41088 -37512
rect -41215 -37592 -41168 -37528
rect -41104 -37592 -41088 -37528
rect -41215 -37608 -41088 -37592
rect -41215 -37672 -41168 -37608
rect -41104 -37672 -41088 -37608
rect -41215 -37688 -41088 -37672
rect -41215 -37752 -41168 -37688
rect -41104 -37752 -41088 -37688
rect -41215 -37768 -41088 -37752
rect -41215 -37832 -41168 -37768
rect -41104 -37832 -41088 -37768
rect -41215 -37848 -41088 -37832
rect -41215 -37912 -41168 -37848
rect -41104 -37912 -41088 -37848
rect -41215 -37928 -41088 -37912
rect -41215 -37992 -41168 -37928
rect -41104 -37992 -41088 -37928
rect -41215 -38008 -41088 -37992
rect -41215 -38072 -41168 -38008
rect -41104 -38072 -41088 -38008
rect -41215 -38088 -41088 -38072
rect -41215 -38152 -41168 -38088
rect -41104 -38152 -41088 -38088
rect -41215 -38168 -41088 -38152
rect -41215 -38232 -41168 -38168
rect -41104 -38232 -41088 -38168
rect -41215 -38248 -41088 -38232
rect -41215 -38312 -41168 -38248
rect -41104 -38312 -41088 -38248
rect -41215 -38328 -41088 -38312
rect -41215 -38392 -41168 -38328
rect -41104 -38392 -41088 -38328
rect -41215 -38408 -41088 -38392
rect -41215 -38472 -41168 -38408
rect -41104 -38472 -41088 -38408
rect -41215 -38488 -41088 -38472
rect -41215 -38552 -41168 -38488
rect -41104 -38552 -41088 -38488
rect -41215 -38568 -41088 -38552
rect -41215 -38632 -41168 -38568
rect -41104 -38632 -41088 -38568
rect -41215 -38648 -41088 -38632
rect -41215 -38712 -41168 -38648
rect -41104 -38712 -41088 -38648
rect -41215 -38728 -41088 -38712
rect -41215 -38792 -41168 -38728
rect -41104 -38792 -41088 -38728
rect -41215 -38808 -41088 -38792
rect -41215 -38872 -41168 -38808
rect -41104 -38872 -41088 -38808
rect -41215 -38888 -41088 -38872
rect -41215 -38952 -41168 -38888
rect -41104 -38952 -41088 -38888
rect -41215 -38968 -41088 -38952
rect -41215 -39032 -41168 -38968
rect -41104 -39032 -41088 -38968
rect -41215 -39048 -41088 -39032
rect -41215 -39112 -41168 -39048
rect -41104 -39112 -41088 -39048
rect -41215 -39128 -41088 -39112
rect -41215 -39192 -41168 -39128
rect -41104 -39192 -41088 -39128
rect -41215 -39208 -41088 -39192
rect -41215 -39272 -41168 -39208
rect -41104 -39272 -41088 -39208
rect -41215 -39288 -41088 -39272
rect -41215 -39352 -41168 -39288
rect -41104 -39352 -41088 -39288
rect -41215 -39368 -41088 -39352
rect -41215 -39432 -41168 -39368
rect -41104 -39432 -41088 -39368
rect -41215 -39448 -41088 -39432
rect -41215 -39512 -41168 -39448
rect -41104 -39512 -41088 -39448
rect -41215 -39528 -41088 -39512
rect -41215 -39592 -41168 -39528
rect -41104 -39592 -41088 -39528
rect -41215 -39608 -41088 -39592
rect -41215 -39672 -41168 -39608
rect -41104 -39672 -41088 -39608
rect -41215 -39688 -41088 -39672
rect -41215 -39752 -41168 -39688
rect -41104 -39752 -41088 -39688
rect -41215 -39768 -41088 -39752
rect -41215 -39832 -41168 -39768
rect -41104 -39832 -41088 -39768
rect -41215 -39848 -41088 -39832
rect -41215 -39912 -41168 -39848
rect -41104 -39912 -41088 -39848
rect -41215 -39928 -41088 -39912
rect -41215 -39992 -41168 -39928
rect -41104 -39992 -41088 -39928
rect -41215 -40008 -41088 -39992
rect -41215 -40072 -41168 -40008
rect -41104 -40072 -41088 -40008
rect -41215 -40088 -41088 -40072
rect -41215 -40152 -41168 -40088
rect -41104 -40152 -41088 -40088
rect -41215 -40168 -41088 -40152
rect -41215 -40232 -41168 -40168
rect -41104 -40232 -41088 -40168
rect -41215 -40248 -41088 -40232
rect -41215 -40312 -41168 -40248
rect -41104 -40312 -41088 -40248
rect -41215 -40328 -41088 -40312
rect -41215 -40392 -41168 -40328
rect -41104 -40392 -41088 -40328
rect -41215 -40408 -41088 -40392
rect -41215 -40472 -41168 -40408
rect -41104 -40472 -41088 -40408
rect -41215 -40488 -41088 -40472
rect -41215 -40552 -41168 -40488
rect -41104 -40552 -41088 -40488
rect -41215 -40568 -41088 -40552
rect -41215 -40632 -41168 -40568
rect -41104 -40632 -41088 -40568
rect -41215 -40648 -41088 -40632
rect -41215 -40712 -41168 -40648
rect -41104 -40712 -41088 -40648
rect -41215 -40728 -41088 -40712
rect -44335 -41139 -44231 -40761
rect -41215 -40792 -41168 -40728
rect -41104 -40792 -41088 -40728
rect -40925 -34848 -35003 -34839
rect -40925 -40752 -40916 -34848
rect -35012 -40752 -35003 -34848
rect -40925 -40761 -35003 -40752
rect -34896 -34872 -34849 -34808
rect -34785 -34872 -34769 -34808
rect -31697 -34839 -31593 -34461
rect -28577 -34492 -28530 -34428
rect -28466 -34492 -28450 -34428
rect -28287 -28548 -22365 -28539
rect -28287 -34452 -28278 -28548
rect -22374 -34452 -22365 -28548
rect -28287 -34461 -22365 -34452
rect -22258 -28572 -22211 -28508
rect -22147 -28572 -22131 -28508
rect -19059 -28539 -18955 -28161
rect -15939 -28192 -15892 -28128
rect -15828 -28192 -15812 -28128
rect -15649 -22248 -9727 -22239
rect -15649 -28152 -15640 -22248
rect -9736 -28152 -9727 -22248
rect -15649 -28161 -9727 -28152
rect -9620 -22272 -9573 -22208
rect -9509 -22272 -9493 -22208
rect -6421 -22239 -6317 -21861
rect -3301 -21892 -3254 -21828
rect -3190 -21892 -3174 -21828
rect -3011 -15948 2911 -15939
rect -3011 -21852 -3002 -15948
rect 2902 -21852 2911 -15948
rect -3011 -21861 2911 -21852
rect 3018 -15972 3065 -15908
rect 3129 -15972 3145 -15908
rect 6217 -15939 6321 -15561
rect 9337 -15592 9384 -15528
rect 9448 -15592 9464 -15528
rect 9627 -9648 15549 -9639
rect 9627 -15552 9636 -9648
rect 15540 -15552 15549 -9648
rect 9627 -15561 15549 -15552
rect 15656 -9672 15703 -9608
rect 15767 -9672 15783 -9608
rect 18855 -9639 18959 -9261
rect 21975 -9292 22022 -9228
rect 22086 -9292 22102 -9228
rect 22265 -3348 28187 -3339
rect 22265 -9252 22274 -3348
rect 28178 -9252 28187 -3348
rect 22265 -9261 28187 -9252
rect 28294 -3372 28341 -3308
rect 28405 -3372 28421 -3308
rect 31493 -3339 31597 -2961
rect 34613 -2992 34660 -2928
rect 34724 -2992 34740 -2928
rect 34903 2952 40825 2961
rect 34903 -2952 34912 2952
rect 40816 -2952 40825 2952
rect 34903 -2961 40825 -2952
rect 40932 2928 40979 2992
rect 41043 2928 41059 2992
rect 44131 2961 44235 3339
rect 47251 3308 47298 3372
rect 47362 3308 47378 3372
rect 47251 3292 47378 3308
rect 47251 3228 47298 3292
rect 47362 3228 47378 3292
rect 47251 3212 47378 3228
rect 47251 3088 47355 3212
rect 47251 3072 47378 3088
rect 47251 3008 47298 3072
rect 47362 3008 47378 3072
rect 47251 2992 47378 3008
rect 40932 2912 41059 2928
rect 40932 2848 40979 2912
rect 41043 2848 41059 2912
rect 40932 2832 41059 2848
rect 40932 2768 40979 2832
rect 41043 2768 41059 2832
rect 40932 2752 41059 2768
rect 40932 2688 40979 2752
rect 41043 2688 41059 2752
rect 40932 2672 41059 2688
rect 40932 2608 40979 2672
rect 41043 2608 41059 2672
rect 40932 2592 41059 2608
rect 40932 2528 40979 2592
rect 41043 2528 41059 2592
rect 40932 2512 41059 2528
rect 40932 2448 40979 2512
rect 41043 2448 41059 2512
rect 40932 2432 41059 2448
rect 40932 2368 40979 2432
rect 41043 2368 41059 2432
rect 40932 2352 41059 2368
rect 40932 2288 40979 2352
rect 41043 2288 41059 2352
rect 40932 2272 41059 2288
rect 40932 2208 40979 2272
rect 41043 2208 41059 2272
rect 40932 2192 41059 2208
rect 40932 2128 40979 2192
rect 41043 2128 41059 2192
rect 40932 2112 41059 2128
rect 40932 2048 40979 2112
rect 41043 2048 41059 2112
rect 40932 2032 41059 2048
rect 40932 1968 40979 2032
rect 41043 1968 41059 2032
rect 40932 1952 41059 1968
rect 40932 1888 40979 1952
rect 41043 1888 41059 1952
rect 40932 1872 41059 1888
rect 40932 1808 40979 1872
rect 41043 1808 41059 1872
rect 40932 1792 41059 1808
rect 40932 1728 40979 1792
rect 41043 1728 41059 1792
rect 40932 1712 41059 1728
rect 40932 1648 40979 1712
rect 41043 1648 41059 1712
rect 40932 1632 41059 1648
rect 40932 1568 40979 1632
rect 41043 1568 41059 1632
rect 40932 1552 41059 1568
rect 40932 1488 40979 1552
rect 41043 1488 41059 1552
rect 40932 1472 41059 1488
rect 40932 1408 40979 1472
rect 41043 1408 41059 1472
rect 40932 1392 41059 1408
rect 40932 1328 40979 1392
rect 41043 1328 41059 1392
rect 40932 1312 41059 1328
rect 40932 1248 40979 1312
rect 41043 1248 41059 1312
rect 40932 1232 41059 1248
rect 40932 1168 40979 1232
rect 41043 1168 41059 1232
rect 40932 1152 41059 1168
rect 40932 1088 40979 1152
rect 41043 1088 41059 1152
rect 40932 1072 41059 1088
rect 40932 1008 40979 1072
rect 41043 1008 41059 1072
rect 40932 992 41059 1008
rect 40932 928 40979 992
rect 41043 928 41059 992
rect 40932 912 41059 928
rect 40932 848 40979 912
rect 41043 848 41059 912
rect 40932 832 41059 848
rect 40932 768 40979 832
rect 41043 768 41059 832
rect 40932 752 41059 768
rect 40932 688 40979 752
rect 41043 688 41059 752
rect 40932 672 41059 688
rect 40932 608 40979 672
rect 41043 608 41059 672
rect 40932 592 41059 608
rect 40932 528 40979 592
rect 41043 528 41059 592
rect 40932 512 41059 528
rect 40932 448 40979 512
rect 41043 448 41059 512
rect 40932 432 41059 448
rect 40932 368 40979 432
rect 41043 368 41059 432
rect 40932 352 41059 368
rect 40932 288 40979 352
rect 41043 288 41059 352
rect 40932 272 41059 288
rect 40932 208 40979 272
rect 41043 208 41059 272
rect 40932 192 41059 208
rect 40932 128 40979 192
rect 41043 128 41059 192
rect 40932 112 41059 128
rect 40932 48 40979 112
rect 41043 48 41059 112
rect 40932 32 41059 48
rect 40932 -32 40979 32
rect 41043 -32 41059 32
rect 40932 -48 41059 -32
rect 40932 -112 40979 -48
rect 41043 -112 41059 -48
rect 40932 -128 41059 -112
rect 40932 -192 40979 -128
rect 41043 -192 41059 -128
rect 40932 -208 41059 -192
rect 40932 -272 40979 -208
rect 41043 -272 41059 -208
rect 40932 -288 41059 -272
rect 40932 -352 40979 -288
rect 41043 -352 41059 -288
rect 40932 -368 41059 -352
rect 40932 -432 40979 -368
rect 41043 -432 41059 -368
rect 40932 -448 41059 -432
rect 40932 -512 40979 -448
rect 41043 -512 41059 -448
rect 40932 -528 41059 -512
rect 40932 -592 40979 -528
rect 41043 -592 41059 -528
rect 40932 -608 41059 -592
rect 40932 -672 40979 -608
rect 41043 -672 41059 -608
rect 40932 -688 41059 -672
rect 40932 -752 40979 -688
rect 41043 -752 41059 -688
rect 40932 -768 41059 -752
rect 40932 -832 40979 -768
rect 41043 -832 41059 -768
rect 40932 -848 41059 -832
rect 40932 -912 40979 -848
rect 41043 -912 41059 -848
rect 40932 -928 41059 -912
rect 40932 -992 40979 -928
rect 41043 -992 41059 -928
rect 40932 -1008 41059 -992
rect 40932 -1072 40979 -1008
rect 41043 -1072 41059 -1008
rect 40932 -1088 41059 -1072
rect 40932 -1152 40979 -1088
rect 41043 -1152 41059 -1088
rect 40932 -1168 41059 -1152
rect 40932 -1232 40979 -1168
rect 41043 -1232 41059 -1168
rect 40932 -1248 41059 -1232
rect 40932 -1312 40979 -1248
rect 41043 -1312 41059 -1248
rect 40932 -1328 41059 -1312
rect 40932 -1392 40979 -1328
rect 41043 -1392 41059 -1328
rect 40932 -1408 41059 -1392
rect 40932 -1472 40979 -1408
rect 41043 -1472 41059 -1408
rect 40932 -1488 41059 -1472
rect 40932 -1552 40979 -1488
rect 41043 -1552 41059 -1488
rect 40932 -1568 41059 -1552
rect 40932 -1632 40979 -1568
rect 41043 -1632 41059 -1568
rect 40932 -1648 41059 -1632
rect 40932 -1712 40979 -1648
rect 41043 -1712 41059 -1648
rect 40932 -1728 41059 -1712
rect 40932 -1792 40979 -1728
rect 41043 -1792 41059 -1728
rect 40932 -1808 41059 -1792
rect 40932 -1872 40979 -1808
rect 41043 -1872 41059 -1808
rect 40932 -1888 41059 -1872
rect 40932 -1952 40979 -1888
rect 41043 -1952 41059 -1888
rect 40932 -1968 41059 -1952
rect 40932 -2032 40979 -1968
rect 41043 -2032 41059 -1968
rect 40932 -2048 41059 -2032
rect 40932 -2112 40979 -2048
rect 41043 -2112 41059 -2048
rect 40932 -2128 41059 -2112
rect 40932 -2192 40979 -2128
rect 41043 -2192 41059 -2128
rect 40932 -2208 41059 -2192
rect 40932 -2272 40979 -2208
rect 41043 -2272 41059 -2208
rect 40932 -2288 41059 -2272
rect 40932 -2352 40979 -2288
rect 41043 -2352 41059 -2288
rect 40932 -2368 41059 -2352
rect 40932 -2432 40979 -2368
rect 41043 -2432 41059 -2368
rect 40932 -2448 41059 -2432
rect 40932 -2512 40979 -2448
rect 41043 -2512 41059 -2448
rect 40932 -2528 41059 -2512
rect 40932 -2592 40979 -2528
rect 41043 -2592 41059 -2528
rect 40932 -2608 41059 -2592
rect 40932 -2672 40979 -2608
rect 41043 -2672 41059 -2608
rect 40932 -2688 41059 -2672
rect 40932 -2752 40979 -2688
rect 41043 -2752 41059 -2688
rect 40932 -2768 41059 -2752
rect 40932 -2832 40979 -2768
rect 41043 -2832 41059 -2768
rect 40932 -2848 41059 -2832
rect 40932 -2912 40979 -2848
rect 41043 -2912 41059 -2848
rect 40932 -2928 41059 -2912
rect 34613 -3008 34740 -2992
rect 34613 -3072 34660 -3008
rect 34724 -3072 34740 -3008
rect 34613 -3088 34740 -3072
rect 34613 -3212 34717 -3088
rect 34613 -3228 34740 -3212
rect 34613 -3292 34660 -3228
rect 34724 -3292 34740 -3228
rect 34613 -3308 34740 -3292
rect 28294 -3388 28421 -3372
rect 28294 -3452 28341 -3388
rect 28405 -3452 28421 -3388
rect 28294 -3468 28421 -3452
rect 28294 -3532 28341 -3468
rect 28405 -3532 28421 -3468
rect 28294 -3548 28421 -3532
rect 28294 -3612 28341 -3548
rect 28405 -3612 28421 -3548
rect 28294 -3628 28421 -3612
rect 28294 -3692 28341 -3628
rect 28405 -3692 28421 -3628
rect 28294 -3708 28421 -3692
rect 28294 -3772 28341 -3708
rect 28405 -3772 28421 -3708
rect 28294 -3788 28421 -3772
rect 28294 -3852 28341 -3788
rect 28405 -3852 28421 -3788
rect 28294 -3868 28421 -3852
rect 28294 -3932 28341 -3868
rect 28405 -3932 28421 -3868
rect 28294 -3948 28421 -3932
rect 28294 -4012 28341 -3948
rect 28405 -4012 28421 -3948
rect 28294 -4028 28421 -4012
rect 28294 -4092 28341 -4028
rect 28405 -4092 28421 -4028
rect 28294 -4108 28421 -4092
rect 28294 -4172 28341 -4108
rect 28405 -4172 28421 -4108
rect 28294 -4188 28421 -4172
rect 28294 -4252 28341 -4188
rect 28405 -4252 28421 -4188
rect 28294 -4268 28421 -4252
rect 28294 -4332 28341 -4268
rect 28405 -4332 28421 -4268
rect 28294 -4348 28421 -4332
rect 28294 -4412 28341 -4348
rect 28405 -4412 28421 -4348
rect 28294 -4428 28421 -4412
rect 28294 -4492 28341 -4428
rect 28405 -4492 28421 -4428
rect 28294 -4508 28421 -4492
rect 28294 -4572 28341 -4508
rect 28405 -4572 28421 -4508
rect 28294 -4588 28421 -4572
rect 28294 -4652 28341 -4588
rect 28405 -4652 28421 -4588
rect 28294 -4668 28421 -4652
rect 28294 -4732 28341 -4668
rect 28405 -4732 28421 -4668
rect 28294 -4748 28421 -4732
rect 28294 -4812 28341 -4748
rect 28405 -4812 28421 -4748
rect 28294 -4828 28421 -4812
rect 28294 -4892 28341 -4828
rect 28405 -4892 28421 -4828
rect 28294 -4908 28421 -4892
rect 28294 -4972 28341 -4908
rect 28405 -4972 28421 -4908
rect 28294 -4988 28421 -4972
rect 28294 -5052 28341 -4988
rect 28405 -5052 28421 -4988
rect 28294 -5068 28421 -5052
rect 28294 -5132 28341 -5068
rect 28405 -5132 28421 -5068
rect 28294 -5148 28421 -5132
rect 28294 -5212 28341 -5148
rect 28405 -5212 28421 -5148
rect 28294 -5228 28421 -5212
rect 28294 -5292 28341 -5228
rect 28405 -5292 28421 -5228
rect 28294 -5308 28421 -5292
rect 28294 -5372 28341 -5308
rect 28405 -5372 28421 -5308
rect 28294 -5388 28421 -5372
rect 28294 -5452 28341 -5388
rect 28405 -5452 28421 -5388
rect 28294 -5468 28421 -5452
rect 28294 -5532 28341 -5468
rect 28405 -5532 28421 -5468
rect 28294 -5548 28421 -5532
rect 28294 -5612 28341 -5548
rect 28405 -5612 28421 -5548
rect 28294 -5628 28421 -5612
rect 28294 -5692 28341 -5628
rect 28405 -5692 28421 -5628
rect 28294 -5708 28421 -5692
rect 28294 -5772 28341 -5708
rect 28405 -5772 28421 -5708
rect 28294 -5788 28421 -5772
rect 28294 -5852 28341 -5788
rect 28405 -5852 28421 -5788
rect 28294 -5868 28421 -5852
rect 28294 -5932 28341 -5868
rect 28405 -5932 28421 -5868
rect 28294 -5948 28421 -5932
rect 28294 -6012 28341 -5948
rect 28405 -6012 28421 -5948
rect 28294 -6028 28421 -6012
rect 28294 -6092 28341 -6028
rect 28405 -6092 28421 -6028
rect 28294 -6108 28421 -6092
rect 28294 -6172 28341 -6108
rect 28405 -6172 28421 -6108
rect 28294 -6188 28421 -6172
rect 28294 -6252 28341 -6188
rect 28405 -6252 28421 -6188
rect 28294 -6268 28421 -6252
rect 28294 -6332 28341 -6268
rect 28405 -6332 28421 -6268
rect 28294 -6348 28421 -6332
rect 28294 -6412 28341 -6348
rect 28405 -6412 28421 -6348
rect 28294 -6428 28421 -6412
rect 28294 -6492 28341 -6428
rect 28405 -6492 28421 -6428
rect 28294 -6508 28421 -6492
rect 28294 -6572 28341 -6508
rect 28405 -6572 28421 -6508
rect 28294 -6588 28421 -6572
rect 28294 -6652 28341 -6588
rect 28405 -6652 28421 -6588
rect 28294 -6668 28421 -6652
rect 28294 -6732 28341 -6668
rect 28405 -6732 28421 -6668
rect 28294 -6748 28421 -6732
rect 28294 -6812 28341 -6748
rect 28405 -6812 28421 -6748
rect 28294 -6828 28421 -6812
rect 28294 -6892 28341 -6828
rect 28405 -6892 28421 -6828
rect 28294 -6908 28421 -6892
rect 28294 -6972 28341 -6908
rect 28405 -6972 28421 -6908
rect 28294 -6988 28421 -6972
rect 28294 -7052 28341 -6988
rect 28405 -7052 28421 -6988
rect 28294 -7068 28421 -7052
rect 28294 -7132 28341 -7068
rect 28405 -7132 28421 -7068
rect 28294 -7148 28421 -7132
rect 28294 -7212 28341 -7148
rect 28405 -7212 28421 -7148
rect 28294 -7228 28421 -7212
rect 28294 -7292 28341 -7228
rect 28405 -7292 28421 -7228
rect 28294 -7308 28421 -7292
rect 28294 -7372 28341 -7308
rect 28405 -7372 28421 -7308
rect 28294 -7388 28421 -7372
rect 28294 -7452 28341 -7388
rect 28405 -7452 28421 -7388
rect 28294 -7468 28421 -7452
rect 28294 -7532 28341 -7468
rect 28405 -7532 28421 -7468
rect 28294 -7548 28421 -7532
rect 28294 -7612 28341 -7548
rect 28405 -7612 28421 -7548
rect 28294 -7628 28421 -7612
rect 28294 -7692 28341 -7628
rect 28405 -7692 28421 -7628
rect 28294 -7708 28421 -7692
rect 28294 -7772 28341 -7708
rect 28405 -7772 28421 -7708
rect 28294 -7788 28421 -7772
rect 28294 -7852 28341 -7788
rect 28405 -7852 28421 -7788
rect 28294 -7868 28421 -7852
rect 28294 -7932 28341 -7868
rect 28405 -7932 28421 -7868
rect 28294 -7948 28421 -7932
rect 28294 -8012 28341 -7948
rect 28405 -8012 28421 -7948
rect 28294 -8028 28421 -8012
rect 28294 -8092 28341 -8028
rect 28405 -8092 28421 -8028
rect 28294 -8108 28421 -8092
rect 28294 -8172 28341 -8108
rect 28405 -8172 28421 -8108
rect 28294 -8188 28421 -8172
rect 28294 -8252 28341 -8188
rect 28405 -8252 28421 -8188
rect 28294 -8268 28421 -8252
rect 28294 -8332 28341 -8268
rect 28405 -8332 28421 -8268
rect 28294 -8348 28421 -8332
rect 28294 -8412 28341 -8348
rect 28405 -8412 28421 -8348
rect 28294 -8428 28421 -8412
rect 28294 -8492 28341 -8428
rect 28405 -8492 28421 -8428
rect 28294 -8508 28421 -8492
rect 28294 -8572 28341 -8508
rect 28405 -8572 28421 -8508
rect 28294 -8588 28421 -8572
rect 28294 -8652 28341 -8588
rect 28405 -8652 28421 -8588
rect 28294 -8668 28421 -8652
rect 28294 -8732 28341 -8668
rect 28405 -8732 28421 -8668
rect 28294 -8748 28421 -8732
rect 28294 -8812 28341 -8748
rect 28405 -8812 28421 -8748
rect 28294 -8828 28421 -8812
rect 28294 -8892 28341 -8828
rect 28405 -8892 28421 -8828
rect 28294 -8908 28421 -8892
rect 28294 -8972 28341 -8908
rect 28405 -8972 28421 -8908
rect 28294 -8988 28421 -8972
rect 28294 -9052 28341 -8988
rect 28405 -9052 28421 -8988
rect 28294 -9068 28421 -9052
rect 28294 -9132 28341 -9068
rect 28405 -9132 28421 -9068
rect 28294 -9148 28421 -9132
rect 28294 -9212 28341 -9148
rect 28405 -9212 28421 -9148
rect 28294 -9228 28421 -9212
rect 21975 -9308 22102 -9292
rect 21975 -9372 22022 -9308
rect 22086 -9372 22102 -9308
rect 21975 -9388 22102 -9372
rect 21975 -9512 22079 -9388
rect 21975 -9528 22102 -9512
rect 21975 -9592 22022 -9528
rect 22086 -9592 22102 -9528
rect 21975 -9608 22102 -9592
rect 15656 -9688 15783 -9672
rect 15656 -9752 15703 -9688
rect 15767 -9752 15783 -9688
rect 15656 -9768 15783 -9752
rect 15656 -9832 15703 -9768
rect 15767 -9832 15783 -9768
rect 15656 -9848 15783 -9832
rect 15656 -9912 15703 -9848
rect 15767 -9912 15783 -9848
rect 15656 -9928 15783 -9912
rect 15656 -9992 15703 -9928
rect 15767 -9992 15783 -9928
rect 15656 -10008 15783 -9992
rect 15656 -10072 15703 -10008
rect 15767 -10072 15783 -10008
rect 15656 -10088 15783 -10072
rect 15656 -10152 15703 -10088
rect 15767 -10152 15783 -10088
rect 15656 -10168 15783 -10152
rect 15656 -10232 15703 -10168
rect 15767 -10232 15783 -10168
rect 15656 -10248 15783 -10232
rect 15656 -10312 15703 -10248
rect 15767 -10312 15783 -10248
rect 15656 -10328 15783 -10312
rect 15656 -10392 15703 -10328
rect 15767 -10392 15783 -10328
rect 15656 -10408 15783 -10392
rect 15656 -10472 15703 -10408
rect 15767 -10472 15783 -10408
rect 15656 -10488 15783 -10472
rect 15656 -10552 15703 -10488
rect 15767 -10552 15783 -10488
rect 15656 -10568 15783 -10552
rect 15656 -10632 15703 -10568
rect 15767 -10632 15783 -10568
rect 15656 -10648 15783 -10632
rect 15656 -10712 15703 -10648
rect 15767 -10712 15783 -10648
rect 15656 -10728 15783 -10712
rect 15656 -10792 15703 -10728
rect 15767 -10792 15783 -10728
rect 15656 -10808 15783 -10792
rect 15656 -10872 15703 -10808
rect 15767 -10872 15783 -10808
rect 15656 -10888 15783 -10872
rect 15656 -10952 15703 -10888
rect 15767 -10952 15783 -10888
rect 15656 -10968 15783 -10952
rect 15656 -11032 15703 -10968
rect 15767 -11032 15783 -10968
rect 15656 -11048 15783 -11032
rect 15656 -11112 15703 -11048
rect 15767 -11112 15783 -11048
rect 15656 -11128 15783 -11112
rect 15656 -11192 15703 -11128
rect 15767 -11192 15783 -11128
rect 15656 -11208 15783 -11192
rect 15656 -11272 15703 -11208
rect 15767 -11272 15783 -11208
rect 15656 -11288 15783 -11272
rect 15656 -11352 15703 -11288
rect 15767 -11352 15783 -11288
rect 15656 -11368 15783 -11352
rect 15656 -11432 15703 -11368
rect 15767 -11432 15783 -11368
rect 15656 -11448 15783 -11432
rect 15656 -11512 15703 -11448
rect 15767 -11512 15783 -11448
rect 15656 -11528 15783 -11512
rect 15656 -11592 15703 -11528
rect 15767 -11592 15783 -11528
rect 15656 -11608 15783 -11592
rect 15656 -11672 15703 -11608
rect 15767 -11672 15783 -11608
rect 15656 -11688 15783 -11672
rect 15656 -11752 15703 -11688
rect 15767 -11752 15783 -11688
rect 15656 -11768 15783 -11752
rect 15656 -11832 15703 -11768
rect 15767 -11832 15783 -11768
rect 15656 -11848 15783 -11832
rect 15656 -11912 15703 -11848
rect 15767 -11912 15783 -11848
rect 15656 -11928 15783 -11912
rect 15656 -11992 15703 -11928
rect 15767 -11992 15783 -11928
rect 15656 -12008 15783 -11992
rect 15656 -12072 15703 -12008
rect 15767 -12072 15783 -12008
rect 15656 -12088 15783 -12072
rect 15656 -12152 15703 -12088
rect 15767 -12152 15783 -12088
rect 15656 -12168 15783 -12152
rect 15656 -12232 15703 -12168
rect 15767 -12232 15783 -12168
rect 15656 -12248 15783 -12232
rect 15656 -12312 15703 -12248
rect 15767 -12312 15783 -12248
rect 15656 -12328 15783 -12312
rect 15656 -12392 15703 -12328
rect 15767 -12392 15783 -12328
rect 15656 -12408 15783 -12392
rect 15656 -12472 15703 -12408
rect 15767 -12472 15783 -12408
rect 15656 -12488 15783 -12472
rect 15656 -12552 15703 -12488
rect 15767 -12552 15783 -12488
rect 15656 -12568 15783 -12552
rect 15656 -12632 15703 -12568
rect 15767 -12632 15783 -12568
rect 15656 -12648 15783 -12632
rect 15656 -12712 15703 -12648
rect 15767 -12712 15783 -12648
rect 15656 -12728 15783 -12712
rect 15656 -12792 15703 -12728
rect 15767 -12792 15783 -12728
rect 15656 -12808 15783 -12792
rect 15656 -12872 15703 -12808
rect 15767 -12872 15783 -12808
rect 15656 -12888 15783 -12872
rect 15656 -12952 15703 -12888
rect 15767 -12952 15783 -12888
rect 15656 -12968 15783 -12952
rect 15656 -13032 15703 -12968
rect 15767 -13032 15783 -12968
rect 15656 -13048 15783 -13032
rect 15656 -13112 15703 -13048
rect 15767 -13112 15783 -13048
rect 15656 -13128 15783 -13112
rect 15656 -13192 15703 -13128
rect 15767 -13192 15783 -13128
rect 15656 -13208 15783 -13192
rect 15656 -13272 15703 -13208
rect 15767 -13272 15783 -13208
rect 15656 -13288 15783 -13272
rect 15656 -13352 15703 -13288
rect 15767 -13352 15783 -13288
rect 15656 -13368 15783 -13352
rect 15656 -13432 15703 -13368
rect 15767 -13432 15783 -13368
rect 15656 -13448 15783 -13432
rect 15656 -13512 15703 -13448
rect 15767 -13512 15783 -13448
rect 15656 -13528 15783 -13512
rect 15656 -13592 15703 -13528
rect 15767 -13592 15783 -13528
rect 15656 -13608 15783 -13592
rect 15656 -13672 15703 -13608
rect 15767 -13672 15783 -13608
rect 15656 -13688 15783 -13672
rect 15656 -13752 15703 -13688
rect 15767 -13752 15783 -13688
rect 15656 -13768 15783 -13752
rect 15656 -13832 15703 -13768
rect 15767 -13832 15783 -13768
rect 15656 -13848 15783 -13832
rect 15656 -13912 15703 -13848
rect 15767 -13912 15783 -13848
rect 15656 -13928 15783 -13912
rect 15656 -13992 15703 -13928
rect 15767 -13992 15783 -13928
rect 15656 -14008 15783 -13992
rect 15656 -14072 15703 -14008
rect 15767 -14072 15783 -14008
rect 15656 -14088 15783 -14072
rect 15656 -14152 15703 -14088
rect 15767 -14152 15783 -14088
rect 15656 -14168 15783 -14152
rect 15656 -14232 15703 -14168
rect 15767 -14232 15783 -14168
rect 15656 -14248 15783 -14232
rect 15656 -14312 15703 -14248
rect 15767 -14312 15783 -14248
rect 15656 -14328 15783 -14312
rect 15656 -14392 15703 -14328
rect 15767 -14392 15783 -14328
rect 15656 -14408 15783 -14392
rect 15656 -14472 15703 -14408
rect 15767 -14472 15783 -14408
rect 15656 -14488 15783 -14472
rect 15656 -14552 15703 -14488
rect 15767 -14552 15783 -14488
rect 15656 -14568 15783 -14552
rect 15656 -14632 15703 -14568
rect 15767 -14632 15783 -14568
rect 15656 -14648 15783 -14632
rect 15656 -14712 15703 -14648
rect 15767 -14712 15783 -14648
rect 15656 -14728 15783 -14712
rect 15656 -14792 15703 -14728
rect 15767 -14792 15783 -14728
rect 15656 -14808 15783 -14792
rect 15656 -14872 15703 -14808
rect 15767 -14872 15783 -14808
rect 15656 -14888 15783 -14872
rect 15656 -14952 15703 -14888
rect 15767 -14952 15783 -14888
rect 15656 -14968 15783 -14952
rect 15656 -15032 15703 -14968
rect 15767 -15032 15783 -14968
rect 15656 -15048 15783 -15032
rect 15656 -15112 15703 -15048
rect 15767 -15112 15783 -15048
rect 15656 -15128 15783 -15112
rect 15656 -15192 15703 -15128
rect 15767 -15192 15783 -15128
rect 15656 -15208 15783 -15192
rect 15656 -15272 15703 -15208
rect 15767 -15272 15783 -15208
rect 15656 -15288 15783 -15272
rect 15656 -15352 15703 -15288
rect 15767 -15352 15783 -15288
rect 15656 -15368 15783 -15352
rect 15656 -15432 15703 -15368
rect 15767 -15432 15783 -15368
rect 15656 -15448 15783 -15432
rect 15656 -15512 15703 -15448
rect 15767 -15512 15783 -15448
rect 15656 -15528 15783 -15512
rect 9337 -15608 9464 -15592
rect 9337 -15672 9384 -15608
rect 9448 -15672 9464 -15608
rect 9337 -15688 9464 -15672
rect 9337 -15812 9441 -15688
rect 9337 -15828 9464 -15812
rect 9337 -15892 9384 -15828
rect 9448 -15892 9464 -15828
rect 9337 -15908 9464 -15892
rect 3018 -15988 3145 -15972
rect 3018 -16052 3065 -15988
rect 3129 -16052 3145 -15988
rect 3018 -16068 3145 -16052
rect 3018 -16132 3065 -16068
rect 3129 -16132 3145 -16068
rect 3018 -16148 3145 -16132
rect 3018 -16212 3065 -16148
rect 3129 -16212 3145 -16148
rect 3018 -16228 3145 -16212
rect 3018 -16292 3065 -16228
rect 3129 -16292 3145 -16228
rect 3018 -16308 3145 -16292
rect 3018 -16372 3065 -16308
rect 3129 -16372 3145 -16308
rect 3018 -16388 3145 -16372
rect 3018 -16452 3065 -16388
rect 3129 -16452 3145 -16388
rect 3018 -16468 3145 -16452
rect 3018 -16532 3065 -16468
rect 3129 -16532 3145 -16468
rect 3018 -16548 3145 -16532
rect 3018 -16612 3065 -16548
rect 3129 -16612 3145 -16548
rect 3018 -16628 3145 -16612
rect 3018 -16692 3065 -16628
rect 3129 -16692 3145 -16628
rect 3018 -16708 3145 -16692
rect 3018 -16772 3065 -16708
rect 3129 -16772 3145 -16708
rect 3018 -16788 3145 -16772
rect 3018 -16852 3065 -16788
rect 3129 -16852 3145 -16788
rect 3018 -16868 3145 -16852
rect 3018 -16932 3065 -16868
rect 3129 -16932 3145 -16868
rect 3018 -16948 3145 -16932
rect 3018 -17012 3065 -16948
rect 3129 -17012 3145 -16948
rect 3018 -17028 3145 -17012
rect 3018 -17092 3065 -17028
rect 3129 -17092 3145 -17028
rect 3018 -17108 3145 -17092
rect 3018 -17172 3065 -17108
rect 3129 -17172 3145 -17108
rect 3018 -17188 3145 -17172
rect 3018 -17252 3065 -17188
rect 3129 -17252 3145 -17188
rect 3018 -17268 3145 -17252
rect 3018 -17332 3065 -17268
rect 3129 -17332 3145 -17268
rect 3018 -17348 3145 -17332
rect 3018 -17412 3065 -17348
rect 3129 -17412 3145 -17348
rect 3018 -17428 3145 -17412
rect 3018 -17492 3065 -17428
rect 3129 -17492 3145 -17428
rect 3018 -17508 3145 -17492
rect 3018 -17572 3065 -17508
rect 3129 -17572 3145 -17508
rect 3018 -17588 3145 -17572
rect 3018 -17652 3065 -17588
rect 3129 -17652 3145 -17588
rect 3018 -17668 3145 -17652
rect 3018 -17732 3065 -17668
rect 3129 -17732 3145 -17668
rect 3018 -17748 3145 -17732
rect 3018 -17812 3065 -17748
rect 3129 -17812 3145 -17748
rect 3018 -17828 3145 -17812
rect 3018 -17892 3065 -17828
rect 3129 -17892 3145 -17828
rect 3018 -17908 3145 -17892
rect 3018 -17972 3065 -17908
rect 3129 -17972 3145 -17908
rect 3018 -17988 3145 -17972
rect 3018 -18052 3065 -17988
rect 3129 -18052 3145 -17988
rect 3018 -18068 3145 -18052
rect 3018 -18132 3065 -18068
rect 3129 -18132 3145 -18068
rect 3018 -18148 3145 -18132
rect 3018 -18212 3065 -18148
rect 3129 -18212 3145 -18148
rect 3018 -18228 3145 -18212
rect 3018 -18292 3065 -18228
rect 3129 -18292 3145 -18228
rect 3018 -18308 3145 -18292
rect 3018 -18372 3065 -18308
rect 3129 -18372 3145 -18308
rect 3018 -18388 3145 -18372
rect 3018 -18452 3065 -18388
rect 3129 -18452 3145 -18388
rect 3018 -18468 3145 -18452
rect 3018 -18532 3065 -18468
rect 3129 -18532 3145 -18468
rect 3018 -18548 3145 -18532
rect 3018 -18612 3065 -18548
rect 3129 -18612 3145 -18548
rect 3018 -18628 3145 -18612
rect 3018 -18692 3065 -18628
rect 3129 -18692 3145 -18628
rect 3018 -18708 3145 -18692
rect 3018 -18772 3065 -18708
rect 3129 -18772 3145 -18708
rect 3018 -18788 3145 -18772
rect 3018 -18852 3065 -18788
rect 3129 -18852 3145 -18788
rect 3018 -18868 3145 -18852
rect 3018 -18932 3065 -18868
rect 3129 -18932 3145 -18868
rect 3018 -18948 3145 -18932
rect 3018 -19012 3065 -18948
rect 3129 -19012 3145 -18948
rect 3018 -19028 3145 -19012
rect 3018 -19092 3065 -19028
rect 3129 -19092 3145 -19028
rect 3018 -19108 3145 -19092
rect 3018 -19172 3065 -19108
rect 3129 -19172 3145 -19108
rect 3018 -19188 3145 -19172
rect 3018 -19252 3065 -19188
rect 3129 -19252 3145 -19188
rect 3018 -19268 3145 -19252
rect 3018 -19332 3065 -19268
rect 3129 -19332 3145 -19268
rect 3018 -19348 3145 -19332
rect 3018 -19412 3065 -19348
rect 3129 -19412 3145 -19348
rect 3018 -19428 3145 -19412
rect 3018 -19492 3065 -19428
rect 3129 -19492 3145 -19428
rect 3018 -19508 3145 -19492
rect 3018 -19572 3065 -19508
rect 3129 -19572 3145 -19508
rect 3018 -19588 3145 -19572
rect 3018 -19652 3065 -19588
rect 3129 -19652 3145 -19588
rect 3018 -19668 3145 -19652
rect 3018 -19732 3065 -19668
rect 3129 -19732 3145 -19668
rect 3018 -19748 3145 -19732
rect 3018 -19812 3065 -19748
rect 3129 -19812 3145 -19748
rect 3018 -19828 3145 -19812
rect 3018 -19892 3065 -19828
rect 3129 -19892 3145 -19828
rect 3018 -19908 3145 -19892
rect 3018 -19972 3065 -19908
rect 3129 -19972 3145 -19908
rect 3018 -19988 3145 -19972
rect 3018 -20052 3065 -19988
rect 3129 -20052 3145 -19988
rect 3018 -20068 3145 -20052
rect 3018 -20132 3065 -20068
rect 3129 -20132 3145 -20068
rect 3018 -20148 3145 -20132
rect 3018 -20212 3065 -20148
rect 3129 -20212 3145 -20148
rect 3018 -20228 3145 -20212
rect 3018 -20292 3065 -20228
rect 3129 -20292 3145 -20228
rect 3018 -20308 3145 -20292
rect 3018 -20372 3065 -20308
rect 3129 -20372 3145 -20308
rect 3018 -20388 3145 -20372
rect 3018 -20452 3065 -20388
rect 3129 -20452 3145 -20388
rect 3018 -20468 3145 -20452
rect 3018 -20532 3065 -20468
rect 3129 -20532 3145 -20468
rect 3018 -20548 3145 -20532
rect 3018 -20612 3065 -20548
rect 3129 -20612 3145 -20548
rect 3018 -20628 3145 -20612
rect 3018 -20692 3065 -20628
rect 3129 -20692 3145 -20628
rect 3018 -20708 3145 -20692
rect 3018 -20772 3065 -20708
rect 3129 -20772 3145 -20708
rect 3018 -20788 3145 -20772
rect 3018 -20852 3065 -20788
rect 3129 -20852 3145 -20788
rect 3018 -20868 3145 -20852
rect 3018 -20932 3065 -20868
rect 3129 -20932 3145 -20868
rect 3018 -20948 3145 -20932
rect 3018 -21012 3065 -20948
rect 3129 -21012 3145 -20948
rect 3018 -21028 3145 -21012
rect 3018 -21092 3065 -21028
rect 3129 -21092 3145 -21028
rect 3018 -21108 3145 -21092
rect 3018 -21172 3065 -21108
rect 3129 -21172 3145 -21108
rect 3018 -21188 3145 -21172
rect 3018 -21252 3065 -21188
rect 3129 -21252 3145 -21188
rect 3018 -21268 3145 -21252
rect 3018 -21332 3065 -21268
rect 3129 -21332 3145 -21268
rect 3018 -21348 3145 -21332
rect 3018 -21412 3065 -21348
rect 3129 -21412 3145 -21348
rect 3018 -21428 3145 -21412
rect 3018 -21492 3065 -21428
rect 3129 -21492 3145 -21428
rect 3018 -21508 3145 -21492
rect 3018 -21572 3065 -21508
rect 3129 -21572 3145 -21508
rect 3018 -21588 3145 -21572
rect 3018 -21652 3065 -21588
rect 3129 -21652 3145 -21588
rect 3018 -21668 3145 -21652
rect 3018 -21732 3065 -21668
rect 3129 -21732 3145 -21668
rect 3018 -21748 3145 -21732
rect 3018 -21812 3065 -21748
rect 3129 -21812 3145 -21748
rect 3018 -21828 3145 -21812
rect -3301 -21908 -3174 -21892
rect -3301 -21972 -3254 -21908
rect -3190 -21972 -3174 -21908
rect -3301 -21988 -3174 -21972
rect -3301 -22112 -3197 -21988
rect -3301 -22128 -3174 -22112
rect -3301 -22192 -3254 -22128
rect -3190 -22192 -3174 -22128
rect -3301 -22208 -3174 -22192
rect -9620 -22288 -9493 -22272
rect -9620 -22352 -9573 -22288
rect -9509 -22352 -9493 -22288
rect -9620 -22368 -9493 -22352
rect -9620 -22432 -9573 -22368
rect -9509 -22432 -9493 -22368
rect -9620 -22448 -9493 -22432
rect -9620 -22512 -9573 -22448
rect -9509 -22512 -9493 -22448
rect -9620 -22528 -9493 -22512
rect -9620 -22592 -9573 -22528
rect -9509 -22592 -9493 -22528
rect -9620 -22608 -9493 -22592
rect -9620 -22672 -9573 -22608
rect -9509 -22672 -9493 -22608
rect -9620 -22688 -9493 -22672
rect -9620 -22752 -9573 -22688
rect -9509 -22752 -9493 -22688
rect -9620 -22768 -9493 -22752
rect -9620 -22832 -9573 -22768
rect -9509 -22832 -9493 -22768
rect -9620 -22848 -9493 -22832
rect -9620 -22912 -9573 -22848
rect -9509 -22912 -9493 -22848
rect -9620 -22928 -9493 -22912
rect -9620 -22992 -9573 -22928
rect -9509 -22992 -9493 -22928
rect -9620 -23008 -9493 -22992
rect -9620 -23072 -9573 -23008
rect -9509 -23072 -9493 -23008
rect -9620 -23088 -9493 -23072
rect -9620 -23152 -9573 -23088
rect -9509 -23152 -9493 -23088
rect -9620 -23168 -9493 -23152
rect -9620 -23232 -9573 -23168
rect -9509 -23232 -9493 -23168
rect -9620 -23248 -9493 -23232
rect -9620 -23312 -9573 -23248
rect -9509 -23312 -9493 -23248
rect -9620 -23328 -9493 -23312
rect -9620 -23392 -9573 -23328
rect -9509 -23392 -9493 -23328
rect -9620 -23408 -9493 -23392
rect -9620 -23472 -9573 -23408
rect -9509 -23472 -9493 -23408
rect -9620 -23488 -9493 -23472
rect -9620 -23552 -9573 -23488
rect -9509 -23552 -9493 -23488
rect -9620 -23568 -9493 -23552
rect -9620 -23632 -9573 -23568
rect -9509 -23632 -9493 -23568
rect -9620 -23648 -9493 -23632
rect -9620 -23712 -9573 -23648
rect -9509 -23712 -9493 -23648
rect -9620 -23728 -9493 -23712
rect -9620 -23792 -9573 -23728
rect -9509 -23792 -9493 -23728
rect -9620 -23808 -9493 -23792
rect -9620 -23872 -9573 -23808
rect -9509 -23872 -9493 -23808
rect -9620 -23888 -9493 -23872
rect -9620 -23952 -9573 -23888
rect -9509 -23952 -9493 -23888
rect -9620 -23968 -9493 -23952
rect -9620 -24032 -9573 -23968
rect -9509 -24032 -9493 -23968
rect -9620 -24048 -9493 -24032
rect -9620 -24112 -9573 -24048
rect -9509 -24112 -9493 -24048
rect -9620 -24128 -9493 -24112
rect -9620 -24192 -9573 -24128
rect -9509 -24192 -9493 -24128
rect -9620 -24208 -9493 -24192
rect -9620 -24272 -9573 -24208
rect -9509 -24272 -9493 -24208
rect -9620 -24288 -9493 -24272
rect -9620 -24352 -9573 -24288
rect -9509 -24352 -9493 -24288
rect -9620 -24368 -9493 -24352
rect -9620 -24432 -9573 -24368
rect -9509 -24432 -9493 -24368
rect -9620 -24448 -9493 -24432
rect -9620 -24512 -9573 -24448
rect -9509 -24512 -9493 -24448
rect -9620 -24528 -9493 -24512
rect -9620 -24592 -9573 -24528
rect -9509 -24592 -9493 -24528
rect -9620 -24608 -9493 -24592
rect -9620 -24672 -9573 -24608
rect -9509 -24672 -9493 -24608
rect -9620 -24688 -9493 -24672
rect -9620 -24752 -9573 -24688
rect -9509 -24752 -9493 -24688
rect -9620 -24768 -9493 -24752
rect -9620 -24832 -9573 -24768
rect -9509 -24832 -9493 -24768
rect -9620 -24848 -9493 -24832
rect -9620 -24912 -9573 -24848
rect -9509 -24912 -9493 -24848
rect -9620 -24928 -9493 -24912
rect -9620 -24992 -9573 -24928
rect -9509 -24992 -9493 -24928
rect -9620 -25008 -9493 -24992
rect -9620 -25072 -9573 -25008
rect -9509 -25072 -9493 -25008
rect -9620 -25088 -9493 -25072
rect -9620 -25152 -9573 -25088
rect -9509 -25152 -9493 -25088
rect -9620 -25168 -9493 -25152
rect -9620 -25232 -9573 -25168
rect -9509 -25232 -9493 -25168
rect -9620 -25248 -9493 -25232
rect -9620 -25312 -9573 -25248
rect -9509 -25312 -9493 -25248
rect -9620 -25328 -9493 -25312
rect -9620 -25392 -9573 -25328
rect -9509 -25392 -9493 -25328
rect -9620 -25408 -9493 -25392
rect -9620 -25472 -9573 -25408
rect -9509 -25472 -9493 -25408
rect -9620 -25488 -9493 -25472
rect -9620 -25552 -9573 -25488
rect -9509 -25552 -9493 -25488
rect -9620 -25568 -9493 -25552
rect -9620 -25632 -9573 -25568
rect -9509 -25632 -9493 -25568
rect -9620 -25648 -9493 -25632
rect -9620 -25712 -9573 -25648
rect -9509 -25712 -9493 -25648
rect -9620 -25728 -9493 -25712
rect -9620 -25792 -9573 -25728
rect -9509 -25792 -9493 -25728
rect -9620 -25808 -9493 -25792
rect -9620 -25872 -9573 -25808
rect -9509 -25872 -9493 -25808
rect -9620 -25888 -9493 -25872
rect -9620 -25952 -9573 -25888
rect -9509 -25952 -9493 -25888
rect -9620 -25968 -9493 -25952
rect -9620 -26032 -9573 -25968
rect -9509 -26032 -9493 -25968
rect -9620 -26048 -9493 -26032
rect -9620 -26112 -9573 -26048
rect -9509 -26112 -9493 -26048
rect -9620 -26128 -9493 -26112
rect -9620 -26192 -9573 -26128
rect -9509 -26192 -9493 -26128
rect -9620 -26208 -9493 -26192
rect -9620 -26272 -9573 -26208
rect -9509 -26272 -9493 -26208
rect -9620 -26288 -9493 -26272
rect -9620 -26352 -9573 -26288
rect -9509 -26352 -9493 -26288
rect -9620 -26368 -9493 -26352
rect -9620 -26432 -9573 -26368
rect -9509 -26432 -9493 -26368
rect -9620 -26448 -9493 -26432
rect -9620 -26512 -9573 -26448
rect -9509 -26512 -9493 -26448
rect -9620 -26528 -9493 -26512
rect -9620 -26592 -9573 -26528
rect -9509 -26592 -9493 -26528
rect -9620 -26608 -9493 -26592
rect -9620 -26672 -9573 -26608
rect -9509 -26672 -9493 -26608
rect -9620 -26688 -9493 -26672
rect -9620 -26752 -9573 -26688
rect -9509 -26752 -9493 -26688
rect -9620 -26768 -9493 -26752
rect -9620 -26832 -9573 -26768
rect -9509 -26832 -9493 -26768
rect -9620 -26848 -9493 -26832
rect -9620 -26912 -9573 -26848
rect -9509 -26912 -9493 -26848
rect -9620 -26928 -9493 -26912
rect -9620 -26992 -9573 -26928
rect -9509 -26992 -9493 -26928
rect -9620 -27008 -9493 -26992
rect -9620 -27072 -9573 -27008
rect -9509 -27072 -9493 -27008
rect -9620 -27088 -9493 -27072
rect -9620 -27152 -9573 -27088
rect -9509 -27152 -9493 -27088
rect -9620 -27168 -9493 -27152
rect -9620 -27232 -9573 -27168
rect -9509 -27232 -9493 -27168
rect -9620 -27248 -9493 -27232
rect -9620 -27312 -9573 -27248
rect -9509 -27312 -9493 -27248
rect -9620 -27328 -9493 -27312
rect -9620 -27392 -9573 -27328
rect -9509 -27392 -9493 -27328
rect -9620 -27408 -9493 -27392
rect -9620 -27472 -9573 -27408
rect -9509 -27472 -9493 -27408
rect -9620 -27488 -9493 -27472
rect -9620 -27552 -9573 -27488
rect -9509 -27552 -9493 -27488
rect -9620 -27568 -9493 -27552
rect -9620 -27632 -9573 -27568
rect -9509 -27632 -9493 -27568
rect -9620 -27648 -9493 -27632
rect -9620 -27712 -9573 -27648
rect -9509 -27712 -9493 -27648
rect -9620 -27728 -9493 -27712
rect -9620 -27792 -9573 -27728
rect -9509 -27792 -9493 -27728
rect -9620 -27808 -9493 -27792
rect -9620 -27872 -9573 -27808
rect -9509 -27872 -9493 -27808
rect -9620 -27888 -9493 -27872
rect -9620 -27952 -9573 -27888
rect -9509 -27952 -9493 -27888
rect -9620 -27968 -9493 -27952
rect -9620 -28032 -9573 -27968
rect -9509 -28032 -9493 -27968
rect -9620 -28048 -9493 -28032
rect -9620 -28112 -9573 -28048
rect -9509 -28112 -9493 -28048
rect -9620 -28128 -9493 -28112
rect -15939 -28208 -15812 -28192
rect -15939 -28272 -15892 -28208
rect -15828 -28272 -15812 -28208
rect -15939 -28288 -15812 -28272
rect -15939 -28412 -15835 -28288
rect -15939 -28428 -15812 -28412
rect -15939 -28492 -15892 -28428
rect -15828 -28492 -15812 -28428
rect -15939 -28508 -15812 -28492
rect -22258 -28588 -22131 -28572
rect -22258 -28652 -22211 -28588
rect -22147 -28652 -22131 -28588
rect -22258 -28668 -22131 -28652
rect -22258 -28732 -22211 -28668
rect -22147 -28732 -22131 -28668
rect -22258 -28748 -22131 -28732
rect -22258 -28812 -22211 -28748
rect -22147 -28812 -22131 -28748
rect -22258 -28828 -22131 -28812
rect -22258 -28892 -22211 -28828
rect -22147 -28892 -22131 -28828
rect -22258 -28908 -22131 -28892
rect -22258 -28972 -22211 -28908
rect -22147 -28972 -22131 -28908
rect -22258 -28988 -22131 -28972
rect -22258 -29052 -22211 -28988
rect -22147 -29052 -22131 -28988
rect -22258 -29068 -22131 -29052
rect -22258 -29132 -22211 -29068
rect -22147 -29132 -22131 -29068
rect -22258 -29148 -22131 -29132
rect -22258 -29212 -22211 -29148
rect -22147 -29212 -22131 -29148
rect -22258 -29228 -22131 -29212
rect -22258 -29292 -22211 -29228
rect -22147 -29292 -22131 -29228
rect -22258 -29308 -22131 -29292
rect -22258 -29372 -22211 -29308
rect -22147 -29372 -22131 -29308
rect -22258 -29388 -22131 -29372
rect -22258 -29452 -22211 -29388
rect -22147 -29452 -22131 -29388
rect -22258 -29468 -22131 -29452
rect -22258 -29532 -22211 -29468
rect -22147 -29532 -22131 -29468
rect -22258 -29548 -22131 -29532
rect -22258 -29612 -22211 -29548
rect -22147 -29612 -22131 -29548
rect -22258 -29628 -22131 -29612
rect -22258 -29692 -22211 -29628
rect -22147 -29692 -22131 -29628
rect -22258 -29708 -22131 -29692
rect -22258 -29772 -22211 -29708
rect -22147 -29772 -22131 -29708
rect -22258 -29788 -22131 -29772
rect -22258 -29852 -22211 -29788
rect -22147 -29852 -22131 -29788
rect -22258 -29868 -22131 -29852
rect -22258 -29932 -22211 -29868
rect -22147 -29932 -22131 -29868
rect -22258 -29948 -22131 -29932
rect -22258 -30012 -22211 -29948
rect -22147 -30012 -22131 -29948
rect -22258 -30028 -22131 -30012
rect -22258 -30092 -22211 -30028
rect -22147 -30092 -22131 -30028
rect -22258 -30108 -22131 -30092
rect -22258 -30172 -22211 -30108
rect -22147 -30172 -22131 -30108
rect -22258 -30188 -22131 -30172
rect -22258 -30252 -22211 -30188
rect -22147 -30252 -22131 -30188
rect -22258 -30268 -22131 -30252
rect -22258 -30332 -22211 -30268
rect -22147 -30332 -22131 -30268
rect -22258 -30348 -22131 -30332
rect -22258 -30412 -22211 -30348
rect -22147 -30412 -22131 -30348
rect -22258 -30428 -22131 -30412
rect -22258 -30492 -22211 -30428
rect -22147 -30492 -22131 -30428
rect -22258 -30508 -22131 -30492
rect -22258 -30572 -22211 -30508
rect -22147 -30572 -22131 -30508
rect -22258 -30588 -22131 -30572
rect -22258 -30652 -22211 -30588
rect -22147 -30652 -22131 -30588
rect -22258 -30668 -22131 -30652
rect -22258 -30732 -22211 -30668
rect -22147 -30732 -22131 -30668
rect -22258 -30748 -22131 -30732
rect -22258 -30812 -22211 -30748
rect -22147 -30812 -22131 -30748
rect -22258 -30828 -22131 -30812
rect -22258 -30892 -22211 -30828
rect -22147 -30892 -22131 -30828
rect -22258 -30908 -22131 -30892
rect -22258 -30972 -22211 -30908
rect -22147 -30972 -22131 -30908
rect -22258 -30988 -22131 -30972
rect -22258 -31052 -22211 -30988
rect -22147 -31052 -22131 -30988
rect -22258 -31068 -22131 -31052
rect -22258 -31132 -22211 -31068
rect -22147 -31132 -22131 -31068
rect -22258 -31148 -22131 -31132
rect -22258 -31212 -22211 -31148
rect -22147 -31212 -22131 -31148
rect -22258 -31228 -22131 -31212
rect -22258 -31292 -22211 -31228
rect -22147 -31292 -22131 -31228
rect -22258 -31308 -22131 -31292
rect -22258 -31372 -22211 -31308
rect -22147 -31372 -22131 -31308
rect -22258 -31388 -22131 -31372
rect -22258 -31452 -22211 -31388
rect -22147 -31452 -22131 -31388
rect -22258 -31468 -22131 -31452
rect -22258 -31532 -22211 -31468
rect -22147 -31532 -22131 -31468
rect -22258 -31548 -22131 -31532
rect -22258 -31612 -22211 -31548
rect -22147 -31612 -22131 -31548
rect -22258 -31628 -22131 -31612
rect -22258 -31692 -22211 -31628
rect -22147 -31692 -22131 -31628
rect -22258 -31708 -22131 -31692
rect -22258 -31772 -22211 -31708
rect -22147 -31772 -22131 -31708
rect -22258 -31788 -22131 -31772
rect -22258 -31852 -22211 -31788
rect -22147 -31852 -22131 -31788
rect -22258 -31868 -22131 -31852
rect -22258 -31932 -22211 -31868
rect -22147 -31932 -22131 -31868
rect -22258 -31948 -22131 -31932
rect -22258 -32012 -22211 -31948
rect -22147 -32012 -22131 -31948
rect -22258 -32028 -22131 -32012
rect -22258 -32092 -22211 -32028
rect -22147 -32092 -22131 -32028
rect -22258 -32108 -22131 -32092
rect -22258 -32172 -22211 -32108
rect -22147 -32172 -22131 -32108
rect -22258 -32188 -22131 -32172
rect -22258 -32252 -22211 -32188
rect -22147 -32252 -22131 -32188
rect -22258 -32268 -22131 -32252
rect -22258 -32332 -22211 -32268
rect -22147 -32332 -22131 -32268
rect -22258 -32348 -22131 -32332
rect -22258 -32412 -22211 -32348
rect -22147 -32412 -22131 -32348
rect -22258 -32428 -22131 -32412
rect -22258 -32492 -22211 -32428
rect -22147 -32492 -22131 -32428
rect -22258 -32508 -22131 -32492
rect -22258 -32572 -22211 -32508
rect -22147 -32572 -22131 -32508
rect -22258 -32588 -22131 -32572
rect -22258 -32652 -22211 -32588
rect -22147 -32652 -22131 -32588
rect -22258 -32668 -22131 -32652
rect -22258 -32732 -22211 -32668
rect -22147 -32732 -22131 -32668
rect -22258 -32748 -22131 -32732
rect -22258 -32812 -22211 -32748
rect -22147 -32812 -22131 -32748
rect -22258 -32828 -22131 -32812
rect -22258 -32892 -22211 -32828
rect -22147 -32892 -22131 -32828
rect -22258 -32908 -22131 -32892
rect -22258 -32972 -22211 -32908
rect -22147 -32972 -22131 -32908
rect -22258 -32988 -22131 -32972
rect -22258 -33052 -22211 -32988
rect -22147 -33052 -22131 -32988
rect -22258 -33068 -22131 -33052
rect -22258 -33132 -22211 -33068
rect -22147 -33132 -22131 -33068
rect -22258 -33148 -22131 -33132
rect -22258 -33212 -22211 -33148
rect -22147 -33212 -22131 -33148
rect -22258 -33228 -22131 -33212
rect -22258 -33292 -22211 -33228
rect -22147 -33292 -22131 -33228
rect -22258 -33308 -22131 -33292
rect -22258 -33372 -22211 -33308
rect -22147 -33372 -22131 -33308
rect -22258 -33388 -22131 -33372
rect -22258 -33452 -22211 -33388
rect -22147 -33452 -22131 -33388
rect -22258 -33468 -22131 -33452
rect -22258 -33532 -22211 -33468
rect -22147 -33532 -22131 -33468
rect -22258 -33548 -22131 -33532
rect -22258 -33612 -22211 -33548
rect -22147 -33612 -22131 -33548
rect -22258 -33628 -22131 -33612
rect -22258 -33692 -22211 -33628
rect -22147 -33692 -22131 -33628
rect -22258 -33708 -22131 -33692
rect -22258 -33772 -22211 -33708
rect -22147 -33772 -22131 -33708
rect -22258 -33788 -22131 -33772
rect -22258 -33852 -22211 -33788
rect -22147 -33852 -22131 -33788
rect -22258 -33868 -22131 -33852
rect -22258 -33932 -22211 -33868
rect -22147 -33932 -22131 -33868
rect -22258 -33948 -22131 -33932
rect -22258 -34012 -22211 -33948
rect -22147 -34012 -22131 -33948
rect -22258 -34028 -22131 -34012
rect -22258 -34092 -22211 -34028
rect -22147 -34092 -22131 -34028
rect -22258 -34108 -22131 -34092
rect -22258 -34172 -22211 -34108
rect -22147 -34172 -22131 -34108
rect -22258 -34188 -22131 -34172
rect -22258 -34252 -22211 -34188
rect -22147 -34252 -22131 -34188
rect -22258 -34268 -22131 -34252
rect -22258 -34332 -22211 -34268
rect -22147 -34332 -22131 -34268
rect -22258 -34348 -22131 -34332
rect -22258 -34412 -22211 -34348
rect -22147 -34412 -22131 -34348
rect -22258 -34428 -22131 -34412
rect -28577 -34508 -28450 -34492
rect -28577 -34572 -28530 -34508
rect -28466 -34572 -28450 -34508
rect -28577 -34588 -28450 -34572
rect -28577 -34712 -28473 -34588
rect -28577 -34728 -28450 -34712
rect -28577 -34792 -28530 -34728
rect -28466 -34792 -28450 -34728
rect -28577 -34808 -28450 -34792
rect -34896 -34888 -34769 -34872
rect -34896 -34952 -34849 -34888
rect -34785 -34952 -34769 -34888
rect -34896 -34968 -34769 -34952
rect -34896 -35032 -34849 -34968
rect -34785 -35032 -34769 -34968
rect -34896 -35048 -34769 -35032
rect -34896 -35112 -34849 -35048
rect -34785 -35112 -34769 -35048
rect -34896 -35128 -34769 -35112
rect -34896 -35192 -34849 -35128
rect -34785 -35192 -34769 -35128
rect -34896 -35208 -34769 -35192
rect -34896 -35272 -34849 -35208
rect -34785 -35272 -34769 -35208
rect -34896 -35288 -34769 -35272
rect -34896 -35352 -34849 -35288
rect -34785 -35352 -34769 -35288
rect -34896 -35368 -34769 -35352
rect -34896 -35432 -34849 -35368
rect -34785 -35432 -34769 -35368
rect -34896 -35448 -34769 -35432
rect -34896 -35512 -34849 -35448
rect -34785 -35512 -34769 -35448
rect -34896 -35528 -34769 -35512
rect -34896 -35592 -34849 -35528
rect -34785 -35592 -34769 -35528
rect -34896 -35608 -34769 -35592
rect -34896 -35672 -34849 -35608
rect -34785 -35672 -34769 -35608
rect -34896 -35688 -34769 -35672
rect -34896 -35752 -34849 -35688
rect -34785 -35752 -34769 -35688
rect -34896 -35768 -34769 -35752
rect -34896 -35832 -34849 -35768
rect -34785 -35832 -34769 -35768
rect -34896 -35848 -34769 -35832
rect -34896 -35912 -34849 -35848
rect -34785 -35912 -34769 -35848
rect -34896 -35928 -34769 -35912
rect -34896 -35992 -34849 -35928
rect -34785 -35992 -34769 -35928
rect -34896 -36008 -34769 -35992
rect -34896 -36072 -34849 -36008
rect -34785 -36072 -34769 -36008
rect -34896 -36088 -34769 -36072
rect -34896 -36152 -34849 -36088
rect -34785 -36152 -34769 -36088
rect -34896 -36168 -34769 -36152
rect -34896 -36232 -34849 -36168
rect -34785 -36232 -34769 -36168
rect -34896 -36248 -34769 -36232
rect -34896 -36312 -34849 -36248
rect -34785 -36312 -34769 -36248
rect -34896 -36328 -34769 -36312
rect -34896 -36392 -34849 -36328
rect -34785 -36392 -34769 -36328
rect -34896 -36408 -34769 -36392
rect -34896 -36472 -34849 -36408
rect -34785 -36472 -34769 -36408
rect -34896 -36488 -34769 -36472
rect -34896 -36552 -34849 -36488
rect -34785 -36552 -34769 -36488
rect -34896 -36568 -34769 -36552
rect -34896 -36632 -34849 -36568
rect -34785 -36632 -34769 -36568
rect -34896 -36648 -34769 -36632
rect -34896 -36712 -34849 -36648
rect -34785 -36712 -34769 -36648
rect -34896 -36728 -34769 -36712
rect -34896 -36792 -34849 -36728
rect -34785 -36792 -34769 -36728
rect -34896 -36808 -34769 -36792
rect -34896 -36872 -34849 -36808
rect -34785 -36872 -34769 -36808
rect -34896 -36888 -34769 -36872
rect -34896 -36952 -34849 -36888
rect -34785 -36952 -34769 -36888
rect -34896 -36968 -34769 -36952
rect -34896 -37032 -34849 -36968
rect -34785 -37032 -34769 -36968
rect -34896 -37048 -34769 -37032
rect -34896 -37112 -34849 -37048
rect -34785 -37112 -34769 -37048
rect -34896 -37128 -34769 -37112
rect -34896 -37192 -34849 -37128
rect -34785 -37192 -34769 -37128
rect -34896 -37208 -34769 -37192
rect -34896 -37272 -34849 -37208
rect -34785 -37272 -34769 -37208
rect -34896 -37288 -34769 -37272
rect -34896 -37352 -34849 -37288
rect -34785 -37352 -34769 -37288
rect -34896 -37368 -34769 -37352
rect -34896 -37432 -34849 -37368
rect -34785 -37432 -34769 -37368
rect -34896 -37448 -34769 -37432
rect -34896 -37512 -34849 -37448
rect -34785 -37512 -34769 -37448
rect -34896 -37528 -34769 -37512
rect -34896 -37592 -34849 -37528
rect -34785 -37592 -34769 -37528
rect -34896 -37608 -34769 -37592
rect -34896 -37672 -34849 -37608
rect -34785 -37672 -34769 -37608
rect -34896 -37688 -34769 -37672
rect -34896 -37752 -34849 -37688
rect -34785 -37752 -34769 -37688
rect -34896 -37768 -34769 -37752
rect -34896 -37832 -34849 -37768
rect -34785 -37832 -34769 -37768
rect -34896 -37848 -34769 -37832
rect -34896 -37912 -34849 -37848
rect -34785 -37912 -34769 -37848
rect -34896 -37928 -34769 -37912
rect -34896 -37992 -34849 -37928
rect -34785 -37992 -34769 -37928
rect -34896 -38008 -34769 -37992
rect -34896 -38072 -34849 -38008
rect -34785 -38072 -34769 -38008
rect -34896 -38088 -34769 -38072
rect -34896 -38152 -34849 -38088
rect -34785 -38152 -34769 -38088
rect -34896 -38168 -34769 -38152
rect -34896 -38232 -34849 -38168
rect -34785 -38232 -34769 -38168
rect -34896 -38248 -34769 -38232
rect -34896 -38312 -34849 -38248
rect -34785 -38312 -34769 -38248
rect -34896 -38328 -34769 -38312
rect -34896 -38392 -34849 -38328
rect -34785 -38392 -34769 -38328
rect -34896 -38408 -34769 -38392
rect -34896 -38472 -34849 -38408
rect -34785 -38472 -34769 -38408
rect -34896 -38488 -34769 -38472
rect -34896 -38552 -34849 -38488
rect -34785 -38552 -34769 -38488
rect -34896 -38568 -34769 -38552
rect -34896 -38632 -34849 -38568
rect -34785 -38632 -34769 -38568
rect -34896 -38648 -34769 -38632
rect -34896 -38712 -34849 -38648
rect -34785 -38712 -34769 -38648
rect -34896 -38728 -34769 -38712
rect -34896 -38792 -34849 -38728
rect -34785 -38792 -34769 -38728
rect -34896 -38808 -34769 -38792
rect -34896 -38872 -34849 -38808
rect -34785 -38872 -34769 -38808
rect -34896 -38888 -34769 -38872
rect -34896 -38952 -34849 -38888
rect -34785 -38952 -34769 -38888
rect -34896 -38968 -34769 -38952
rect -34896 -39032 -34849 -38968
rect -34785 -39032 -34769 -38968
rect -34896 -39048 -34769 -39032
rect -34896 -39112 -34849 -39048
rect -34785 -39112 -34769 -39048
rect -34896 -39128 -34769 -39112
rect -34896 -39192 -34849 -39128
rect -34785 -39192 -34769 -39128
rect -34896 -39208 -34769 -39192
rect -34896 -39272 -34849 -39208
rect -34785 -39272 -34769 -39208
rect -34896 -39288 -34769 -39272
rect -34896 -39352 -34849 -39288
rect -34785 -39352 -34769 -39288
rect -34896 -39368 -34769 -39352
rect -34896 -39432 -34849 -39368
rect -34785 -39432 -34769 -39368
rect -34896 -39448 -34769 -39432
rect -34896 -39512 -34849 -39448
rect -34785 -39512 -34769 -39448
rect -34896 -39528 -34769 -39512
rect -34896 -39592 -34849 -39528
rect -34785 -39592 -34769 -39528
rect -34896 -39608 -34769 -39592
rect -34896 -39672 -34849 -39608
rect -34785 -39672 -34769 -39608
rect -34896 -39688 -34769 -39672
rect -34896 -39752 -34849 -39688
rect -34785 -39752 -34769 -39688
rect -34896 -39768 -34769 -39752
rect -34896 -39832 -34849 -39768
rect -34785 -39832 -34769 -39768
rect -34896 -39848 -34769 -39832
rect -34896 -39912 -34849 -39848
rect -34785 -39912 -34769 -39848
rect -34896 -39928 -34769 -39912
rect -34896 -39992 -34849 -39928
rect -34785 -39992 -34769 -39928
rect -34896 -40008 -34769 -39992
rect -34896 -40072 -34849 -40008
rect -34785 -40072 -34769 -40008
rect -34896 -40088 -34769 -40072
rect -34896 -40152 -34849 -40088
rect -34785 -40152 -34769 -40088
rect -34896 -40168 -34769 -40152
rect -34896 -40232 -34849 -40168
rect -34785 -40232 -34769 -40168
rect -34896 -40248 -34769 -40232
rect -34896 -40312 -34849 -40248
rect -34785 -40312 -34769 -40248
rect -34896 -40328 -34769 -40312
rect -34896 -40392 -34849 -40328
rect -34785 -40392 -34769 -40328
rect -34896 -40408 -34769 -40392
rect -34896 -40472 -34849 -40408
rect -34785 -40472 -34769 -40408
rect -34896 -40488 -34769 -40472
rect -34896 -40552 -34849 -40488
rect -34785 -40552 -34769 -40488
rect -34896 -40568 -34769 -40552
rect -34896 -40632 -34849 -40568
rect -34785 -40632 -34769 -40568
rect -34896 -40648 -34769 -40632
rect -34896 -40712 -34849 -40648
rect -34785 -40712 -34769 -40648
rect -34896 -40728 -34769 -40712
rect -41215 -40808 -41088 -40792
rect -41215 -40872 -41168 -40808
rect -41104 -40872 -41088 -40808
rect -41215 -40888 -41088 -40872
rect -41215 -41012 -41111 -40888
rect -41215 -41028 -41088 -41012
rect -41215 -41092 -41168 -41028
rect -41104 -41092 -41088 -41028
rect -41215 -41108 -41088 -41092
rect -47244 -41148 -41322 -41139
rect -47244 -47052 -47235 -41148
rect -41331 -47052 -41322 -41148
rect -47244 -47061 -41322 -47052
rect -41215 -41172 -41168 -41108
rect -41104 -41172 -41088 -41108
rect -38016 -41139 -37912 -40761
rect -34896 -40792 -34849 -40728
rect -34785 -40792 -34769 -40728
rect -34606 -34848 -28684 -34839
rect -34606 -40752 -34597 -34848
rect -28693 -40752 -28684 -34848
rect -34606 -40761 -28684 -40752
rect -28577 -34872 -28530 -34808
rect -28466 -34872 -28450 -34808
rect -25378 -34839 -25274 -34461
rect -22258 -34492 -22211 -34428
rect -22147 -34492 -22131 -34428
rect -21968 -28548 -16046 -28539
rect -21968 -34452 -21959 -28548
rect -16055 -34452 -16046 -28548
rect -21968 -34461 -16046 -34452
rect -15939 -28572 -15892 -28508
rect -15828 -28572 -15812 -28508
rect -12740 -28539 -12636 -28161
rect -9620 -28192 -9573 -28128
rect -9509 -28192 -9493 -28128
rect -9330 -22248 -3408 -22239
rect -9330 -28152 -9321 -22248
rect -3417 -28152 -3408 -22248
rect -9330 -28161 -3408 -28152
rect -3301 -22272 -3254 -22208
rect -3190 -22272 -3174 -22208
rect -102 -22239 2 -21861
rect 3018 -21892 3065 -21828
rect 3129 -21892 3145 -21828
rect 3308 -15948 9230 -15939
rect 3308 -21852 3317 -15948
rect 9221 -21852 9230 -15948
rect 3308 -21861 9230 -21852
rect 9337 -15972 9384 -15908
rect 9448 -15972 9464 -15908
rect 12536 -15939 12640 -15561
rect 15656 -15592 15703 -15528
rect 15767 -15592 15783 -15528
rect 15946 -9648 21868 -9639
rect 15946 -15552 15955 -9648
rect 21859 -15552 21868 -9648
rect 15946 -15561 21868 -15552
rect 21975 -9672 22022 -9608
rect 22086 -9672 22102 -9608
rect 25174 -9639 25278 -9261
rect 28294 -9292 28341 -9228
rect 28405 -9292 28421 -9228
rect 28584 -3348 34506 -3339
rect 28584 -9252 28593 -3348
rect 34497 -9252 34506 -3348
rect 28584 -9261 34506 -9252
rect 34613 -3372 34660 -3308
rect 34724 -3372 34740 -3308
rect 37812 -3339 37916 -2961
rect 40932 -2992 40979 -2928
rect 41043 -2992 41059 -2928
rect 41222 2952 47144 2961
rect 41222 -2952 41231 2952
rect 47135 -2952 47144 2952
rect 41222 -2961 47144 -2952
rect 47251 2928 47298 2992
rect 47362 2928 47378 2992
rect 47251 2912 47378 2928
rect 47251 2848 47298 2912
rect 47362 2848 47378 2912
rect 47251 2832 47378 2848
rect 47251 2768 47298 2832
rect 47362 2768 47378 2832
rect 47251 2752 47378 2768
rect 47251 2688 47298 2752
rect 47362 2688 47378 2752
rect 47251 2672 47378 2688
rect 47251 2608 47298 2672
rect 47362 2608 47378 2672
rect 47251 2592 47378 2608
rect 47251 2528 47298 2592
rect 47362 2528 47378 2592
rect 47251 2512 47378 2528
rect 47251 2448 47298 2512
rect 47362 2448 47378 2512
rect 47251 2432 47378 2448
rect 47251 2368 47298 2432
rect 47362 2368 47378 2432
rect 47251 2352 47378 2368
rect 47251 2288 47298 2352
rect 47362 2288 47378 2352
rect 47251 2272 47378 2288
rect 47251 2208 47298 2272
rect 47362 2208 47378 2272
rect 47251 2192 47378 2208
rect 47251 2128 47298 2192
rect 47362 2128 47378 2192
rect 47251 2112 47378 2128
rect 47251 2048 47298 2112
rect 47362 2048 47378 2112
rect 47251 2032 47378 2048
rect 47251 1968 47298 2032
rect 47362 1968 47378 2032
rect 47251 1952 47378 1968
rect 47251 1888 47298 1952
rect 47362 1888 47378 1952
rect 47251 1872 47378 1888
rect 47251 1808 47298 1872
rect 47362 1808 47378 1872
rect 47251 1792 47378 1808
rect 47251 1728 47298 1792
rect 47362 1728 47378 1792
rect 47251 1712 47378 1728
rect 47251 1648 47298 1712
rect 47362 1648 47378 1712
rect 47251 1632 47378 1648
rect 47251 1568 47298 1632
rect 47362 1568 47378 1632
rect 47251 1552 47378 1568
rect 47251 1488 47298 1552
rect 47362 1488 47378 1552
rect 47251 1472 47378 1488
rect 47251 1408 47298 1472
rect 47362 1408 47378 1472
rect 47251 1392 47378 1408
rect 47251 1328 47298 1392
rect 47362 1328 47378 1392
rect 47251 1312 47378 1328
rect 47251 1248 47298 1312
rect 47362 1248 47378 1312
rect 47251 1232 47378 1248
rect 47251 1168 47298 1232
rect 47362 1168 47378 1232
rect 47251 1152 47378 1168
rect 47251 1088 47298 1152
rect 47362 1088 47378 1152
rect 47251 1072 47378 1088
rect 47251 1008 47298 1072
rect 47362 1008 47378 1072
rect 47251 992 47378 1008
rect 47251 928 47298 992
rect 47362 928 47378 992
rect 47251 912 47378 928
rect 47251 848 47298 912
rect 47362 848 47378 912
rect 47251 832 47378 848
rect 47251 768 47298 832
rect 47362 768 47378 832
rect 47251 752 47378 768
rect 47251 688 47298 752
rect 47362 688 47378 752
rect 47251 672 47378 688
rect 47251 608 47298 672
rect 47362 608 47378 672
rect 47251 592 47378 608
rect 47251 528 47298 592
rect 47362 528 47378 592
rect 47251 512 47378 528
rect 47251 448 47298 512
rect 47362 448 47378 512
rect 47251 432 47378 448
rect 47251 368 47298 432
rect 47362 368 47378 432
rect 47251 352 47378 368
rect 47251 288 47298 352
rect 47362 288 47378 352
rect 47251 272 47378 288
rect 47251 208 47298 272
rect 47362 208 47378 272
rect 47251 192 47378 208
rect 47251 128 47298 192
rect 47362 128 47378 192
rect 47251 112 47378 128
rect 47251 48 47298 112
rect 47362 48 47378 112
rect 47251 32 47378 48
rect 47251 -32 47298 32
rect 47362 -32 47378 32
rect 47251 -48 47378 -32
rect 47251 -112 47298 -48
rect 47362 -112 47378 -48
rect 47251 -128 47378 -112
rect 47251 -192 47298 -128
rect 47362 -192 47378 -128
rect 47251 -208 47378 -192
rect 47251 -272 47298 -208
rect 47362 -272 47378 -208
rect 47251 -288 47378 -272
rect 47251 -352 47298 -288
rect 47362 -352 47378 -288
rect 47251 -368 47378 -352
rect 47251 -432 47298 -368
rect 47362 -432 47378 -368
rect 47251 -448 47378 -432
rect 47251 -512 47298 -448
rect 47362 -512 47378 -448
rect 47251 -528 47378 -512
rect 47251 -592 47298 -528
rect 47362 -592 47378 -528
rect 47251 -608 47378 -592
rect 47251 -672 47298 -608
rect 47362 -672 47378 -608
rect 47251 -688 47378 -672
rect 47251 -752 47298 -688
rect 47362 -752 47378 -688
rect 47251 -768 47378 -752
rect 47251 -832 47298 -768
rect 47362 -832 47378 -768
rect 47251 -848 47378 -832
rect 47251 -912 47298 -848
rect 47362 -912 47378 -848
rect 47251 -928 47378 -912
rect 47251 -992 47298 -928
rect 47362 -992 47378 -928
rect 47251 -1008 47378 -992
rect 47251 -1072 47298 -1008
rect 47362 -1072 47378 -1008
rect 47251 -1088 47378 -1072
rect 47251 -1152 47298 -1088
rect 47362 -1152 47378 -1088
rect 47251 -1168 47378 -1152
rect 47251 -1232 47298 -1168
rect 47362 -1232 47378 -1168
rect 47251 -1248 47378 -1232
rect 47251 -1312 47298 -1248
rect 47362 -1312 47378 -1248
rect 47251 -1328 47378 -1312
rect 47251 -1392 47298 -1328
rect 47362 -1392 47378 -1328
rect 47251 -1408 47378 -1392
rect 47251 -1472 47298 -1408
rect 47362 -1472 47378 -1408
rect 47251 -1488 47378 -1472
rect 47251 -1552 47298 -1488
rect 47362 -1552 47378 -1488
rect 47251 -1568 47378 -1552
rect 47251 -1632 47298 -1568
rect 47362 -1632 47378 -1568
rect 47251 -1648 47378 -1632
rect 47251 -1712 47298 -1648
rect 47362 -1712 47378 -1648
rect 47251 -1728 47378 -1712
rect 47251 -1792 47298 -1728
rect 47362 -1792 47378 -1728
rect 47251 -1808 47378 -1792
rect 47251 -1872 47298 -1808
rect 47362 -1872 47378 -1808
rect 47251 -1888 47378 -1872
rect 47251 -1952 47298 -1888
rect 47362 -1952 47378 -1888
rect 47251 -1968 47378 -1952
rect 47251 -2032 47298 -1968
rect 47362 -2032 47378 -1968
rect 47251 -2048 47378 -2032
rect 47251 -2112 47298 -2048
rect 47362 -2112 47378 -2048
rect 47251 -2128 47378 -2112
rect 47251 -2192 47298 -2128
rect 47362 -2192 47378 -2128
rect 47251 -2208 47378 -2192
rect 47251 -2272 47298 -2208
rect 47362 -2272 47378 -2208
rect 47251 -2288 47378 -2272
rect 47251 -2352 47298 -2288
rect 47362 -2352 47378 -2288
rect 47251 -2368 47378 -2352
rect 47251 -2432 47298 -2368
rect 47362 -2432 47378 -2368
rect 47251 -2448 47378 -2432
rect 47251 -2512 47298 -2448
rect 47362 -2512 47378 -2448
rect 47251 -2528 47378 -2512
rect 47251 -2592 47298 -2528
rect 47362 -2592 47378 -2528
rect 47251 -2608 47378 -2592
rect 47251 -2672 47298 -2608
rect 47362 -2672 47378 -2608
rect 47251 -2688 47378 -2672
rect 47251 -2752 47298 -2688
rect 47362 -2752 47378 -2688
rect 47251 -2768 47378 -2752
rect 47251 -2832 47298 -2768
rect 47362 -2832 47378 -2768
rect 47251 -2848 47378 -2832
rect 47251 -2912 47298 -2848
rect 47362 -2912 47378 -2848
rect 47251 -2928 47378 -2912
rect 40932 -3008 41059 -2992
rect 40932 -3072 40979 -3008
rect 41043 -3072 41059 -3008
rect 40932 -3088 41059 -3072
rect 40932 -3212 41036 -3088
rect 40932 -3228 41059 -3212
rect 40932 -3292 40979 -3228
rect 41043 -3292 41059 -3228
rect 40932 -3308 41059 -3292
rect 34613 -3388 34740 -3372
rect 34613 -3452 34660 -3388
rect 34724 -3452 34740 -3388
rect 34613 -3468 34740 -3452
rect 34613 -3532 34660 -3468
rect 34724 -3532 34740 -3468
rect 34613 -3548 34740 -3532
rect 34613 -3612 34660 -3548
rect 34724 -3612 34740 -3548
rect 34613 -3628 34740 -3612
rect 34613 -3692 34660 -3628
rect 34724 -3692 34740 -3628
rect 34613 -3708 34740 -3692
rect 34613 -3772 34660 -3708
rect 34724 -3772 34740 -3708
rect 34613 -3788 34740 -3772
rect 34613 -3852 34660 -3788
rect 34724 -3852 34740 -3788
rect 34613 -3868 34740 -3852
rect 34613 -3932 34660 -3868
rect 34724 -3932 34740 -3868
rect 34613 -3948 34740 -3932
rect 34613 -4012 34660 -3948
rect 34724 -4012 34740 -3948
rect 34613 -4028 34740 -4012
rect 34613 -4092 34660 -4028
rect 34724 -4092 34740 -4028
rect 34613 -4108 34740 -4092
rect 34613 -4172 34660 -4108
rect 34724 -4172 34740 -4108
rect 34613 -4188 34740 -4172
rect 34613 -4252 34660 -4188
rect 34724 -4252 34740 -4188
rect 34613 -4268 34740 -4252
rect 34613 -4332 34660 -4268
rect 34724 -4332 34740 -4268
rect 34613 -4348 34740 -4332
rect 34613 -4412 34660 -4348
rect 34724 -4412 34740 -4348
rect 34613 -4428 34740 -4412
rect 34613 -4492 34660 -4428
rect 34724 -4492 34740 -4428
rect 34613 -4508 34740 -4492
rect 34613 -4572 34660 -4508
rect 34724 -4572 34740 -4508
rect 34613 -4588 34740 -4572
rect 34613 -4652 34660 -4588
rect 34724 -4652 34740 -4588
rect 34613 -4668 34740 -4652
rect 34613 -4732 34660 -4668
rect 34724 -4732 34740 -4668
rect 34613 -4748 34740 -4732
rect 34613 -4812 34660 -4748
rect 34724 -4812 34740 -4748
rect 34613 -4828 34740 -4812
rect 34613 -4892 34660 -4828
rect 34724 -4892 34740 -4828
rect 34613 -4908 34740 -4892
rect 34613 -4972 34660 -4908
rect 34724 -4972 34740 -4908
rect 34613 -4988 34740 -4972
rect 34613 -5052 34660 -4988
rect 34724 -5052 34740 -4988
rect 34613 -5068 34740 -5052
rect 34613 -5132 34660 -5068
rect 34724 -5132 34740 -5068
rect 34613 -5148 34740 -5132
rect 34613 -5212 34660 -5148
rect 34724 -5212 34740 -5148
rect 34613 -5228 34740 -5212
rect 34613 -5292 34660 -5228
rect 34724 -5292 34740 -5228
rect 34613 -5308 34740 -5292
rect 34613 -5372 34660 -5308
rect 34724 -5372 34740 -5308
rect 34613 -5388 34740 -5372
rect 34613 -5452 34660 -5388
rect 34724 -5452 34740 -5388
rect 34613 -5468 34740 -5452
rect 34613 -5532 34660 -5468
rect 34724 -5532 34740 -5468
rect 34613 -5548 34740 -5532
rect 34613 -5612 34660 -5548
rect 34724 -5612 34740 -5548
rect 34613 -5628 34740 -5612
rect 34613 -5692 34660 -5628
rect 34724 -5692 34740 -5628
rect 34613 -5708 34740 -5692
rect 34613 -5772 34660 -5708
rect 34724 -5772 34740 -5708
rect 34613 -5788 34740 -5772
rect 34613 -5852 34660 -5788
rect 34724 -5852 34740 -5788
rect 34613 -5868 34740 -5852
rect 34613 -5932 34660 -5868
rect 34724 -5932 34740 -5868
rect 34613 -5948 34740 -5932
rect 34613 -6012 34660 -5948
rect 34724 -6012 34740 -5948
rect 34613 -6028 34740 -6012
rect 34613 -6092 34660 -6028
rect 34724 -6092 34740 -6028
rect 34613 -6108 34740 -6092
rect 34613 -6172 34660 -6108
rect 34724 -6172 34740 -6108
rect 34613 -6188 34740 -6172
rect 34613 -6252 34660 -6188
rect 34724 -6252 34740 -6188
rect 34613 -6268 34740 -6252
rect 34613 -6332 34660 -6268
rect 34724 -6332 34740 -6268
rect 34613 -6348 34740 -6332
rect 34613 -6412 34660 -6348
rect 34724 -6412 34740 -6348
rect 34613 -6428 34740 -6412
rect 34613 -6492 34660 -6428
rect 34724 -6492 34740 -6428
rect 34613 -6508 34740 -6492
rect 34613 -6572 34660 -6508
rect 34724 -6572 34740 -6508
rect 34613 -6588 34740 -6572
rect 34613 -6652 34660 -6588
rect 34724 -6652 34740 -6588
rect 34613 -6668 34740 -6652
rect 34613 -6732 34660 -6668
rect 34724 -6732 34740 -6668
rect 34613 -6748 34740 -6732
rect 34613 -6812 34660 -6748
rect 34724 -6812 34740 -6748
rect 34613 -6828 34740 -6812
rect 34613 -6892 34660 -6828
rect 34724 -6892 34740 -6828
rect 34613 -6908 34740 -6892
rect 34613 -6972 34660 -6908
rect 34724 -6972 34740 -6908
rect 34613 -6988 34740 -6972
rect 34613 -7052 34660 -6988
rect 34724 -7052 34740 -6988
rect 34613 -7068 34740 -7052
rect 34613 -7132 34660 -7068
rect 34724 -7132 34740 -7068
rect 34613 -7148 34740 -7132
rect 34613 -7212 34660 -7148
rect 34724 -7212 34740 -7148
rect 34613 -7228 34740 -7212
rect 34613 -7292 34660 -7228
rect 34724 -7292 34740 -7228
rect 34613 -7308 34740 -7292
rect 34613 -7372 34660 -7308
rect 34724 -7372 34740 -7308
rect 34613 -7388 34740 -7372
rect 34613 -7452 34660 -7388
rect 34724 -7452 34740 -7388
rect 34613 -7468 34740 -7452
rect 34613 -7532 34660 -7468
rect 34724 -7532 34740 -7468
rect 34613 -7548 34740 -7532
rect 34613 -7612 34660 -7548
rect 34724 -7612 34740 -7548
rect 34613 -7628 34740 -7612
rect 34613 -7692 34660 -7628
rect 34724 -7692 34740 -7628
rect 34613 -7708 34740 -7692
rect 34613 -7772 34660 -7708
rect 34724 -7772 34740 -7708
rect 34613 -7788 34740 -7772
rect 34613 -7852 34660 -7788
rect 34724 -7852 34740 -7788
rect 34613 -7868 34740 -7852
rect 34613 -7932 34660 -7868
rect 34724 -7932 34740 -7868
rect 34613 -7948 34740 -7932
rect 34613 -8012 34660 -7948
rect 34724 -8012 34740 -7948
rect 34613 -8028 34740 -8012
rect 34613 -8092 34660 -8028
rect 34724 -8092 34740 -8028
rect 34613 -8108 34740 -8092
rect 34613 -8172 34660 -8108
rect 34724 -8172 34740 -8108
rect 34613 -8188 34740 -8172
rect 34613 -8252 34660 -8188
rect 34724 -8252 34740 -8188
rect 34613 -8268 34740 -8252
rect 34613 -8332 34660 -8268
rect 34724 -8332 34740 -8268
rect 34613 -8348 34740 -8332
rect 34613 -8412 34660 -8348
rect 34724 -8412 34740 -8348
rect 34613 -8428 34740 -8412
rect 34613 -8492 34660 -8428
rect 34724 -8492 34740 -8428
rect 34613 -8508 34740 -8492
rect 34613 -8572 34660 -8508
rect 34724 -8572 34740 -8508
rect 34613 -8588 34740 -8572
rect 34613 -8652 34660 -8588
rect 34724 -8652 34740 -8588
rect 34613 -8668 34740 -8652
rect 34613 -8732 34660 -8668
rect 34724 -8732 34740 -8668
rect 34613 -8748 34740 -8732
rect 34613 -8812 34660 -8748
rect 34724 -8812 34740 -8748
rect 34613 -8828 34740 -8812
rect 34613 -8892 34660 -8828
rect 34724 -8892 34740 -8828
rect 34613 -8908 34740 -8892
rect 34613 -8972 34660 -8908
rect 34724 -8972 34740 -8908
rect 34613 -8988 34740 -8972
rect 34613 -9052 34660 -8988
rect 34724 -9052 34740 -8988
rect 34613 -9068 34740 -9052
rect 34613 -9132 34660 -9068
rect 34724 -9132 34740 -9068
rect 34613 -9148 34740 -9132
rect 34613 -9212 34660 -9148
rect 34724 -9212 34740 -9148
rect 34613 -9228 34740 -9212
rect 28294 -9308 28421 -9292
rect 28294 -9372 28341 -9308
rect 28405 -9372 28421 -9308
rect 28294 -9388 28421 -9372
rect 28294 -9512 28398 -9388
rect 28294 -9528 28421 -9512
rect 28294 -9592 28341 -9528
rect 28405 -9592 28421 -9528
rect 28294 -9608 28421 -9592
rect 21975 -9688 22102 -9672
rect 21975 -9752 22022 -9688
rect 22086 -9752 22102 -9688
rect 21975 -9768 22102 -9752
rect 21975 -9832 22022 -9768
rect 22086 -9832 22102 -9768
rect 21975 -9848 22102 -9832
rect 21975 -9912 22022 -9848
rect 22086 -9912 22102 -9848
rect 21975 -9928 22102 -9912
rect 21975 -9992 22022 -9928
rect 22086 -9992 22102 -9928
rect 21975 -10008 22102 -9992
rect 21975 -10072 22022 -10008
rect 22086 -10072 22102 -10008
rect 21975 -10088 22102 -10072
rect 21975 -10152 22022 -10088
rect 22086 -10152 22102 -10088
rect 21975 -10168 22102 -10152
rect 21975 -10232 22022 -10168
rect 22086 -10232 22102 -10168
rect 21975 -10248 22102 -10232
rect 21975 -10312 22022 -10248
rect 22086 -10312 22102 -10248
rect 21975 -10328 22102 -10312
rect 21975 -10392 22022 -10328
rect 22086 -10392 22102 -10328
rect 21975 -10408 22102 -10392
rect 21975 -10472 22022 -10408
rect 22086 -10472 22102 -10408
rect 21975 -10488 22102 -10472
rect 21975 -10552 22022 -10488
rect 22086 -10552 22102 -10488
rect 21975 -10568 22102 -10552
rect 21975 -10632 22022 -10568
rect 22086 -10632 22102 -10568
rect 21975 -10648 22102 -10632
rect 21975 -10712 22022 -10648
rect 22086 -10712 22102 -10648
rect 21975 -10728 22102 -10712
rect 21975 -10792 22022 -10728
rect 22086 -10792 22102 -10728
rect 21975 -10808 22102 -10792
rect 21975 -10872 22022 -10808
rect 22086 -10872 22102 -10808
rect 21975 -10888 22102 -10872
rect 21975 -10952 22022 -10888
rect 22086 -10952 22102 -10888
rect 21975 -10968 22102 -10952
rect 21975 -11032 22022 -10968
rect 22086 -11032 22102 -10968
rect 21975 -11048 22102 -11032
rect 21975 -11112 22022 -11048
rect 22086 -11112 22102 -11048
rect 21975 -11128 22102 -11112
rect 21975 -11192 22022 -11128
rect 22086 -11192 22102 -11128
rect 21975 -11208 22102 -11192
rect 21975 -11272 22022 -11208
rect 22086 -11272 22102 -11208
rect 21975 -11288 22102 -11272
rect 21975 -11352 22022 -11288
rect 22086 -11352 22102 -11288
rect 21975 -11368 22102 -11352
rect 21975 -11432 22022 -11368
rect 22086 -11432 22102 -11368
rect 21975 -11448 22102 -11432
rect 21975 -11512 22022 -11448
rect 22086 -11512 22102 -11448
rect 21975 -11528 22102 -11512
rect 21975 -11592 22022 -11528
rect 22086 -11592 22102 -11528
rect 21975 -11608 22102 -11592
rect 21975 -11672 22022 -11608
rect 22086 -11672 22102 -11608
rect 21975 -11688 22102 -11672
rect 21975 -11752 22022 -11688
rect 22086 -11752 22102 -11688
rect 21975 -11768 22102 -11752
rect 21975 -11832 22022 -11768
rect 22086 -11832 22102 -11768
rect 21975 -11848 22102 -11832
rect 21975 -11912 22022 -11848
rect 22086 -11912 22102 -11848
rect 21975 -11928 22102 -11912
rect 21975 -11992 22022 -11928
rect 22086 -11992 22102 -11928
rect 21975 -12008 22102 -11992
rect 21975 -12072 22022 -12008
rect 22086 -12072 22102 -12008
rect 21975 -12088 22102 -12072
rect 21975 -12152 22022 -12088
rect 22086 -12152 22102 -12088
rect 21975 -12168 22102 -12152
rect 21975 -12232 22022 -12168
rect 22086 -12232 22102 -12168
rect 21975 -12248 22102 -12232
rect 21975 -12312 22022 -12248
rect 22086 -12312 22102 -12248
rect 21975 -12328 22102 -12312
rect 21975 -12392 22022 -12328
rect 22086 -12392 22102 -12328
rect 21975 -12408 22102 -12392
rect 21975 -12472 22022 -12408
rect 22086 -12472 22102 -12408
rect 21975 -12488 22102 -12472
rect 21975 -12552 22022 -12488
rect 22086 -12552 22102 -12488
rect 21975 -12568 22102 -12552
rect 21975 -12632 22022 -12568
rect 22086 -12632 22102 -12568
rect 21975 -12648 22102 -12632
rect 21975 -12712 22022 -12648
rect 22086 -12712 22102 -12648
rect 21975 -12728 22102 -12712
rect 21975 -12792 22022 -12728
rect 22086 -12792 22102 -12728
rect 21975 -12808 22102 -12792
rect 21975 -12872 22022 -12808
rect 22086 -12872 22102 -12808
rect 21975 -12888 22102 -12872
rect 21975 -12952 22022 -12888
rect 22086 -12952 22102 -12888
rect 21975 -12968 22102 -12952
rect 21975 -13032 22022 -12968
rect 22086 -13032 22102 -12968
rect 21975 -13048 22102 -13032
rect 21975 -13112 22022 -13048
rect 22086 -13112 22102 -13048
rect 21975 -13128 22102 -13112
rect 21975 -13192 22022 -13128
rect 22086 -13192 22102 -13128
rect 21975 -13208 22102 -13192
rect 21975 -13272 22022 -13208
rect 22086 -13272 22102 -13208
rect 21975 -13288 22102 -13272
rect 21975 -13352 22022 -13288
rect 22086 -13352 22102 -13288
rect 21975 -13368 22102 -13352
rect 21975 -13432 22022 -13368
rect 22086 -13432 22102 -13368
rect 21975 -13448 22102 -13432
rect 21975 -13512 22022 -13448
rect 22086 -13512 22102 -13448
rect 21975 -13528 22102 -13512
rect 21975 -13592 22022 -13528
rect 22086 -13592 22102 -13528
rect 21975 -13608 22102 -13592
rect 21975 -13672 22022 -13608
rect 22086 -13672 22102 -13608
rect 21975 -13688 22102 -13672
rect 21975 -13752 22022 -13688
rect 22086 -13752 22102 -13688
rect 21975 -13768 22102 -13752
rect 21975 -13832 22022 -13768
rect 22086 -13832 22102 -13768
rect 21975 -13848 22102 -13832
rect 21975 -13912 22022 -13848
rect 22086 -13912 22102 -13848
rect 21975 -13928 22102 -13912
rect 21975 -13992 22022 -13928
rect 22086 -13992 22102 -13928
rect 21975 -14008 22102 -13992
rect 21975 -14072 22022 -14008
rect 22086 -14072 22102 -14008
rect 21975 -14088 22102 -14072
rect 21975 -14152 22022 -14088
rect 22086 -14152 22102 -14088
rect 21975 -14168 22102 -14152
rect 21975 -14232 22022 -14168
rect 22086 -14232 22102 -14168
rect 21975 -14248 22102 -14232
rect 21975 -14312 22022 -14248
rect 22086 -14312 22102 -14248
rect 21975 -14328 22102 -14312
rect 21975 -14392 22022 -14328
rect 22086 -14392 22102 -14328
rect 21975 -14408 22102 -14392
rect 21975 -14472 22022 -14408
rect 22086 -14472 22102 -14408
rect 21975 -14488 22102 -14472
rect 21975 -14552 22022 -14488
rect 22086 -14552 22102 -14488
rect 21975 -14568 22102 -14552
rect 21975 -14632 22022 -14568
rect 22086 -14632 22102 -14568
rect 21975 -14648 22102 -14632
rect 21975 -14712 22022 -14648
rect 22086 -14712 22102 -14648
rect 21975 -14728 22102 -14712
rect 21975 -14792 22022 -14728
rect 22086 -14792 22102 -14728
rect 21975 -14808 22102 -14792
rect 21975 -14872 22022 -14808
rect 22086 -14872 22102 -14808
rect 21975 -14888 22102 -14872
rect 21975 -14952 22022 -14888
rect 22086 -14952 22102 -14888
rect 21975 -14968 22102 -14952
rect 21975 -15032 22022 -14968
rect 22086 -15032 22102 -14968
rect 21975 -15048 22102 -15032
rect 21975 -15112 22022 -15048
rect 22086 -15112 22102 -15048
rect 21975 -15128 22102 -15112
rect 21975 -15192 22022 -15128
rect 22086 -15192 22102 -15128
rect 21975 -15208 22102 -15192
rect 21975 -15272 22022 -15208
rect 22086 -15272 22102 -15208
rect 21975 -15288 22102 -15272
rect 21975 -15352 22022 -15288
rect 22086 -15352 22102 -15288
rect 21975 -15368 22102 -15352
rect 21975 -15432 22022 -15368
rect 22086 -15432 22102 -15368
rect 21975 -15448 22102 -15432
rect 21975 -15512 22022 -15448
rect 22086 -15512 22102 -15448
rect 21975 -15528 22102 -15512
rect 15656 -15608 15783 -15592
rect 15656 -15672 15703 -15608
rect 15767 -15672 15783 -15608
rect 15656 -15688 15783 -15672
rect 15656 -15812 15760 -15688
rect 15656 -15828 15783 -15812
rect 15656 -15892 15703 -15828
rect 15767 -15892 15783 -15828
rect 15656 -15908 15783 -15892
rect 9337 -15988 9464 -15972
rect 9337 -16052 9384 -15988
rect 9448 -16052 9464 -15988
rect 9337 -16068 9464 -16052
rect 9337 -16132 9384 -16068
rect 9448 -16132 9464 -16068
rect 9337 -16148 9464 -16132
rect 9337 -16212 9384 -16148
rect 9448 -16212 9464 -16148
rect 9337 -16228 9464 -16212
rect 9337 -16292 9384 -16228
rect 9448 -16292 9464 -16228
rect 9337 -16308 9464 -16292
rect 9337 -16372 9384 -16308
rect 9448 -16372 9464 -16308
rect 9337 -16388 9464 -16372
rect 9337 -16452 9384 -16388
rect 9448 -16452 9464 -16388
rect 9337 -16468 9464 -16452
rect 9337 -16532 9384 -16468
rect 9448 -16532 9464 -16468
rect 9337 -16548 9464 -16532
rect 9337 -16612 9384 -16548
rect 9448 -16612 9464 -16548
rect 9337 -16628 9464 -16612
rect 9337 -16692 9384 -16628
rect 9448 -16692 9464 -16628
rect 9337 -16708 9464 -16692
rect 9337 -16772 9384 -16708
rect 9448 -16772 9464 -16708
rect 9337 -16788 9464 -16772
rect 9337 -16852 9384 -16788
rect 9448 -16852 9464 -16788
rect 9337 -16868 9464 -16852
rect 9337 -16932 9384 -16868
rect 9448 -16932 9464 -16868
rect 9337 -16948 9464 -16932
rect 9337 -17012 9384 -16948
rect 9448 -17012 9464 -16948
rect 9337 -17028 9464 -17012
rect 9337 -17092 9384 -17028
rect 9448 -17092 9464 -17028
rect 9337 -17108 9464 -17092
rect 9337 -17172 9384 -17108
rect 9448 -17172 9464 -17108
rect 9337 -17188 9464 -17172
rect 9337 -17252 9384 -17188
rect 9448 -17252 9464 -17188
rect 9337 -17268 9464 -17252
rect 9337 -17332 9384 -17268
rect 9448 -17332 9464 -17268
rect 9337 -17348 9464 -17332
rect 9337 -17412 9384 -17348
rect 9448 -17412 9464 -17348
rect 9337 -17428 9464 -17412
rect 9337 -17492 9384 -17428
rect 9448 -17492 9464 -17428
rect 9337 -17508 9464 -17492
rect 9337 -17572 9384 -17508
rect 9448 -17572 9464 -17508
rect 9337 -17588 9464 -17572
rect 9337 -17652 9384 -17588
rect 9448 -17652 9464 -17588
rect 9337 -17668 9464 -17652
rect 9337 -17732 9384 -17668
rect 9448 -17732 9464 -17668
rect 9337 -17748 9464 -17732
rect 9337 -17812 9384 -17748
rect 9448 -17812 9464 -17748
rect 9337 -17828 9464 -17812
rect 9337 -17892 9384 -17828
rect 9448 -17892 9464 -17828
rect 9337 -17908 9464 -17892
rect 9337 -17972 9384 -17908
rect 9448 -17972 9464 -17908
rect 9337 -17988 9464 -17972
rect 9337 -18052 9384 -17988
rect 9448 -18052 9464 -17988
rect 9337 -18068 9464 -18052
rect 9337 -18132 9384 -18068
rect 9448 -18132 9464 -18068
rect 9337 -18148 9464 -18132
rect 9337 -18212 9384 -18148
rect 9448 -18212 9464 -18148
rect 9337 -18228 9464 -18212
rect 9337 -18292 9384 -18228
rect 9448 -18292 9464 -18228
rect 9337 -18308 9464 -18292
rect 9337 -18372 9384 -18308
rect 9448 -18372 9464 -18308
rect 9337 -18388 9464 -18372
rect 9337 -18452 9384 -18388
rect 9448 -18452 9464 -18388
rect 9337 -18468 9464 -18452
rect 9337 -18532 9384 -18468
rect 9448 -18532 9464 -18468
rect 9337 -18548 9464 -18532
rect 9337 -18612 9384 -18548
rect 9448 -18612 9464 -18548
rect 9337 -18628 9464 -18612
rect 9337 -18692 9384 -18628
rect 9448 -18692 9464 -18628
rect 9337 -18708 9464 -18692
rect 9337 -18772 9384 -18708
rect 9448 -18772 9464 -18708
rect 9337 -18788 9464 -18772
rect 9337 -18852 9384 -18788
rect 9448 -18852 9464 -18788
rect 9337 -18868 9464 -18852
rect 9337 -18932 9384 -18868
rect 9448 -18932 9464 -18868
rect 9337 -18948 9464 -18932
rect 9337 -19012 9384 -18948
rect 9448 -19012 9464 -18948
rect 9337 -19028 9464 -19012
rect 9337 -19092 9384 -19028
rect 9448 -19092 9464 -19028
rect 9337 -19108 9464 -19092
rect 9337 -19172 9384 -19108
rect 9448 -19172 9464 -19108
rect 9337 -19188 9464 -19172
rect 9337 -19252 9384 -19188
rect 9448 -19252 9464 -19188
rect 9337 -19268 9464 -19252
rect 9337 -19332 9384 -19268
rect 9448 -19332 9464 -19268
rect 9337 -19348 9464 -19332
rect 9337 -19412 9384 -19348
rect 9448 -19412 9464 -19348
rect 9337 -19428 9464 -19412
rect 9337 -19492 9384 -19428
rect 9448 -19492 9464 -19428
rect 9337 -19508 9464 -19492
rect 9337 -19572 9384 -19508
rect 9448 -19572 9464 -19508
rect 9337 -19588 9464 -19572
rect 9337 -19652 9384 -19588
rect 9448 -19652 9464 -19588
rect 9337 -19668 9464 -19652
rect 9337 -19732 9384 -19668
rect 9448 -19732 9464 -19668
rect 9337 -19748 9464 -19732
rect 9337 -19812 9384 -19748
rect 9448 -19812 9464 -19748
rect 9337 -19828 9464 -19812
rect 9337 -19892 9384 -19828
rect 9448 -19892 9464 -19828
rect 9337 -19908 9464 -19892
rect 9337 -19972 9384 -19908
rect 9448 -19972 9464 -19908
rect 9337 -19988 9464 -19972
rect 9337 -20052 9384 -19988
rect 9448 -20052 9464 -19988
rect 9337 -20068 9464 -20052
rect 9337 -20132 9384 -20068
rect 9448 -20132 9464 -20068
rect 9337 -20148 9464 -20132
rect 9337 -20212 9384 -20148
rect 9448 -20212 9464 -20148
rect 9337 -20228 9464 -20212
rect 9337 -20292 9384 -20228
rect 9448 -20292 9464 -20228
rect 9337 -20308 9464 -20292
rect 9337 -20372 9384 -20308
rect 9448 -20372 9464 -20308
rect 9337 -20388 9464 -20372
rect 9337 -20452 9384 -20388
rect 9448 -20452 9464 -20388
rect 9337 -20468 9464 -20452
rect 9337 -20532 9384 -20468
rect 9448 -20532 9464 -20468
rect 9337 -20548 9464 -20532
rect 9337 -20612 9384 -20548
rect 9448 -20612 9464 -20548
rect 9337 -20628 9464 -20612
rect 9337 -20692 9384 -20628
rect 9448 -20692 9464 -20628
rect 9337 -20708 9464 -20692
rect 9337 -20772 9384 -20708
rect 9448 -20772 9464 -20708
rect 9337 -20788 9464 -20772
rect 9337 -20852 9384 -20788
rect 9448 -20852 9464 -20788
rect 9337 -20868 9464 -20852
rect 9337 -20932 9384 -20868
rect 9448 -20932 9464 -20868
rect 9337 -20948 9464 -20932
rect 9337 -21012 9384 -20948
rect 9448 -21012 9464 -20948
rect 9337 -21028 9464 -21012
rect 9337 -21092 9384 -21028
rect 9448 -21092 9464 -21028
rect 9337 -21108 9464 -21092
rect 9337 -21172 9384 -21108
rect 9448 -21172 9464 -21108
rect 9337 -21188 9464 -21172
rect 9337 -21252 9384 -21188
rect 9448 -21252 9464 -21188
rect 9337 -21268 9464 -21252
rect 9337 -21332 9384 -21268
rect 9448 -21332 9464 -21268
rect 9337 -21348 9464 -21332
rect 9337 -21412 9384 -21348
rect 9448 -21412 9464 -21348
rect 9337 -21428 9464 -21412
rect 9337 -21492 9384 -21428
rect 9448 -21492 9464 -21428
rect 9337 -21508 9464 -21492
rect 9337 -21572 9384 -21508
rect 9448 -21572 9464 -21508
rect 9337 -21588 9464 -21572
rect 9337 -21652 9384 -21588
rect 9448 -21652 9464 -21588
rect 9337 -21668 9464 -21652
rect 9337 -21732 9384 -21668
rect 9448 -21732 9464 -21668
rect 9337 -21748 9464 -21732
rect 9337 -21812 9384 -21748
rect 9448 -21812 9464 -21748
rect 9337 -21828 9464 -21812
rect 3018 -21908 3145 -21892
rect 3018 -21972 3065 -21908
rect 3129 -21972 3145 -21908
rect 3018 -21988 3145 -21972
rect 3018 -22112 3122 -21988
rect 3018 -22128 3145 -22112
rect 3018 -22192 3065 -22128
rect 3129 -22192 3145 -22128
rect 3018 -22208 3145 -22192
rect -3301 -22288 -3174 -22272
rect -3301 -22352 -3254 -22288
rect -3190 -22352 -3174 -22288
rect -3301 -22368 -3174 -22352
rect -3301 -22432 -3254 -22368
rect -3190 -22432 -3174 -22368
rect -3301 -22448 -3174 -22432
rect -3301 -22512 -3254 -22448
rect -3190 -22512 -3174 -22448
rect -3301 -22528 -3174 -22512
rect -3301 -22592 -3254 -22528
rect -3190 -22592 -3174 -22528
rect -3301 -22608 -3174 -22592
rect -3301 -22672 -3254 -22608
rect -3190 -22672 -3174 -22608
rect -3301 -22688 -3174 -22672
rect -3301 -22752 -3254 -22688
rect -3190 -22752 -3174 -22688
rect -3301 -22768 -3174 -22752
rect -3301 -22832 -3254 -22768
rect -3190 -22832 -3174 -22768
rect -3301 -22848 -3174 -22832
rect -3301 -22912 -3254 -22848
rect -3190 -22912 -3174 -22848
rect -3301 -22928 -3174 -22912
rect -3301 -22992 -3254 -22928
rect -3190 -22992 -3174 -22928
rect -3301 -23008 -3174 -22992
rect -3301 -23072 -3254 -23008
rect -3190 -23072 -3174 -23008
rect -3301 -23088 -3174 -23072
rect -3301 -23152 -3254 -23088
rect -3190 -23152 -3174 -23088
rect -3301 -23168 -3174 -23152
rect -3301 -23232 -3254 -23168
rect -3190 -23232 -3174 -23168
rect -3301 -23248 -3174 -23232
rect -3301 -23312 -3254 -23248
rect -3190 -23312 -3174 -23248
rect -3301 -23328 -3174 -23312
rect -3301 -23392 -3254 -23328
rect -3190 -23392 -3174 -23328
rect -3301 -23408 -3174 -23392
rect -3301 -23472 -3254 -23408
rect -3190 -23472 -3174 -23408
rect -3301 -23488 -3174 -23472
rect -3301 -23552 -3254 -23488
rect -3190 -23552 -3174 -23488
rect -3301 -23568 -3174 -23552
rect -3301 -23632 -3254 -23568
rect -3190 -23632 -3174 -23568
rect -3301 -23648 -3174 -23632
rect -3301 -23712 -3254 -23648
rect -3190 -23712 -3174 -23648
rect -3301 -23728 -3174 -23712
rect -3301 -23792 -3254 -23728
rect -3190 -23792 -3174 -23728
rect -3301 -23808 -3174 -23792
rect -3301 -23872 -3254 -23808
rect -3190 -23872 -3174 -23808
rect -3301 -23888 -3174 -23872
rect -3301 -23952 -3254 -23888
rect -3190 -23952 -3174 -23888
rect -3301 -23968 -3174 -23952
rect -3301 -24032 -3254 -23968
rect -3190 -24032 -3174 -23968
rect -3301 -24048 -3174 -24032
rect -3301 -24112 -3254 -24048
rect -3190 -24112 -3174 -24048
rect -3301 -24128 -3174 -24112
rect -3301 -24192 -3254 -24128
rect -3190 -24192 -3174 -24128
rect -3301 -24208 -3174 -24192
rect -3301 -24272 -3254 -24208
rect -3190 -24272 -3174 -24208
rect -3301 -24288 -3174 -24272
rect -3301 -24352 -3254 -24288
rect -3190 -24352 -3174 -24288
rect -3301 -24368 -3174 -24352
rect -3301 -24432 -3254 -24368
rect -3190 -24432 -3174 -24368
rect -3301 -24448 -3174 -24432
rect -3301 -24512 -3254 -24448
rect -3190 -24512 -3174 -24448
rect -3301 -24528 -3174 -24512
rect -3301 -24592 -3254 -24528
rect -3190 -24592 -3174 -24528
rect -3301 -24608 -3174 -24592
rect -3301 -24672 -3254 -24608
rect -3190 -24672 -3174 -24608
rect -3301 -24688 -3174 -24672
rect -3301 -24752 -3254 -24688
rect -3190 -24752 -3174 -24688
rect -3301 -24768 -3174 -24752
rect -3301 -24832 -3254 -24768
rect -3190 -24832 -3174 -24768
rect -3301 -24848 -3174 -24832
rect -3301 -24912 -3254 -24848
rect -3190 -24912 -3174 -24848
rect -3301 -24928 -3174 -24912
rect -3301 -24992 -3254 -24928
rect -3190 -24992 -3174 -24928
rect -3301 -25008 -3174 -24992
rect -3301 -25072 -3254 -25008
rect -3190 -25072 -3174 -25008
rect -3301 -25088 -3174 -25072
rect -3301 -25152 -3254 -25088
rect -3190 -25152 -3174 -25088
rect -3301 -25168 -3174 -25152
rect -3301 -25232 -3254 -25168
rect -3190 -25232 -3174 -25168
rect -3301 -25248 -3174 -25232
rect -3301 -25312 -3254 -25248
rect -3190 -25312 -3174 -25248
rect -3301 -25328 -3174 -25312
rect -3301 -25392 -3254 -25328
rect -3190 -25392 -3174 -25328
rect -3301 -25408 -3174 -25392
rect -3301 -25472 -3254 -25408
rect -3190 -25472 -3174 -25408
rect -3301 -25488 -3174 -25472
rect -3301 -25552 -3254 -25488
rect -3190 -25552 -3174 -25488
rect -3301 -25568 -3174 -25552
rect -3301 -25632 -3254 -25568
rect -3190 -25632 -3174 -25568
rect -3301 -25648 -3174 -25632
rect -3301 -25712 -3254 -25648
rect -3190 -25712 -3174 -25648
rect -3301 -25728 -3174 -25712
rect -3301 -25792 -3254 -25728
rect -3190 -25792 -3174 -25728
rect -3301 -25808 -3174 -25792
rect -3301 -25872 -3254 -25808
rect -3190 -25872 -3174 -25808
rect -3301 -25888 -3174 -25872
rect -3301 -25952 -3254 -25888
rect -3190 -25952 -3174 -25888
rect -3301 -25968 -3174 -25952
rect -3301 -26032 -3254 -25968
rect -3190 -26032 -3174 -25968
rect -3301 -26048 -3174 -26032
rect -3301 -26112 -3254 -26048
rect -3190 -26112 -3174 -26048
rect -3301 -26128 -3174 -26112
rect -3301 -26192 -3254 -26128
rect -3190 -26192 -3174 -26128
rect -3301 -26208 -3174 -26192
rect -3301 -26272 -3254 -26208
rect -3190 -26272 -3174 -26208
rect -3301 -26288 -3174 -26272
rect -3301 -26352 -3254 -26288
rect -3190 -26352 -3174 -26288
rect -3301 -26368 -3174 -26352
rect -3301 -26432 -3254 -26368
rect -3190 -26432 -3174 -26368
rect -3301 -26448 -3174 -26432
rect -3301 -26512 -3254 -26448
rect -3190 -26512 -3174 -26448
rect -3301 -26528 -3174 -26512
rect -3301 -26592 -3254 -26528
rect -3190 -26592 -3174 -26528
rect -3301 -26608 -3174 -26592
rect -3301 -26672 -3254 -26608
rect -3190 -26672 -3174 -26608
rect -3301 -26688 -3174 -26672
rect -3301 -26752 -3254 -26688
rect -3190 -26752 -3174 -26688
rect -3301 -26768 -3174 -26752
rect -3301 -26832 -3254 -26768
rect -3190 -26832 -3174 -26768
rect -3301 -26848 -3174 -26832
rect -3301 -26912 -3254 -26848
rect -3190 -26912 -3174 -26848
rect -3301 -26928 -3174 -26912
rect -3301 -26992 -3254 -26928
rect -3190 -26992 -3174 -26928
rect -3301 -27008 -3174 -26992
rect -3301 -27072 -3254 -27008
rect -3190 -27072 -3174 -27008
rect -3301 -27088 -3174 -27072
rect -3301 -27152 -3254 -27088
rect -3190 -27152 -3174 -27088
rect -3301 -27168 -3174 -27152
rect -3301 -27232 -3254 -27168
rect -3190 -27232 -3174 -27168
rect -3301 -27248 -3174 -27232
rect -3301 -27312 -3254 -27248
rect -3190 -27312 -3174 -27248
rect -3301 -27328 -3174 -27312
rect -3301 -27392 -3254 -27328
rect -3190 -27392 -3174 -27328
rect -3301 -27408 -3174 -27392
rect -3301 -27472 -3254 -27408
rect -3190 -27472 -3174 -27408
rect -3301 -27488 -3174 -27472
rect -3301 -27552 -3254 -27488
rect -3190 -27552 -3174 -27488
rect -3301 -27568 -3174 -27552
rect -3301 -27632 -3254 -27568
rect -3190 -27632 -3174 -27568
rect -3301 -27648 -3174 -27632
rect -3301 -27712 -3254 -27648
rect -3190 -27712 -3174 -27648
rect -3301 -27728 -3174 -27712
rect -3301 -27792 -3254 -27728
rect -3190 -27792 -3174 -27728
rect -3301 -27808 -3174 -27792
rect -3301 -27872 -3254 -27808
rect -3190 -27872 -3174 -27808
rect -3301 -27888 -3174 -27872
rect -3301 -27952 -3254 -27888
rect -3190 -27952 -3174 -27888
rect -3301 -27968 -3174 -27952
rect -3301 -28032 -3254 -27968
rect -3190 -28032 -3174 -27968
rect -3301 -28048 -3174 -28032
rect -3301 -28112 -3254 -28048
rect -3190 -28112 -3174 -28048
rect -3301 -28128 -3174 -28112
rect -9620 -28208 -9493 -28192
rect -9620 -28272 -9573 -28208
rect -9509 -28272 -9493 -28208
rect -9620 -28288 -9493 -28272
rect -9620 -28412 -9516 -28288
rect -9620 -28428 -9493 -28412
rect -9620 -28492 -9573 -28428
rect -9509 -28492 -9493 -28428
rect -9620 -28508 -9493 -28492
rect -15939 -28588 -15812 -28572
rect -15939 -28652 -15892 -28588
rect -15828 -28652 -15812 -28588
rect -15939 -28668 -15812 -28652
rect -15939 -28732 -15892 -28668
rect -15828 -28732 -15812 -28668
rect -15939 -28748 -15812 -28732
rect -15939 -28812 -15892 -28748
rect -15828 -28812 -15812 -28748
rect -15939 -28828 -15812 -28812
rect -15939 -28892 -15892 -28828
rect -15828 -28892 -15812 -28828
rect -15939 -28908 -15812 -28892
rect -15939 -28972 -15892 -28908
rect -15828 -28972 -15812 -28908
rect -15939 -28988 -15812 -28972
rect -15939 -29052 -15892 -28988
rect -15828 -29052 -15812 -28988
rect -15939 -29068 -15812 -29052
rect -15939 -29132 -15892 -29068
rect -15828 -29132 -15812 -29068
rect -15939 -29148 -15812 -29132
rect -15939 -29212 -15892 -29148
rect -15828 -29212 -15812 -29148
rect -15939 -29228 -15812 -29212
rect -15939 -29292 -15892 -29228
rect -15828 -29292 -15812 -29228
rect -15939 -29308 -15812 -29292
rect -15939 -29372 -15892 -29308
rect -15828 -29372 -15812 -29308
rect -15939 -29388 -15812 -29372
rect -15939 -29452 -15892 -29388
rect -15828 -29452 -15812 -29388
rect -15939 -29468 -15812 -29452
rect -15939 -29532 -15892 -29468
rect -15828 -29532 -15812 -29468
rect -15939 -29548 -15812 -29532
rect -15939 -29612 -15892 -29548
rect -15828 -29612 -15812 -29548
rect -15939 -29628 -15812 -29612
rect -15939 -29692 -15892 -29628
rect -15828 -29692 -15812 -29628
rect -15939 -29708 -15812 -29692
rect -15939 -29772 -15892 -29708
rect -15828 -29772 -15812 -29708
rect -15939 -29788 -15812 -29772
rect -15939 -29852 -15892 -29788
rect -15828 -29852 -15812 -29788
rect -15939 -29868 -15812 -29852
rect -15939 -29932 -15892 -29868
rect -15828 -29932 -15812 -29868
rect -15939 -29948 -15812 -29932
rect -15939 -30012 -15892 -29948
rect -15828 -30012 -15812 -29948
rect -15939 -30028 -15812 -30012
rect -15939 -30092 -15892 -30028
rect -15828 -30092 -15812 -30028
rect -15939 -30108 -15812 -30092
rect -15939 -30172 -15892 -30108
rect -15828 -30172 -15812 -30108
rect -15939 -30188 -15812 -30172
rect -15939 -30252 -15892 -30188
rect -15828 -30252 -15812 -30188
rect -15939 -30268 -15812 -30252
rect -15939 -30332 -15892 -30268
rect -15828 -30332 -15812 -30268
rect -15939 -30348 -15812 -30332
rect -15939 -30412 -15892 -30348
rect -15828 -30412 -15812 -30348
rect -15939 -30428 -15812 -30412
rect -15939 -30492 -15892 -30428
rect -15828 -30492 -15812 -30428
rect -15939 -30508 -15812 -30492
rect -15939 -30572 -15892 -30508
rect -15828 -30572 -15812 -30508
rect -15939 -30588 -15812 -30572
rect -15939 -30652 -15892 -30588
rect -15828 -30652 -15812 -30588
rect -15939 -30668 -15812 -30652
rect -15939 -30732 -15892 -30668
rect -15828 -30732 -15812 -30668
rect -15939 -30748 -15812 -30732
rect -15939 -30812 -15892 -30748
rect -15828 -30812 -15812 -30748
rect -15939 -30828 -15812 -30812
rect -15939 -30892 -15892 -30828
rect -15828 -30892 -15812 -30828
rect -15939 -30908 -15812 -30892
rect -15939 -30972 -15892 -30908
rect -15828 -30972 -15812 -30908
rect -15939 -30988 -15812 -30972
rect -15939 -31052 -15892 -30988
rect -15828 -31052 -15812 -30988
rect -15939 -31068 -15812 -31052
rect -15939 -31132 -15892 -31068
rect -15828 -31132 -15812 -31068
rect -15939 -31148 -15812 -31132
rect -15939 -31212 -15892 -31148
rect -15828 -31212 -15812 -31148
rect -15939 -31228 -15812 -31212
rect -15939 -31292 -15892 -31228
rect -15828 -31292 -15812 -31228
rect -15939 -31308 -15812 -31292
rect -15939 -31372 -15892 -31308
rect -15828 -31372 -15812 -31308
rect -15939 -31388 -15812 -31372
rect -15939 -31452 -15892 -31388
rect -15828 -31452 -15812 -31388
rect -15939 -31468 -15812 -31452
rect -15939 -31532 -15892 -31468
rect -15828 -31532 -15812 -31468
rect -15939 -31548 -15812 -31532
rect -15939 -31612 -15892 -31548
rect -15828 -31612 -15812 -31548
rect -15939 -31628 -15812 -31612
rect -15939 -31692 -15892 -31628
rect -15828 -31692 -15812 -31628
rect -15939 -31708 -15812 -31692
rect -15939 -31772 -15892 -31708
rect -15828 -31772 -15812 -31708
rect -15939 -31788 -15812 -31772
rect -15939 -31852 -15892 -31788
rect -15828 -31852 -15812 -31788
rect -15939 -31868 -15812 -31852
rect -15939 -31932 -15892 -31868
rect -15828 -31932 -15812 -31868
rect -15939 -31948 -15812 -31932
rect -15939 -32012 -15892 -31948
rect -15828 -32012 -15812 -31948
rect -15939 -32028 -15812 -32012
rect -15939 -32092 -15892 -32028
rect -15828 -32092 -15812 -32028
rect -15939 -32108 -15812 -32092
rect -15939 -32172 -15892 -32108
rect -15828 -32172 -15812 -32108
rect -15939 -32188 -15812 -32172
rect -15939 -32252 -15892 -32188
rect -15828 -32252 -15812 -32188
rect -15939 -32268 -15812 -32252
rect -15939 -32332 -15892 -32268
rect -15828 -32332 -15812 -32268
rect -15939 -32348 -15812 -32332
rect -15939 -32412 -15892 -32348
rect -15828 -32412 -15812 -32348
rect -15939 -32428 -15812 -32412
rect -15939 -32492 -15892 -32428
rect -15828 -32492 -15812 -32428
rect -15939 -32508 -15812 -32492
rect -15939 -32572 -15892 -32508
rect -15828 -32572 -15812 -32508
rect -15939 -32588 -15812 -32572
rect -15939 -32652 -15892 -32588
rect -15828 -32652 -15812 -32588
rect -15939 -32668 -15812 -32652
rect -15939 -32732 -15892 -32668
rect -15828 -32732 -15812 -32668
rect -15939 -32748 -15812 -32732
rect -15939 -32812 -15892 -32748
rect -15828 -32812 -15812 -32748
rect -15939 -32828 -15812 -32812
rect -15939 -32892 -15892 -32828
rect -15828 -32892 -15812 -32828
rect -15939 -32908 -15812 -32892
rect -15939 -32972 -15892 -32908
rect -15828 -32972 -15812 -32908
rect -15939 -32988 -15812 -32972
rect -15939 -33052 -15892 -32988
rect -15828 -33052 -15812 -32988
rect -15939 -33068 -15812 -33052
rect -15939 -33132 -15892 -33068
rect -15828 -33132 -15812 -33068
rect -15939 -33148 -15812 -33132
rect -15939 -33212 -15892 -33148
rect -15828 -33212 -15812 -33148
rect -15939 -33228 -15812 -33212
rect -15939 -33292 -15892 -33228
rect -15828 -33292 -15812 -33228
rect -15939 -33308 -15812 -33292
rect -15939 -33372 -15892 -33308
rect -15828 -33372 -15812 -33308
rect -15939 -33388 -15812 -33372
rect -15939 -33452 -15892 -33388
rect -15828 -33452 -15812 -33388
rect -15939 -33468 -15812 -33452
rect -15939 -33532 -15892 -33468
rect -15828 -33532 -15812 -33468
rect -15939 -33548 -15812 -33532
rect -15939 -33612 -15892 -33548
rect -15828 -33612 -15812 -33548
rect -15939 -33628 -15812 -33612
rect -15939 -33692 -15892 -33628
rect -15828 -33692 -15812 -33628
rect -15939 -33708 -15812 -33692
rect -15939 -33772 -15892 -33708
rect -15828 -33772 -15812 -33708
rect -15939 -33788 -15812 -33772
rect -15939 -33852 -15892 -33788
rect -15828 -33852 -15812 -33788
rect -15939 -33868 -15812 -33852
rect -15939 -33932 -15892 -33868
rect -15828 -33932 -15812 -33868
rect -15939 -33948 -15812 -33932
rect -15939 -34012 -15892 -33948
rect -15828 -34012 -15812 -33948
rect -15939 -34028 -15812 -34012
rect -15939 -34092 -15892 -34028
rect -15828 -34092 -15812 -34028
rect -15939 -34108 -15812 -34092
rect -15939 -34172 -15892 -34108
rect -15828 -34172 -15812 -34108
rect -15939 -34188 -15812 -34172
rect -15939 -34252 -15892 -34188
rect -15828 -34252 -15812 -34188
rect -15939 -34268 -15812 -34252
rect -15939 -34332 -15892 -34268
rect -15828 -34332 -15812 -34268
rect -15939 -34348 -15812 -34332
rect -15939 -34412 -15892 -34348
rect -15828 -34412 -15812 -34348
rect -15939 -34428 -15812 -34412
rect -22258 -34508 -22131 -34492
rect -22258 -34572 -22211 -34508
rect -22147 -34572 -22131 -34508
rect -22258 -34588 -22131 -34572
rect -22258 -34712 -22154 -34588
rect -22258 -34728 -22131 -34712
rect -22258 -34792 -22211 -34728
rect -22147 -34792 -22131 -34728
rect -22258 -34808 -22131 -34792
rect -28577 -34888 -28450 -34872
rect -28577 -34952 -28530 -34888
rect -28466 -34952 -28450 -34888
rect -28577 -34968 -28450 -34952
rect -28577 -35032 -28530 -34968
rect -28466 -35032 -28450 -34968
rect -28577 -35048 -28450 -35032
rect -28577 -35112 -28530 -35048
rect -28466 -35112 -28450 -35048
rect -28577 -35128 -28450 -35112
rect -28577 -35192 -28530 -35128
rect -28466 -35192 -28450 -35128
rect -28577 -35208 -28450 -35192
rect -28577 -35272 -28530 -35208
rect -28466 -35272 -28450 -35208
rect -28577 -35288 -28450 -35272
rect -28577 -35352 -28530 -35288
rect -28466 -35352 -28450 -35288
rect -28577 -35368 -28450 -35352
rect -28577 -35432 -28530 -35368
rect -28466 -35432 -28450 -35368
rect -28577 -35448 -28450 -35432
rect -28577 -35512 -28530 -35448
rect -28466 -35512 -28450 -35448
rect -28577 -35528 -28450 -35512
rect -28577 -35592 -28530 -35528
rect -28466 -35592 -28450 -35528
rect -28577 -35608 -28450 -35592
rect -28577 -35672 -28530 -35608
rect -28466 -35672 -28450 -35608
rect -28577 -35688 -28450 -35672
rect -28577 -35752 -28530 -35688
rect -28466 -35752 -28450 -35688
rect -28577 -35768 -28450 -35752
rect -28577 -35832 -28530 -35768
rect -28466 -35832 -28450 -35768
rect -28577 -35848 -28450 -35832
rect -28577 -35912 -28530 -35848
rect -28466 -35912 -28450 -35848
rect -28577 -35928 -28450 -35912
rect -28577 -35992 -28530 -35928
rect -28466 -35992 -28450 -35928
rect -28577 -36008 -28450 -35992
rect -28577 -36072 -28530 -36008
rect -28466 -36072 -28450 -36008
rect -28577 -36088 -28450 -36072
rect -28577 -36152 -28530 -36088
rect -28466 -36152 -28450 -36088
rect -28577 -36168 -28450 -36152
rect -28577 -36232 -28530 -36168
rect -28466 -36232 -28450 -36168
rect -28577 -36248 -28450 -36232
rect -28577 -36312 -28530 -36248
rect -28466 -36312 -28450 -36248
rect -28577 -36328 -28450 -36312
rect -28577 -36392 -28530 -36328
rect -28466 -36392 -28450 -36328
rect -28577 -36408 -28450 -36392
rect -28577 -36472 -28530 -36408
rect -28466 -36472 -28450 -36408
rect -28577 -36488 -28450 -36472
rect -28577 -36552 -28530 -36488
rect -28466 -36552 -28450 -36488
rect -28577 -36568 -28450 -36552
rect -28577 -36632 -28530 -36568
rect -28466 -36632 -28450 -36568
rect -28577 -36648 -28450 -36632
rect -28577 -36712 -28530 -36648
rect -28466 -36712 -28450 -36648
rect -28577 -36728 -28450 -36712
rect -28577 -36792 -28530 -36728
rect -28466 -36792 -28450 -36728
rect -28577 -36808 -28450 -36792
rect -28577 -36872 -28530 -36808
rect -28466 -36872 -28450 -36808
rect -28577 -36888 -28450 -36872
rect -28577 -36952 -28530 -36888
rect -28466 -36952 -28450 -36888
rect -28577 -36968 -28450 -36952
rect -28577 -37032 -28530 -36968
rect -28466 -37032 -28450 -36968
rect -28577 -37048 -28450 -37032
rect -28577 -37112 -28530 -37048
rect -28466 -37112 -28450 -37048
rect -28577 -37128 -28450 -37112
rect -28577 -37192 -28530 -37128
rect -28466 -37192 -28450 -37128
rect -28577 -37208 -28450 -37192
rect -28577 -37272 -28530 -37208
rect -28466 -37272 -28450 -37208
rect -28577 -37288 -28450 -37272
rect -28577 -37352 -28530 -37288
rect -28466 -37352 -28450 -37288
rect -28577 -37368 -28450 -37352
rect -28577 -37432 -28530 -37368
rect -28466 -37432 -28450 -37368
rect -28577 -37448 -28450 -37432
rect -28577 -37512 -28530 -37448
rect -28466 -37512 -28450 -37448
rect -28577 -37528 -28450 -37512
rect -28577 -37592 -28530 -37528
rect -28466 -37592 -28450 -37528
rect -28577 -37608 -28450 -37592
rect -28577 -37672 -28530 -37608
rect -28466 -37672 -28450 -37608
rect -28577 -37688 -28450 -37672
rect -28577 -37752 -28530 -37688
rect -28466 -37752 -28450 -37688
rect -28577 -37768 -28450 -37752
rect -28577 -37832 -28530 -37768
rect -28466 -37832 -28450 -37768
rect -28577 -37848 -28450 -37832
rect -28577 -37912 -28530 -37848
rect -28466 -37912 -28450 -37848
rect -28577 -37928 -28450 -37912
rect -28577 -37992 -28530 -37928
rect -28466 -37992 -28450 -37928
rect -28577 -38008 -28450 -37992
rect -28577 -38072 -28530 -38008
rect -28466 -38072 -28450 -38008
rect -28577 -38088 -28450 -38072
rect -28577 -38152 -28530 -38088
rect -28466 -38152 -28450 -38088
rect -28577 -38168 -28450 -38152
rect -28577 -38232 -28530 -38168
rect -28466 -38232 -28450 -38168
rect -28577 -38248 -28450 -38232
rect -28577 -38312 -28530 -38248
rect -28466 -38312 -28450 -38248
rect -28577 -38328 -28450 -38312
rect -28577 -38392 -28530 -38328
rect -28466 -38392 -28450 -38328
rect -28577 -38408 -28450 -38392
rect -28577 -38472 -28530 -38408
rect -28466 -38472 -28450 -38408
rect -28577 -38488 -28450 -38472
rect -28577 -38552 -28530 -38488
rect -28466 -38552 -28450 -38488
rect -28577 -38568 -28450 -38552
rect -28577 -38632 -28530 -38568
rect -28466 -38632 -28450 -38568
rect -28577 -38648 -28450 -38632
rect -28577 -38712 -28530 -38648
rect -28466 -38712 -28450 -38648
rect -28577 -38728 -28450 -38712
rect -28577 -38792 -28530 -38728
rect -28466 -38792 -28450 -38728
rect -28577 -38808 -28450 -38792
rect -28577 -38872 -28530 -38808
rect -28466 -38872 -28450 -38808
rect -28577 -38888 -28450 -38872
rect -28577 -38952 -28530 -38888
rect -28466 -38952 -28450 -38888
rect -28577 -38968 -28450 -38952
rect -28577 -39032 -28530 -38968
rect -28466 -39032 -28450 -38968
rect -28577 -39048 -28450 -39032
rect -28577 -39112 -28530 -39048
rect -28466 -39112 -28450 -39048
rect -28577 -39128 -28450 -39112
rect -28577 -39192 -28530 -39128
rect -28466 -39192 -28450 -39128
rect -28577 -39208 -28450 -39192
rect -28577 -39272 -28530 -39208
rect -28466 -39272 -28450 -39208
rect -28577 -39288 -28450 -39272
rect -28577 -39352 -28530 -39288
rect -28466 -39352 -28450 -39288
rect -28577 -39368 -28450 -39352
rect -28577 -39432 -28530 -39368
rect -28466 -39432 -28450 -39368
rect -28577 -39448 -28450 -39432
rect -28577 -39512 -28530 -39448
rect -28466 -39512 -28450 -39448
rect -28577 -39528 -28450 -39512
rect -28577 -39592 -28530 -39528
rect -28466 -39592 -28450 -39528
rect -28577 -39608 -28450 -39592
rect -28577 -39672 -28530 -39608
rect -28466 -39672 -28450 -39608
rect -28577 -39688 -28450 -39672
rect -28577 -39752 -28530 -39688
rect -28466 -39752 -28450 -39688
rect -28577 -39768 -28450 -39752
rect -28577 -39832 -28530 -39768
rect -28466 -39832 -28450 -39768
rect -28577 -39848 -28450 -39832
rect -28577 -39912 -28530 -39848
rect -28466 -39912 -28450 -39848
rect -28577 -39928 -28450 -39912
rect -28577 -39992 -28530 -39928
rect -28466 -39992 -28450 -39928
rect -28577 -40008 -28450 -39992
rect -28577 -40072 -28530 -40008
rect -28466 -40072 -28450 -40008
rect -28577 -40088 -28450 -40072
rect -28577 -40152 -28530 -40088
rect -28466 -40152 -28450 -40088
rect -28577 -40168 -28450 -40152
rect -28577 -40232 -28530 -40168
rect -28466 -40232 -28450 -40168
rect -28577 -40248 -28450 -40232
rect -28577 -40312 -28530 -40248
rect -28466 -40312 -28450 -40248
rect -28577 -40328 -28450 -40312
rect -28577 -40392 -28530 -40328
rect -28466 -40392 -28450 -40328
rect -28577 -40408 -28450 -40392
rect -28577 -40472 -28530 -40408
rect -28466 -40472 -28450 -40408
rect -28577 -40488 -28450 -40472
rect -28577 -40552 -28530 -40488
rect -28466 -40552 -28450 -40488
rect -28577 -40568 -28450 -40552
rect -28577 -40632 -28530 -40568
rect -28466 -40632 -28450 -40568
rect -28577 -40648 -28450 -40632
rect -28577 -40712 -28530 -40648
rect -28466 -40712 -28450 -40648
rect -28577 -40728 -28450 -40712
rect -34896 -40808 -34769 -40792
rect -34896 -40872 -34849 -40808
rect -34785 -40872 -34769 -40808
rect -34896 -40888 -34769 -40872
rect -34896 -41012 -34792 -40888
rect -34896 -41028 -34769 -41012
rect -34896 -41092 -34849 -41028
rect -34785 -41092 -34769 -41028
rect -34896 -41108 -34769 -41092
rect -41215 -41188 -41088 -41172
rect -41215 -41252 -41168 -41188
rect -41104 -41252 -41088 -41188
rect -41215 -41268 -41088 -41252
rect -41215 -41332 -41168 -41268
rect -41104 -41332 -41088 -41268
rect -41215 -41348 -41088 -41332
rect -41215 -41412 -41168 -41348
rect -41104 -41412 -41088 -41348
rect -41215 -41428 -41088 -41412
rect -41215 -41492 -41168 -41428
rect -41104 -41492 -41088 -41428
rect -41215 -41508 -41088 -41492
rect -41215 -41572 -41168 -41508
rect -41104 -41572 -41088 -41508
rect -41215 -41588 -41088 -41572
rect -41215 -41652 -41168 -41588
rect -41104 -41652 -41088 -41588
rect -41215 -41668 -41088 -41652
rect -41215 -41732 -41168 -41668
rect -41104 -41732 -41088 -41668
rect -41215 -41748 -41088 -41732
rect -41215 -41812 -41168 -41748
rect -41104 -41812 -41088 -41748
rect -41215 -41828 -41088 -41812
rect -41215 -41892 -41168 -41828
rect -41104 -41892 -41088 -41828
rect -41215 -41908 -41088 -41892
rect -41215 -41972 -41168 -41908
rect -41104 -41972 -41088 -41908
rect -41215 -41988 -41088 -41972
rect -41215 -42052 -41168 -41988
rect -41104 -42052 -41088 -41988
rect -41215 -42068 -41088 -42052
rect -41215 -42132 -41168 -42068
rect -41104 -42132 -41088 -42068
rect -41215 -42148 -41088 -42132
rect -41215 -42212 -41168 -42148
rect -41104 -42212 -41088 -42148
rect -41215 -42228 -41088 -42212
rect -41215 -42292 -41168 -42228
rect -41104 -42292 -41088 -42228
rect -41215 -42308 -41088 -42292
rect -41215 -42372 -41168 -42308
rect -41104 -42372 -41088 -42308
rect -41215 -42388 -41088 -42372
rect -41215 -42452 -41168 -42388
rect -41104 -42452 -41088 -42388
rect -41215 -42468 -41088 -42452
rect -41215 -42532 -41168 -42468
rect -41104 -42532 -41088 -42468
rect -41215 -42548 -41088 -42532
rect -41215 -42612 -41168 -42548
rect -41104 -42612 -41088 -42548
rect -41215 -42628 -41088 -42612
rect -41215 -42692 -41168 -42628
rect -41104 -42692 -41088 -42628
rect -41215 -42708 -41088 -42692
rect -41215 -42772 -41168 -42708
rect -41104 -42772 -41088 -42708
rect -41215 -42788 -41088 -42772
rect -41215 -42852 -41168 -42788
rect -41104 -42852 -41088 -42788
rect -41215 -42868 -41088 -42852
rect -41215 -42932 -41168 -42868
rect -41104 -42932 -41088 -42868
rect -41215 -42948 -41088 -42932
rect -41215 -43012 -41168 -42948
rect -41104 -43012 -41088 -42948
rect -41215 -43028 -41088 -43012
rect -41215 -43092 -41168 -43028
rect -41104 -43092 -41088 -43028
rect -41215 -43108 -41088 -43092
rect -41215 -43172 -41168 -43108
rect -41104 -43172 -41088 -43108
rect -41215 -43188 -41088 -43172
rect -41215 -43252 -41168 -43188
rect -41104 -43252 -41088 -43188
rect -41215 -43268 -41088 -43252
rect -41215 -43332 -41168 -43268
rect -41104 -43332 -41088 -43268
rect -41215 -43348 -41088 -43332
rect -41215 -43412 -41168 -43348
rect -41104 -43412 -41088 -43348
rect -41215 -43428 -41088 -43412
rect -41215 -43492 -41168 -43428
rect -41104 -43492 -41088 -43428
rect -41215 -43508 -41088 -43492
rect -41215 -43572 -41168 -43508
rect -41104 -43572 -41088 -43508
rect -41215 -43588 -41088 -43572
rect -41215 -43652 -41168 -43588
rect -41104 -43652 -41088 -43588
rect -41215 -43668 -41088 -43652
rect -41215 -43732 -41168 -43668
rect -41104 -43732 -41088 -43668
rect -41215 -43748 -41088 -43732
rect -41215 -43812 -41168 -43748
rect -41104 -43812 -41088 -43748
rect -41215 -43828 -41088 -43812
rect -41215 -43892 -41168 -43828
rect -41104 -43892 -41088 -43828
rect -41215 -43908 -41088 -43892
rect -41215 -43972 -41168 -43908
rect -41104 -43972 -41088 -43908
rect -41215 -43988 -41088 -43972
rect -41215 -44052 -41168 -43988
rect -41104 -44052 -41088 -43988
rect -41215 -44068 -41088 -44052
rect -41215 -44132 -41168 -44068
rect -41104 -44132 -41088 -44068
rect -41215 -44148 -41088 -44132
rect -41215 -44212 -41168 -44148
rect -41104 -44212 -41088 -44148
rect -41215 -44228 -41088 -44212
rect -41215 -44292 -41168 -44228
rect -41104 -44292 -41088 -44228
rect -41215 -44308 -41088 -44292
rect -41215 -44372 -41168 -44308
rect -41104 -44372 -41088 -44308
rect -41215 -44388 -41088 -44372
rect -41215 -44452 -41168 -44388
rect -41104 -44452 -41088 -44388
rect -41215 -44468 -41088 -44452
rect -41215 -44532 -41168 -44468
rect -41104 -44532 -41088 -44468
rect -41215 -44548 -41088 -44532
rect -41215 -44612 -41168 -44548
rect -41104 -44612 -41088 -44548
rect -41215 -44628 -41088 -44612
rect -41215 -44692 -41168 -44628
rect -41104 -44692 -41088 -44628
rect -41215 -44708 -41088 -44692
rect -41215 -44772 -41168 -44708
rect -41104 -44772 -41088 -44708
rect -41215 -44788 -41088 -44772
rect -41215 -44852 -41168 -44788
rect -41104 -44852 -41088 -44788
rect -41215 -44868 -41088 -44852
rect -41215 -44932 -41168 -44868
rect -41104 -44932 -41088 -44868
rect -41215 -44948 -41088 -44932
rect -41215 -45012 -41168 -44948
rect -41104 -45012 -41088 -44948
rect -41215 -45028 -41088 -45012
rect -41215 -45092 -41168 -45028
rect -41104 -45092 -41088 -45028
rect -41215 -45108 -41088 -45092
rect -41215 -45172 -41168 -45108
rect -41104 -45172 -41088 -45108
rect -41215 -45188 -41088 -45172
rect -41215 -45252 -41168 -45188
rect -41104 -45252 -41088 -45188
rect -41215 -45268 -41088 -45252
rect -41215 -45332 -41168 -45268
rect -41104 -45332 -41088 -45268
rect -41215 -45348 -41088 -45332
rect -41215 -45412 -41168 -45348
rect -41104 -45412 -41088 -45348
rect -41215 -45428 -41088 -45412
rect -41215 -45492 -41168 -45428
rect -41104 -45492 -41088 -45428
rect -41215 -45508 -41088 -45492
rect -41215 -45572 -41168 -45508
rect -41104 -45572 -41088 -45508
rect -41215 -45588 -41088 -45572
rect -41215 -45652 -41168 -45588
rect -41104 -45652 -41088 -45588
rect -41215 -45668 -41088 -45652
rect -41215 -45732 -41168 -45668
rect -41104 -45732 -41088 -45668
rect -41215 -45748 -41088 -45732
rect -41215 -45812 -41168 -45748
rect -41104 -45812 -41088 -45748
rect -41215 -45828 -41088 -45812
rect -41215 -45892 -41168 -45828
rect -41104 -45892 -41088 -45828
rect -41215 -45908 -41088 -45892
rect -41215 -45972 -41168 -45908
rect -41104 -45972 -41088 -45908
rect -41215 -45988 -41088 -45972
rect -41215 -46052 -41168 -45988
rect -41104 -46052 -41088 -45988
rect -41215 -46068 -41088 -46052
rect -41215 -46132 -41168 -46068
rect -41104 -46132 -41088 -46068
rect -41215 -46148 -41088 -46132
rect -41215 -46212 -41168 -46148
rect -41104 -46212 -41088 -46148
rect -41215 -46228 -41088 -46212
rect -41215 -46292 -41168 -46228
rect -41104 -46292 -41088 -46228
rect -41215 -46308 -41088 -46292
rect -41215 -46372 -41168 -46308
rect -41104 -46372 -41088 -46308
rect -41215 -46388 -41088 -46372
rect -41215 -46452 -41168 -46388
rect -41104 -46452 -41088 -46388
rect -41215 -46468 -41088 -46452
rect -41215 -46532 -41168 -46468
rect -41104 -46532 -41088 -46468
rect -41215 -46548 -41088 -46532
rect -41215 -46612 -41168 -46548
rect -41104 -46612 -41088 -46548
rect -41215 -46628 -41088 -46612
rect -41215 -46692 -41168 -46628
rect -41104 -46692 -41088 -46628
rect -41215 -46708 -41088 -46692
rect -41215 -46772 -41168 -46708
rect -41104 -46772 -41088 -46708
rect -41215 -46788 -41088 -46772
rect -41215 -46852 -41168 -46788
rect -41104 -46852 -41088 -46788
rect -41215 -46868 -41088 -46852
rect -41215 -46932 -41168 -46868
rect -41104 -46932 -41088 -46868
rect -41215 -46948 -41088 -46932
rect -41215 -47012 -41168 -46948
rect -41104 -47012 -41088 -46948
rect -41215 -47028 -41088 -47012
rect -44335 -47250 -44231 -47061
rect -41215 -47092 -41168 -47028
rect -41104 -47092 -41088 -47028
rect -40925 -41148 -35003 -41139
rect -40925 -47052 -40916 -41148
rect -35012 -47052 -35003 -41148
rect -40925 -47061 -35003 -47052
rect -34896 -41172 -34849 -41108
rect -34785 -41172 -34769 -41108
rect -31697 -41139 -31593 -40761
rect -28577 -40792 -28530 -40728
rect -28466 -40792 -28450 -40728
rect -28287 -34848 -22365 -34839
rect -28287 -40752 -28278 -34848
rect -22374 -40752 -22365 -34848
rect -28287 -40761 -22365 -40752
rect -22258 -34872 -22211 -34808
rect -22147 -34872 -22131 -34808
rect -19059 -34839 -18955 -34461
rect -15939 -34492 -15892 -34428
rect -15828 -34492 -15812 -34428
rect -15649 -28548 -9727 -28539
rect -15649 -34452 -15640 -28548
rect -9736 -34452 -9727 -28548
rect -15649 -34461 -9727 -34452
rect -9620 -28572 -9573 -28508
rect -9509 -28572 -9493 -28508
rect -6421 -28539 -6317 -28161
rect -3301 -28192 -3254 -28128
rect -3190 -28192 -3174 -28128
rect -3011 -22248 2911 -22239
rect -3011 -28152 -3002 -22248
rect 2902 -28152 2911 -22248
rect -3011 -28161 2911 -28152
rect 3018 -22272 3065 -22208
rect 3129 -22272 3145 -22208
rect 6217 -22239 6321 -21861
rect 9337 -21892 9384 -21828
rect 9448 -21892 9464 -21828
rect 9627 -15948 15549 -15939
rect 9627 -21852 9636 -15948
rect 15540 -21852 15549 -15948
rect 9627 -21861 15549 -21852
rect 15656 -15972 15703 -15908
rect 15767 -15972 15783 -15908
rect 18855 -15939 18959 -15561
rect 21975 -15592 22022 -15528
rect 22086 -15592 22102 -15528
rect 22265 -9648 28187 -9639
rect 22265 -15552 22274 -9648
rect 28178 -15552 28187 -9648
rect 22265 -15561 28187 -15552
rect 28294 -9672 28341 -9608
rect 28405 -9672 28421 -9608
rect 31493 -9639 31597 -9261
rect 34613 -9292 34660 -9228
rect 34724 -9292 34740 -9228
rect 34903 -3348 40825 -3339
rect 34903 -9252 34912 -3348
rect 40816 -9252 40825 -3348
rect 34903 -9261 40825 -9252
rect 40932 -3372 40979 -3308
rect 41043 -3372 41059 -3308
rect 44131 -3339 44235 -2961
rect 47251 -2992 47298 -2928
rect 47362 -2992 47378 -2928
rect 47251 -3008 47378 -2992
rect 47251 -3072 47298 -3008
rect 47362 -3072 47378 -3008
rect 47251 -3088 47378 -3072
rect 47251 -3212 47355 -3088
rect 47251 -3228 47378 -3212
rect 47251 -3292 47298 -3228
rect 47362 -3292 47378 -3228
rect 47251 -3308 47378 -3292
rect 40932 -3388 41059 -3372
rect 40932 -3452 40979 -3388
rect 41043 -3452 41059 -3388
rect 40932 -3468 41059 -3452
rect 40932 -3532 40979 -3468
rect 41043 -3532 41059 -3468
rect 40932 -3548 41059 -3532
rect 40932 -3612 40979 -3548
rect 41043 -3612 41059 -3548
rect 40932 -3628 41059 -3612
rect 40932 -3692 40979 -3628
rect 41043 -3692 41059 -3628
rect 40932 -3708 41059 -3692
rect 40932 -3772 40979 -3708
rect 41043 -3772 41059 -3708
rect 40932 -3788 41059 -3772
rect 40932 -3852 40979 -3788
rect 41043 -3852 41059 -3788
rect 40932 -3868 41059 -3852
rect 40932 -3932 40979 -3868
rect 41043 -3932 41059 -3868
rect 40932 -3948 41059 -3932
rect 40932 -4012 40979 -3948
rect 41043 -4012 41059 -3948
rect 40932 -4028 41059 -4012
rect 40932 -4092 40979 -4028
rect 41043 -4092 41059 -4028
rect 40932 -4108 41059 -4092
rect 40932 -4172 40979 -4108
rect 41043 -4172 41059 -4108
rect 40932 -4188 41059 -4172
rect 40932 -4252 40979 -4188
rect 41043 -4252 41059 -4188
rect 40932 -4268 41059 -4252
rect 40932 -4332 40979 -4268
rect 41043 -4332 41059 -4268
rect 40932 -4348 41059 -4332
rect 40932 -4412 40979 -4348
rect 41043 -4412 41059 -4348
rect 40932 -4428 41059 -4412
rect 40932 -4492 40979 -4428
rect 41043 -4492 41059 -4428
rect 40932 -4508 41059 -4492
rect 40932 -4572 40979 -4508
rect 41043 -4572 41059 -4508
rect 40932 -4588 41059 -4572
rect 40932 -4652 40979 -4588
rect 41043 -4652 41059 -4588
rect 40932 -4668 41059 -4652
rect 40932 -4732 40979 -4668
rect 41043 -4732 41059 -4668
rect 40932 -4748 41059 -4732
rect 40932 -4812 40979 -4748
rect 41043 -4812 41059 -4748
rect 40932 -4828 41059 -4812
rect 40932 -4892 40979 -4828
rect 41043 -4892 41059 -4828
rect 40932 -4908 41059 -4892
rect 40932 -4972 40979 -4908
rect 41043 -4972 41059 -4908
rect 40932 -4988 41059 -4972
rect 40932 -5052 40979 -4988
rect 41043 -5052 41059 -4988
rect 40932 -5068 41059 -5052
rect 40932 -5132 40979 -5068
rect 41043 -5132 41059 -5068
rect 40932 -5148 41059 -5132
rect 40932 -5212 40979 -5148
rect 41043 -5212 41059 -5148
rect 40932 -5228 41059 -5212
rect 40932 -5292 40979 -5228
rect 41043 -5292 41059 -5228
rect 40932 -5308 41059 -5292
rect 40932 -5372 40979 -5308
rect 41043 -5372 41059 -5308
rect 40932 -5388 41059 -5372
rect 40932 -5452 40979 -5388
rect 41043 -5452 41059 -5388
rect 40932 -5468 41059 -5452
rect 40932 -5532 40979 -5468
rect 41043 -5532 41059 -5468
rect 40932 -5548 41059 -5532
rect 40932 -5612 40979 -5548
rect 41043 -5612 41059 -5548
rect 40932 -5628 41059 -5612
rect 40932 -5692 40979 -5628
rect 41043 -5692 41059 -5628
rect 40932 -5708 41059 -5692
rect 40932 -5772 40979 -5708
rect 41043 -5772 41059 -5708
rect 40932 -5788 41059 -5772
rect 40932 -5852 40979 -5788
rect 41043 -5852 41059 -5788
rect 40932 -5868 41059 -5852
rect 40932 -5932 40979 -5868
rect 41043 -5932 41059 -5868
rect 40932 -5948 41059 -5932
rect 40932 -6012 40979 -5948
rect 41043 -6012 41059 -5948
rect 40932 -6028 41059 -6012
rect 40932 -6092 40979 -6028
rect 41043 -6092 41059 -6028
rect 40932 -6108 41059 -6092
rect 40932 -6172 40979 -6108
rect 41043 -6172 41059 -6108
rect 40932 -6188 41059 -6172
rect 40932 -6252 40979 -6188
rect 41043 -6252 41059 -6188
rect 40932 -6268 41059 -6252
rect 40932 -6332 40979 -6268
rect 41043 -6332 41059 -6268
rect 40932 -6348 41059 -6332
rect 40932 -6412 40979 -6348
rect 41043 -6412 41059 -6348
rect 40932 -6428 41059 -6412
rect 40932 -6492 40979 -6428
rect 41043 -6492 41059 -6428
rect 40932 -6508 41059 -6492
rect 40932 -6572 40979 -6508
rect 41043 -6572 41059 -6508
rect 40932 -6588 41059 -6572
rect 40932 -6652 40979 -6588
rect 41043 -6652 41059 -6588
rect 40932 -6668 41059 -6652
rect 40932 -6732 40979 -6668
rect 41043 -6732 41059 -6668
rect 40932 -6748 41059 -6732
rect 40932 -6812 40979 -6748
rect 41043 -6812 41059 -6748
rect 40932 -6828 41059 -6812
rect 40932 -6892 40979 -6828
rect 41043 -6892 41059 -6828
rect 40932 -6908 41059 -6892
rect 40932 -6972 40979 -6908
rect 41043 -6972 41059 -6908
rect 40932 -6988 41059 -6972
rect 40932 -7052 40979 -6988
rect 41043 -7052 41059 -6988
rect 40932 -7068 41059 -7052
rect 40932 -7132 40979 -7068
rect 41043 -7132 41059 -7068
rect 40932 -7148 41059 -7132
rect 40932 -7212 40979 -7148
rect 41043 -7212 41059 -7148
rect 40932 -7228 41059 -7212
rect 40932 -7292 40979 -7228
rect 41043 -7292 41059 -7228
rect 40932 -7308 41059 -7292
rect 40932 -7372 40979 -7308
rect 41043 -7372 41059 -7308
rect 40932 -7388 41059 -7372
rect 40932 -7452 40979 -7388
rect 41043 -7452 41059 -7388
rect 40932 -7468 41059 -7452
rect 40932 -7532 40979 -7468
rect 41043 -7532 41059 -7468
rect 40932 -7548 41059 -7532
rect 40932 -7612 40979 -7548
rect 41043 -7612 41059 -7548
rect 40932 -7628 41059 -7612
rect 40932 -7692 40979 -7628
rect 41043 -7692 41059 -7628
rect 40932 -7708 41059 -7692
rect 40932 -7772 40979 -7708
rect 41043 -7772 41059 -7708
rect 40932 -7788 41059 -7772
rect 40932 -7852 40979 -7788
rect 41043 -7852 41059 -7788
rect 40932 -7868 41059 -7852
rect 40932 -7932 40979 -7868
rect 41043 -7932 41059 -7868
rect 40932 -7948 41059 -7932
rect 40932 -8012 40979 -7948
rect 41043 -8012 41059 -7948
rect 40932 -8028 41059 -8012
rect 40932 -8092 40979 -8028
rect 41043 -8092 41059 -8028
rect 40932 -8108 41059 -8092
rect 40932 -8172 40979 -8108
rect 41043 -8172 41059 -8108
rect 40932 -8188 41059 -8172
rect 40932 -8252 40979 -8188
rect 41043 -8252 41059 -8188
rect 40932 -8268 41059 -8252
rect 40932 -8332 40979 -8268
rect 41043 -8332 41059 -8268
rect 40932 -8348 41059 -8332
rect 40932 -8412 40979 -8348
rect 41043 -8412 41059 -8348
rect 40932 -8428 41059 -8412
rect 40932 -8492 40979 -8428
rect 41043 -8492 41059 -8428
rect 40932 -8508 41059 -8492
rect 40932 -8572 40979 -8508
rect 41043 -8572 41059 -8508
rect 40932 -8588 41059 -8572
rect 40932 -8652 40979 -8588
rect 41043 -8652 41059 -8588
rect 40932 -8668 41059 -8652
rect 40932 -8732 40979 -8668
rect 41043 -8732 41059 -8668
rect 40932 -8748 41059 -8732
rect 40932 -8812 40979 -8748
rect 41043 -8812 41059 -8748
rect 40932 -8828 41059 -8812
rect 40932 -8892 40979 -8828
rect 41043 -8892 41059 -8828
rect 40932 -8908 41059 -8892
rect 40932 -8972 40979 -8908
rect 41043 -8972 41059 -8908
rect 40932 -8988 41059 -8972
rect 40932 -9052 40979 -8988
rect 41043 -9052 41059 -8988
rect 40932 -9068 41059 -9052
rect 40932 -9132 40979 -9068
rect 41043 -9132 41059 -9068
rect 40932 -9148 41059 -9132
rect 40932 -9212 40979 -9148
rect 41043 -9212 41059 -9148
rect 40932 -9228 41059 -9212
rect 34613 -9308 34740 -9292
rect 34613 -9372 34660 -9308
rect 34724 -9372 34740 -9308
rect 34613 -9388 34740 -9372
rect 34613 -9512 34717 -9388
rect 34613 -9528 34740 -9512
rect 34613 -9592 34660 -9528
rect 34724 -9592 34740 -9528
rect 34613 -9608 34740 -9592
rect 28294 -9688 28421 -9672
rect 28294 -9752 28341 -9688
rect 28405 -9752 28421 -9688
rect 28294 -9768 28421 -9752
rect 28294 -9832 28341 -9768
rect 28405 -9832 28421 -9768
rect 28294 -9848 28421 -9832
rect 28294 -9912 28341 -9848
rect 28405 -9912 28421 -9848
rect 28294 -9928 28421 -9912
rect 28294 -9992 28341 -9928
rect 28405 -9992 28421 -9928
rect 28294 -10008 28421 -9992
rect 28294 -10072 28341 -10008
rect 28405 -10072 28421 -10008
rect 28294 -10088 28421 -10072
rect 28294 -10152 28341 -10088
rect 28405 -10152 28421 -10088
rect 28294 -10168 28421 -10152
rect 28294 -10232 28341 -10168
rect 28405 -10232 28421 -10168
rect 28294 -10248 28421 -10232
rect 28294 -10312 28341 -10248
rect 28405 -10312 28421 -10248
rect 28294 -10328 28421 -10312
rect 28294 -10392 28341 -10328
rect 28405 -10392 28421 -10328
rect 28294 -10408 28421 -10392
rect 28294 -10472 28341 -10408
rect 28405 -10472 28421 -10408
rect 28294 -10488 28421 -10472
rect 28294 -10552 28341 -10488
rect 28405 -10552 28421 -10488
rect 28294 -10568 28421 -10552
rect 28294 -10632 28341 -10568
rect 28405 -10632 28421 -10568
rect 28294 -10648 28421 -10632
rect 28294 -10712 28341 -10648
rect 28405 -10712 28421 -10648
rect 28294 -10728 28421 -10712
rect 28294 -10792 28341 -10728
rect 28405 -10792 28421 -10728
rect 28294 -10808 28421 -10792
rect 28294 -10872 28341 -10808
rect 28405 -10872 28421 -10808
rect 28294 -10888 28421 -10872
rect 28294 -10952 28341 -10888
rect 28405 -10952 28421 -10888
rect 28294 -10968 28421 -10952
rect 28294 -11032 28341 -10968
rect 28405 -11032 28421 -10968
rect 28294 -11048 28421 -11032
rect 28294 -11112 28341 -11048
rect 28405 -11112 28421 -11048
rect 28294 -11128 28421 -11112
rect 28294 -11192 28341 -11128
rect 28405 -11192 28421 -11128
rect 28294 -11208 28421 -11192
rect 28294 -11272 28341 -11208
rect 28405 -11272 28421 -11208
rect 28294 -11288 28421 -11272
rect 28294 -11352 28341 -11288
rect 28405 -11352 28421 -11288
rect 28294 -11368 28421 -11352
rect 28294 -11432 28341 -11368
rect 28405 -11432 28421 -11368
rect 28294 -11448 28421 -11432
rect 28294 -11512 28341 -11448
rect 28405 -11512 28421 -11448
rect 28294 -11528 28421 -11512
rect 28294 -11592 28341 -11528
rect 28405 -11592 28421 -11528
rect 28294 -11608 28421 -11592
rect 28294 -11672 28341 -11608
rect 28405 -11672 28421 -11608
rect 28294 -11688 28421 -11672
rect 28294 -11752 28341 -11688
rect 28405 -11752 28421 -11688
rect 28294 -11768 28421 -11752
rect 28294 -11832 28341 -11768
rect 28405 -11832 28421 -11768
rect 28294 -11848 28421 -11832
rect 28294 -11912 28341 -11848
rect 28405 -11912 28421 -11848
rect 28294 -11928 28421 -11912
rect 28294 -11992 28341 -11928
rect 28405 -11992 28421 -11928
rect 28294 -12008 28421 -11992
rect 28294 -12072 28341 -12008
rect 28405 -12072 28421 -12008
rect 28294 -12088 28421 -12072
rect 28294 -12152 28341 -12088
rect 28405 -12152 28421 -12088
rect 28294 -12168 28421 -12152
rect 28294 -12232 28341 -12168
rect 28405 -12232 28421 -12168
rect 28294 -12248 28421 -12232
rect 28294 -12312 28341 -12248
rect 28405 -12312 28421 -12248
rect 28294 -12328 28421 -12312
rect 28294 -12392 28341 -12328
rect 28405 -12392 28421 -12328
rect 28294 -12408 28421 -12392
rect 28294 -12472 28341 -12408
rect 28405 -12472 28421 -12408
rect 28294 -12488 28421 -12472
rect 28294 -12552 28341 -12488
rect 28405 -12552 28421 -12488
rect 28294 -12568 28421 -12552
rect 28294 -12632 28341 -12568
rect 28405 -12632 28421 -12568
rect 28294 -12648 28421 -12632
rect 28294 -12712 28341 -12648
rect 28405 -12712 28421 -12648
rect 28294 -12728 28421 -12712
rect 28294 -12792 28341 -12728
rect 28405 -12792 28421 -12728
rect 28294 -12808 28421 -12792
rect 28294 -12872 28341 -12808
rect 28405 -12872 28421 -12808
rect 28294 -12888 28421 -12872
rect 28294 -12952 28341 -12888
rect 28405 -12952 28421 -12888
rect 28294 -12968 28421 -12952
rect 28294 -13032 28341 -12968
rect 28405 -13032 28421 -12968
rect 28294 -13048 28421 -13032
rect 28294 -13112 28341 -13048
rect 28405 -13112 28421 -13048
rect 28294 -13128 28421 -13112
rect 28294 -13192 28341 -13128
rect 28405 -13192 28421 -13128
rect 28294 -13208 28421 -13192
rect 28294 -13272 28341 -13208
rect 28405 -13272 28421 -13208
rect 28294 -13288 28421 -13272
rect 28294 -13352 28341 -13288
rect 28405 -13352 28421 -13288
rect 28294 -13368 28421 -13352
rect 28294 -13432 28341 -13368
rect 28405 -13432 28421 -13368
rect 28294 -13448 28421 -13432
rect 28294 -13512 28341 -13448
rect 28405 -13512 28421 -13448
rect 28294 -13528 28421 -13512
rect 28294 -13592 28341 -13528
rect 28405 -13592 28421 -13528
rect 28294 -13608 28421 -13592
rect 28294 -13672 28341 -13608
rect 28405 -13672 28421 -13608
rect 28294 -13688 28421 -13672
rect 28294 -13752 28341 -13688
rect 28405 -13752 28421 -13688
rect 28294 -13768 28421 -13752
rect 28294 -13832 28341 -13768
rect 28405 -13832 28421 -13768
rect 28294 -13848 28421 -13832
rect 28294 -13912 28341 -13848
rect 28405 -13912 28421 -13848
rect 28294 -13928 28421 -13912
rect 28294 -13992 28341 -13928
rect 28405 -13992 28421 -13928
rect 28294 -14008 28421 -13992
rect 28294 -14072 28341 -14008
rect 28405 -14072 28421 -14008
rect 28294 -14088 28421 -14072
rect 28294 -14152 28341 -14088
rect 28405 -14152 28421 -14088
rect 28294 -14168 28421 -14152
rect 28294 -14232 28341 -14168
rect 28405 -14232 28421 -14168
rect 28294 -14248 28421 -14232
rect 28294 -14312 28341 -14248
rect 28405 -14312 28421 -14248
rect 28294 -14328 28421 -14312
rect 28294 -14392 28341 -14328
rect 28405 -14392 28421 -14328
rect 28294 -14408 28421 -14392
rect 28294 -14472 28341 -14408
rect 28405 -14472 28421 -14408
rect 28294 -14488 28421 -14472
rect 28294 -14552 28341 -14488
rect 28405 -14552 28421 -14488
rect 28294 -14568 28421 -14552
rect 28294 -14632 28341 -14568
rect 28405 -14632 28421 -14568
rect 28294 -14648 28421 -14632
rect 28294 -14712 28341 -14648
rect 28405 -14712 28421 -14648
rect 28294 -14728 28421 -14712
rect 28294 -14792 28341 -14728
rect 28405 -14792 28421 -14728
rect 28294 -14808 28421 -14792
rect 28294 -14872 28341 -14808
rect 28405 -14872 28421 -14808
rect 28294 -14888 28421 -14872
rect 28294 -14952 28341 -14888
rect 28405 -14952 28421 -14888
rect 28294 -14968 28421 -14952
rect 28294 -15032 28341 -14968
rect 28405 -15032 28421 -14968
rect 28294 -15048 28421 -15032
rect 28294 -15112 28341 -15048
rect 28405 -15112 28421 -15048
rect 28294 -15128 28421 -15112
rect 28294 -15192 28341 -15128
rect 28405 -15192 28421 -15128
rect 28294 -15208 28421 -15192
rect 28294 -15272 28341 -15208
rect 28405 -15272 28421 -15208
rect 28294 -15288 28421 -15272
rect 28294 -15352 28341 -15288
rect 28405 -15352 28421 -15288
rect 28294 -15368 28421 -15352
rect 28294 -15432 28341 -15368
rect 28405 -15432 28421 -15368
rect 28294 -15448 28421 -15432
rect 28294 -15512 28341 -15448
rect 28405 -15512 28421 -15448
rect 28294 -15528 28421 -15512
rect 21975 -15608 22102 -15592
rect 21975 -15672 22022 -15608
rect 22086 -15672 22102 -15608
rect 21975 -15688 22102 -15672
rect 21975 -15812 22079 -15688
rect 21975 -15828 22102 -15812
rect 21975 -15892 22022 -15828
rect 22086 -15892 22102 -15828
rect 21975 -15908 22102 -15892
rect 15656 -15988 15783 -15972
rect 15656 -16052 15703 -15988
rect 15767 -16052 15783 -15988
rect 15656 -16068 15783 -16052
rect 15656 -16132 15703 -16068
rect 15767 -16132 15783 -16068
rect 15656 -16148 15783 -16132
rect 15656 -16212 15703 -16148
rect 15767 -16212 15783 -16148
rect 15656 -16228 15783 -16212
rect 15656 -16292 15703 -16228
rect 15767 -16292 15783 -16228
rect 15656 -16308 15783 -16292
rect 15656 -16372 15703 -16308
rect 15767 -16372 15783 -16308
rect 15656 -16388 15783 -16372
rect 15656 -16452 15703 -16388
rect 15767 -16452 15783 -16388
rect 15656 -16468 15783 -16452
rect 15656 -16532 15703 -16468
rect 15767 -16532 15783 -16468
rect 15656 -16548 15783 -16532
rect 15656 -16612 15703 -16548
rect 15767 -16612 15783 -16548
rect 15656 -16628 15783 -16612
rect 15656 -16692 15703 -16628
rect 15767 -16692 15783 -16628
rect 15656 -16708 15783 -16692
rect 15656 -16772 15703 -16708
rect 15767 -16772 15783 -16708
rect 15656 -16788 15783 -16772
rect 15656 -16852 15703 -16788
rect 15767 -16852 15783 -16788
rect 15656 -16868 15783 -16852
rect 15656 -16932 15703 -16868
rect 15767 -16932 15783 -16868
rect 15656 -16948 15783 -16932
rect 15656 -17012 15703 -16948
rect 15767 -17012 15783 -16948
rect 15656 -17028 15783 -17012
rect 15656 -17092 15703 -17028
rect 15767 -17092 15783 -17028
rect 15656 -17108 15783 -17092
rect 15656 -17172 15703 -17108
rect 15767 -17172 15783 -17108
rect 15656 -17188 15783 -17172
rect 15656 -17252 15703 -17188
rect 15767 -17252 15783 -17188
rect 15656 -17268 15783 -17252
rect 15656 -17332 15703 -17268
rect 15767 -17332 15783 -17268
rect 15656 -17348 15783 -17332
rect 15656 -17412 15703 -17348
rect 15767 -17412 15783 -17348
rect 15656 -17428 15783 -17412
rect 15656 -17492 15703 -17428
rect 15767 -17492 15783 -17428
rect 15656 -17508 15783 -17492
rect 15656 -17572 15703 -17508
rect 15767 -17572 15783 -17508
rect 15656 -17588 15783 -17572
rect 15656 -17652 15703 -17588
rect 15767 -17652 15783 -17588
rect 15656 -17668 15783 -17652
rect 15656 -17732 15703 -17668
rect 15767 -17732 15783 -17668
rect 15656 -17748 15783 -17732
rect 15656 -17812 15703 -17748
rect 15767 -17812 15783 -17748
rect 15656 -17828 15783 -17812
rect 15656 -17892 15703 -17828
rect 15767 -17892 15783 -17828
rect 15656 -17908 15783 -17892
rect 15656 -17972 15703 -17908
rect 15767 -17972 15783 -17908
rect 15656 -17988 15783 -17972
rect 15656 -18052 15703 -17988
rect 15767 -18052 15783 -17988
rect 15656 -18068 15783 -18052
rect 15656 -18132 15703 -18068
rect 15767 -18132 15783 -18068
rect 15656 -18148 15783 -18132
rect 15656 -18212 15703 -18148
rect 15767 -18212 15783 -18148
rect 15656 -18228 15783 -18212
rect 15656 -18292 15703 -18228
rect 15767 -18292 15783 -18228
rect 15656 -18308 15783 -18292
rect 15656 -18372 15703 -18308
rect 15767 -18372 15783 -18308
rect 15656 -18388 15783 -18372
rect 15656 -18452 15703 -18388
rect 15767 -18452 15783 -18388
rect 15656 -18468 15783 -18452
rect 15656 -18532 15703 -18468
rect 15767 -18532 15783 -18468
rect 15656 -18548 15783 -18532
rect 15656 -18612 15703 -18548
rect 15767 -18612 15783 -18548
rect 15656 -18628 15783 -18612
rect 15656 -18692 15703 -18628
rect 15767 -18692 15783 -18628
rect 15656 -18708 15783 -18692
rect 15656 -18772 15703 -18708
rect 15767 -18772 15783 -18708
rect 15656 -18788 15783 -18772
rect 15656 -18852 15703 -18788
rect 15767 -18852 15783 -18788
rect 15656 -18868 15783 -18852
rect 15656 -18932 15703 -18868
rect 15767 -18932 15783 -18868
rect 15656 -18948 15783 -18932
rect 15656 -19012 15703 -18948
rect 15767 -19012 15783 -18948
rect 15656 -19028 15783 -19012
rect 15656 -19092 15703 -19028
rect 15767 -19092 15783 -19028
rect 15656 -19108 15783 -19092
rect 15656 -19172 15703 -19108
rect 15767 -19172 15783 -19108
rect 15656 -19188 15783 -19172
rect 15656 -19252 15703 -19188
rect 15767 -19252 15783 -19188
rect 15656 -19268 15783 -19252
rect 15656 -19332 15703 -19268
rect 15767 -19332 15783 -19268
rect 15656 -19348 15783 -19332
rect 15656 -19412 15703 -19348
rect 15767 -19412 15783 -19348
rect 15656 -19428 15783 -19412
rect 15656 -19492 15703 -19428
rect 15767 -19492 15783 -19428
rect 15656 -19508 15783 -19492
rect 15656 -19572 15703 -19508
rect 15767 -19572 15783 -19508
rect 15656 -19588 15783 -19572
rect 15656 -19652 15703 -19588
rect 15767 -19652 15783 -19588
rect 15656 -19668 15783 -19652
rect 15656 -19732 15703 -19668
rect 15767 -19732 15783 -19668
rect 15656 -19748 15783 -19732
rect 15656 -19812 15703 -19748
rect 15767 -19812 15783 -19748
rect 15656 -19828 15783 -19812
rect 15656 -19892 15703 -19828
rect 15767 -19892 15783 -19828
rect 15656 -19908 15783 -19892
rect 15656 -19972 15703 -19908
rect 15767 -19972 15783 -19908
rect 15656 -19988 15783 -19972
rect 15656 -20052 15703 -19988
rect 15767 -20052 15783 -19988
rect 15656 -20068 15783 -20052
rect 15656 -20132 15703 -20068
rect 15767 -20132 15783 -20068
rect 15656 -20148 15783 -20132
rect 15656 -20212 15703 -20148
rect 15767 -20212 15783 -20148
rect 15656 -20228 15783 -20212
rect 15656 -20292 15703 -20228
rect 15767 -20292 15783 -20228
rect 15656 -20308 15783 -20292
rect 15656 -20372 15703 -20308
rect 15767 -20372 15783 -20308
rect 15656 -20388 15783 -20372
rect 15656 -20452 15703 -20388
rect 15767 -20452 15783 -20388
rect 15656 -20468 15783 -20452
rect 15656 -20532 15703 -20468
rect 15767 -20532 15783 -20468
rect 15656 -20548 15783 -20532
rect 15656 -20612 15703 -20548
rect 15767 -20612 15783 -20548
rect 15656 -20628 15783 -20612
rect 15656 -20692 15703 -20628
rect 15767 -20692 15783 -20628
rect 15656 -20708 15783 -20692
rect 15656 -20772 15703 -20708
rect 15767 -20772 15783 -20708
rect 15656 -20788 15783 -20772
rect 15656 -20852 15703 -20788
rect 15767 -20852 15783 -20788
rect 15656 -20868 15783 -20852
rect 15656 -20932 15703 -20868
rect 15767 -20932 15783 -20868
rect 15656 -20948 15783 -20932
rect 15656 -21012 15703 -20948
rect 15767 -21012 15783 -20948
rect 15656 -21028 15783 -21012
rect 15656 -21092 15703 -21028
rect 15767 -21092 15783 -21028
rect 15656 -21108 15783 -21092
rect 15656 -21172 15703 -21108
rect 15767 -21172 15783 -21108
rect 15656 -21188 15783 -21172
rect 15656 -21252 15703 -21188
rect 15767 -21252 15783 -21188
rect 15656 -21268 15783 -21252
rect 15656 -21332 15703 -21268
rect 15767 -21332 15783 -21268
rect 15656 -21348 15783 -21332
rect 15656 -21412 15703 -21348
rect 15767 -21412 15783 -21348
rect 15656 -21428 15783 -21412
rect 15656 -21492 15703 -21428
rect 15767 -21492 15783 -21428
rect 15656 -21508 15783 -21492
rect 15656 -21572 15703 -21508
rect 15767 -21572 15783 -21508
rect 15656 -21588 15783 -21572
rect 15656 -21652 15703 -21588
rect 15767 -21652 15783 -21588
rect 15656 -21668 15783 -21652
rect 15656 -21732 15703 -21668
rect 15767 -21732 15783 -21668
rect 15656 -21748 15783 -21732
rect 15656 -21812 15703 -21748
rect 15767 -21812 15783 -21748
rect 15656 -21828 15783 -21812
rect 9337 -21908 9464 -21892
rect 9337 -21972 9384 -21908
rect 9448 -21972 9464 -21908
rect 9337 -21988 9464 -21972
rect 9337 -22112 9441 -21988
rect 9337 -22128 9464 -22112
rect 9337 -22192 9384 -22128
rect 9448 -22192 9464 -22128
rect 9337 -22208 9464 -22192
rect 3018 -22288 3145 -22272
rect 3018 -22352 3065 -22288
rect 3129 -22352 3145 -22288
rect 3018 -22368 3145 -22352
rect 3018 -22432 3065 -22368
rect 3129 -22432 3145 -22368
rect 3018 -22448 3145 -22432
rect 3018 -22512 3065 -22448
rect 3129 -22512 3145 -22448
rect 3018 -22528 3145 -22512
rect 3018 -22592 3065 -22528
rect 3129 -22592 3145 -22528
rect 3018 -22608 3145 -22592
rect 3018 -22672 3065 -22608
rect 3129 -22672 3145 -22608
rect 3018 -22688 3145 -22672
rect 3018 -22752 3065 -22688
rect 3129 -22752 3145 -22688
rect 3018 -22768 3145 -22752
rect 3018 -22832 3065 -22768
rect 3129 -22832 3145 -22768
rect 3018 -22848 3145 -22832
rect 3018 -22912 3065 -22848
rect 3129 -22912 3145 -22848
rect 3018 -22928 3145 -22912
rect 3018 -22992 3065 -22928
rect 3129 -22992 3145 -22928
rect 3018 -23008 3145 -22992
rect 3018 -23072 3065 -23008
rect 3129 -23072 3145 -23008
rect 3018 -23088 3145 -23072
rect 3018 -23152 3065 -23088
rect 3129 -23152 3145 -23088
rect 3018 -23168 3145 -23152
rect 3018 -23232 3065 -23168
rect 3129 -23232 3145 -23168
rect 3018 -23248 3145 -23232
rect 3018 -23312 3065 -23248
rect 3129 -23312 3145 -23248
rect 3018 -23328 3145 -23312
rect 3018 -23392 3065 -23328
rect 3129 -23392 3145 -23328
rect 3018 -23408 3145 -23392
rect 3018 -23472 3065 -23408
rect 3129 -23472 3145 -23408
rect 3018 -23488 3145 -23472
rect 3018 -23552 3065 -23488
rect 3129 -23552 3145 -23488
rect 3018 -23568 3145 -23552
rect 3018 -23632 3065 -23568
rect 3129 -23632 3145 -23568
rect 3018 -23648 3145 -23632
rect 3018 -23712 3065 -23648
rect 3129 -23712 3145 -23648
rect 3018 -23728 3145 -23712
rect 3018 -23792 3065 -23728
rect 3129 -23792 3145 -23728
rect 3018 -23808 3145 -23792
rect 3018 -23872 3065 -23808
rect 3129 -23872 3145 -23808
rect 3018 -23888 3145 -23872
rect 3018 -23952 3065 -23888
rect 3129 -23952 3145 -23888
rect 3018 -23968 3145 -23952
rect 3018 -24032 3065 -23968
rect 3129 -24032 3145 -23968
rect 3018 -24048 3145 -24032
rect 3018 -24112 3065 -24048
rect 3129 -24112 3145 -24048
rect 3018 -24128 3145 -24112
rect 3018 -24192 3065 -24128
rect 3129 -24192 3145 -24128
rect 3018 -24208 3145 -24192
rect 3018 -24272 3065 -24208
rect 3129 -24272 3145 -24208
rect 3018 -24288 3145 -24272
rect 3018 -24352 3065 -24288
rect 3129 -24352 3145 -24288
rect 3018 -24368 3145 -24352
rect 3018 -24432 3065 -24368
rect 3129 -24432 3145 -24368
rect 3018 -24448 3145 -24432
rect 3018 -24512 3065 -24448
rect 3129 -24512 3145 -24448
rect 3018 -24528 3145 -24512
rect 3018 -24592 3065 -24528
rect 3129 -24592 3145 -24528
rect 3018 -24608 3145 -24592
rect 3018 -24672 3065 -24608
rect 3129 -24672 3145 -24608
rect 3018 -24688 3145 -24672
rect 3018 -24752 3065 -24688
rect 3129 -24752 3145 -24688
rect 3018 -24768 3145 -24752
rect 3018 -24832 3065 -24768
rect 3129 -24832 3145 -24768
rect 3018 -24848 3145 -24832
rect 3018 -24912 3065 -24848
rect 3129 -24912 3145 -24848
rect 3018 -24928 3145 -24912
rect 3018 -24992 3065 -24928
rect 3129 -24992 3145 -24928
rect 3018 -25008 3145 -24992
rect 3018 -25072 3065 -25008
rect 3129 -25072 3145 -25008
rect 3018 -25088 3145 -25072
rect 3018 -25152 3065 -25088
rect 3129 -25152 3145 -25088
rect 3018 -25168 3145 -25152
rect 3018 -25232 3065 -25168
rect 3129 -25232 3145 -25168
rect 3018 -25248 3145 -25232
rect 3018 -25312 3065 -25248
rect 3129 -25312 3145 -25248
rect 3018 -25328 3145 -25312
rect 3018 -25392 3065 -25328
rect 3129 -25392 3145 -25328
rect 3018 -25408 3145 -25392
rect 3018 -25472 3065 -25408
rect 3129 -25472 3145 -25408
rect 3018 -25488 3145 -25472
rect 3018 -25552 3065 -25488
rect 3129 -25552 3145 -25488
rect 3018 -25568 3145 -25552
rect 3018 -25632 3065 -25568
rect 3129 -25632 3145 -25568
rect 3018 -25648 3145 -25632
rect 3018 -25712 3065 -25648
rect 3129 -25712 3145 -25648
rect 3018 -25728 3145 -25712
rect 3018 -25792 3065 -25728
rect 3129 -25792 3145 -25728
rect 3018 -25808 3145 -25792
rect 3018 -25872 3065 -25808
rect 3129 -25872 3145 -25808
rect 3018 -25888 3145 -25872
rect 3018 -25952 3065 -25888
rect 3129 -25952 3145 -25888
rect 3018 -25968 3145 -25952
rect 3018 -26032 3065 -25968
rect 3129 -26032 3145 -25968
rect 3018 -26048 3145 -26032
rect 3018 -26112 3065 -26048
rect 3129 -26112 3145 -26048
rect 3018 -26128 3145 -26112
rect 3018 -26192 3065 -26128
rect 3129 -26192 3145 -26128
rect 3018 -26208 3145 -26192
rect 3018 -26272 3065 -26208
rect 3129 -26272 3145 -26208
rect 3018 -26288 3145 -26272
rect 3018 -26352 3065 -26288
rect 3129 -26352 3145 -26288
rect 3018 -26368 3145 -26352
rect 3018 -26432 3065 -26368
rect 3129 -26432 3145 -26368
rect 3018 -26448 3145 -26432
rect 3018 -26512 3065 -26448
rect 3129 -26512 3145 -26448
rect 3018 -26528 3145 -26512
rect 3018 -26592 3065 -26528
rect 3129 -26592 3145 -26528
rect 3018 -26608 3145 -26592
rect 3018 -26672 3065 -26608
rect 3129 -26672 3145 -26608
rect 3018 -26688 3145 -26672
rect 3018 -26752 3065 -26688
rect 3129 -26752 3145 -26688
rect 3018 -26768 3145 -26752
rect 3018 -26832 3065 -26768
rect 3129 -26832 3145 -26768
rect 3018 -26848 3145 -26832
rect 3018 -26912 3065 -26848
rect 3129 -26912 3145 -26848
rect 3018 -26928 3145 -26912
rect 3018 -26992 3065 -26928
rect 3129 -26992 3145 -26928
rect 3018 -27008 3145 -26992
rect 3018 -27072 3065 -27008
rect 3129 -27072 3145 -27008
rect 3018 -27088 3145 -27072
rect 3018 -27152 3065 -27088
rect 3129 -27152 3145 -27088
rect 3018 -27168 3145 -27152
rect 3018 -27232 3065 -27168
rect 3129 -27232 3145 -27168
rect 3018 -27248 3145 -27232
rect 3018 -27312 3065 -27248
rect 3129 -27312 3145 -27248
rect 3018 -27328 3145 -27312
rect 3018 -27392 3065 -27328
rect 3129 -27392 3145 -27328
rect 3018 -27408 3145 -27392
rect 3018 -27472 3065 -27408
rect 3129 -27472 3145 -27408
rect 3018 -27488 3145 -27472
rect 3018 -27552 3065 -27488
rect 3129 -27552 3145 -27488
rect 3018 -27568 3145 -27552
rect 3018 -27632 3065 -27568
rect 3129 -27632 3145 -27568
rect 3018 -27648 3145 -27632
rect 3018 -27712 3065 -27648
rect 3129 -27712 3145 -27648
rect 3018 -27728 3145 -27712
rect 3018 -27792 3065 -27728
rect 3129 -27792 3145 -27728
rect 3018 -27808 3145 -27792
rect 3018 -27872 3065 -27808
rect 3129 -27872 3145 -27808
rect 3018 -27888 3145 -27872
rect 3018 -27952 3065 -27888
rect 3129 -27952 3145 -27888
rect 3018 -27968 3145 -27952
rect 3018 -28032 3065 -27968
rect 3129 -28032 3145 -27968
rect 3018 -28048 3145 -28032
rect 3018 -28112 3065 -28048
rect 3129 -28112 3145 -28048
rect 3018 -28128 3145 -28112
rect -3301 -28208 -3174 -28192
rect -3301 -28272 -3254 -28208
rect -3190 -28272 -3174 -28208
rect -3301 -28288 -3174 -28272
rect -3301 -28412 -3197 -28288
rect -3301 -28428 -3174 -28412
rect -3301 -28492 -3254 -28428
rect -3190 -28492 -3174 -28428
rect -3301 -28508 -3174 -28492
rect -9620 -28588 -9493 -28572
rect -9620 -28652 -9573 -28588
rect -9509 -28652 -9493 -28588
rect -9620 -28668 -9493 -28652
rect -9620 -28732 -9573 -28668
rect -9509 -28732 -9493 -28668
rect -9620 -28748 -9493 -28732
rect -9620 -28812 -9573 -28748
rect -9509 -28812 -9493 -28748
rect -9620 -28828 -9493 -28812
rect -9620 -28892 -9573 -28828
rect -9509 -28892 -9493 -28828
rect -9620 -28908 -9493 -28892
rect -9620 -28972 -9573 -28908
rect -9509 -28972 -9493 -28908
rect -9620 -28988 -9493 -28972
rect -9620 -29052 -9573 -28988
rect -9509 -29052 -9493 -28988
rect -9620 -29068 -9493 -29052
rect -9620 -29132 -9573 -29068
rect -9509 -29132 -9493 -29068
rect -9620 -29148 -9493 -29132
rect -9620 -29212 -9573 -29148
rect -9509 -29212 -9493 -29148
rect -9620 -29228 -9493 -29212
rect -9620 -29292 -9573 -29228
rect -9509 -29292 -9493 -29228
rect -9620 -29308 -9493 -29292
rect -9620 -29372 -9573 -29308
rect -9509 -29372 -9493 -29308
rect -9620 -29388 -9493 -29372
rect -9620 -29452 -9573 -29388
rect -9509 -29452 -9493 -29388
rect -9620 -29468 -9493 -29452
rect -9620 -29532 -9573 -29468
rect -9509 -29532 -9493 -29468
rect -9620 -29548 -9493 -29532
rect -9620 -29612 -9573 -29548
rect -9509 -29612 -9493 -29548
rect -9620 -29628 -9493 -29612
rect -9620 -29692 -9573 -29628
rect -9509 -29692 -9493 -29628
rect -9620 -29708 -9493 -29692
rect -9620 -29772 -9573 -29708
rect -9509 -29772 -9493 -29708
rect -9620 -29788 -9493 -29772
rect -9620 -29852 -9573 -29788
rect -9509 -29852 -9493 -29788
rect -9620 -29868 -9493 -29852
rect -9620 -29932 -9573 -29868
rect -9509 -29932 -9493 -29868
rect -9620 -29948 -9493 -29932
rect -9620 -30012 -9573 -29948
rect -9509 -30012 -9493 -29948
rect -9620 -30028 -9493 -30012
rect -9620 -30092 -9573 -30028
rect -9509 -30092 -9493 -30028
rect -9620 -30108 -9493 -30092
rect -9620 -30172 -9573 -30108
rect -9509 -30172 -9493 -30108
rect -9620 -30188 -9493 -30172
rect -9620 -30252 -9573 -30188
rect -9509 -30252 -9493 -30188
rect -9620 -30268 -9493 -30252
rect -9620 -30332 -9573 -30268
rect -9509 -30332 -9493 -30268
rect -9620 -30348 -9493 -30332
rect -9620 -30412 -9573 -30348
rect -9509 -30412 -9493 -30348
rect -9620 -30428 -9493 -30412
rect -9620 -30492 -9573 -30428
rect -9509 -30492 -9493 -30428
rect -9620 -30508 -9493 -30492
rect -9620 -30572 -9573 -30508
rect -9509 -30572 -9493 -30508
rect -9620 -30588 -9493 -30572
rect -9620 -30652 -9573 -30588
rect -9509 -30652 -9493 -30588
rect -9620 -30668 -9493 -30652
rect -9620 -30732 -9573 -30668
rect -9509 -30732 -9493 -30668
rect -9620 -30748 -9493 -30732
rect -9620 -30812 -9573 -30748
rect -9509 -30812 -9493 -30748
rect -9620 -30828 -9493 -30812
rect -9620 -30892 -9573 -30828
rect -9509 -30892 -9493 -30828
rect -9620 -30908 -9493 -30892
rect -9620 -30972 -9573 -30908
rect -9509 -30972 -9493 -30908
rect -9620 -30988 -9493 -30972
rect -9620 -31052 -9573 -30988
rect -9509 -31052 -9493 -30988
rect -9620 -31068 -9493 -31052
rect -9620 -31132 -9573 -31068
rect -9509 -31132 -9493 -31068
rect -9620 -31148 -9493 -31132
rect -9620 -31212 -9573 -31148
rect -9509 -31212 -9493 -31148
rect -9620 -31228 -9493 -31212
rect -9620 -31292 -9573 -31228
rect -9509 -31292 -9493 -31228
rect -9620 -31308 -9493 -31292
rect -9620 -31372 -9573 -31308
rect -9509 -31372 -9493 -31308
rect -9620 -31388 -9493 -31372
rect -9620 -31452 -9573 -31388
rect -9509 -31452 -9493 -31388
rect -9620 -31468 -9493 -31452
rect -9620 -31532 -9573 -31468
rect -9509 -31532 -9493 -31468
rect -9620 -31548 -9493 -31532
rect -9620 -31612 -9573 -31548
rect -9509 -31612 -9493 -31548
rect -9620 -31628 -9493 -31612
rect -9620 -31692 -9573 -31628
rect -9509 -31692 -9493 -31628
rect -9620 -31708 -9493 -31692
rect -9620 -31772 -9573 -31708
rect -9509 -31772 -9493 -31708
rect -9620 -31788 -9493 -31772
rect -9620 -31852 -9573 -31788
rect -9509 -31852 -9493 -31788
rect -9620 -31868 -9493 -31852
rect -9620 -31932 -9573 -31868
rect -9509 -31932 -9493 -31868
rect -9620 -31948 -9493 -31932
rect -9620 -32012 -9573 -31948
rect -9509 -32012 -9493 -31948
rect -9620 -32028 -9493 -32012
rect -9620 -32092 -9573 -32028
rect -9509 -32092 -9493 -32028
rect -9620 -32108 -9493 -32092
rect -9620 -32172 -9573 -32108
rect -9509 -32172 -9493 -32108
rect -9620 -32188 -9493 -32172
rect -9620 -32252 -9573 -32188
rect -9509 -32252 -9493 -32188
rect -9620 -32268 -9493 -32252
rect -9620 -32332 -9573 -32268
rect -9509 -32332 -9493 -32268
rect -9620 -32348 -9493 -32332
rect -9620 -32412 -9573 -32348
rect -9509 -32412 -9493 -32348
rect -9620 -32428 -9493 -32412
rect -9620 -32492 -9573 -32428
rect -9509 -32492 -9493 -32428
rect -9620 -32508 -9493 -32492
rect -9620 -32572 -9573 -32508
rect -9509 -32572 -9493 -32508
rect -9620 -32588 -9493 -32572
rect -9620 -32652 -9573 -32588
rect -9509 -32652 -9493 -32588
rect -9620 -32668 -9493 -32652
rect -9620 -32732 -9573 -32668
rect -9509 -32732 -9493 -32668
rect -9620 -32748 -9493 -32732
rect -9620 -32812 -9573 -32748
rect -9509 -32812 -9493 -32748
rect -9620 -32828 -9493 -32812
rect -9620 -32892 -9573 -32828
rect -9509 -32892 -9493 -32828
rect -9620 -32908 -9493 -32892
rect -9620 -32972 -9573 -32908
rect -9509 -32972 -9493 -32908
rect -9620 -32988 -9493 -32972
rect -9620 -33052 -9573 -32988
rect -9509 -33052 -9493 -32988
rect -9620 -33068 -9493 -33052
rect -9620 -33132 -9573 -33068
rect -9509 -33132 -9493 -33068
rect -9620 -33148 -9493 -33132
rect -9620 -33212 -9573 -33148
rect -9509 -33212 -9493 -33148
rect -9620 -33228 -9493 -33212
rect -9620 -33292 -9573 -33228
rect -9509 -33292 -9493 -33228
rect -9620 -33308 -9493 -33292
rect -9620 -33372 -9573 -33308
rect -9509 -33372 -9493 -33308
rect -9620 -33388 -9493 -33372
rect -9620 -33452 -9573 -33388
rect -9509 -33452 -9493 -33388
rect -9620 -33468 -9493 -33452
rect -9620 -33532 -9573 -33468
rect -9509 -33532 -9493 -33468
rect -9620 -33548 -9493 -33532
rect -9620 -33612 -9573 -33548
rect -9509 -33612 -9493 -33548
rect -9620 -33628 -9493 -33612
rect -9620 -33692 -9573 -33628
rect -9509 -33692 -9493 -33628
rect -9620 -33708 -9493 -33692
rect -9620 -33772 -9573 -33708
rect -9509 -33772 -9493 -33708
rect -9620 -33788 -9493 -33772
rect -9620 -33852 -9573 -33788
rect -9509 -33852 -9493 -33788
rect -9620 -33868 -9493 -33852
rect -9620 -33932 -9573 -33868
rect -9509 -33932 -9493 -33868
rect -9620 -33948 -9493 -33932
rect -9620 -34012 -9573 -33948
rect -9509 -34012 -9493 -33948
rect -9620 -34028 -9493 -34012
rect -9620 -34092 -9573 -34028
rect -9509 -34092 -9493 -34028
rect -9620 -34108 -9493 -34092
rect -9620 -34172 -9573 -34108
rect -9509 -34172 -9493 -34108
rect -9620 -34188 -9493 -34172
rect -9620 -34252 -9573 -34188
rect -9509 -34252 -9493 -34188
rect -9620 -34268 -9493 -34252
rect -9620 -34332 -9573 -34268
rect -9509 -34332 -9493 -34268
rect -9620 -34348 -9493 -34332
rect -9620 -34412 -9573 -34348
rect -9509 -34412 -9493 -34348
rect -9620 -34428 -9493 -34412
rect -15939 -34508 -15812 -34492
rect -15939 -34572 -15892 -34508
rect -15828 -34572 -15812 -34508
rect -15939 -34588 -15812 -34572
rect -15939 -34712 -15835 -34588
rect -15939 -34728 -15812 -34712
rect -15939 -34792 -15892 -34728
rect -15828 -34792 -15812 -34728
rect -15939 -34808 -15812 -34792
rect -22258 -34888 -22131 -34872
rect -22258 -34952 -22211 -34888
rect -22147 -34952 -22131 -34888
rect -22258 -34968 -22131 -34952
rect -22258 -35032 -22211 -34968
rect -22147 -35032 -22131 -34968
rect -22258 -35048 -22131 -35032
rect -22258 -35112 -22211 -35048
rect -22147 -35112 -22131 -35048
rect -22258 -35128 -22131 -35112
rect -22258 -35192 -22211 -35128
rect -22147 -35192 -22131 -35128
rect -22258 -35208 -22131 -35192
rect -22258 -35272 -22211 -35208
rect -22147 -35272 -22131 -35208
rect -22258 -35288 -22131 -35272
rect -22258 -35352 -22211 -35288
rect -22147 -35352 -22131 -35288
rect -22258 -35368 -22131 -35352
rect -22258 -35432 -22211 -35368
rect -22147 -35432 -22131 -35368
rect -22258 -35448 -22131 -35432
rect -22258 -35512 -22211 -35448
rect -22147 -35512 -22131 -35448
rect -22258 -35528 -22131 -35512
rect -22258 -35592 -22211 -35528
rect -22147 -35592 -22131 -35528
rect -22258 -35608 -22131 -35592
rect -22258 -35672 -22211 -35608
rect -22147 -35672 -22131 -35608
rect -22258 -35688 -22131 -35672
rect -22258 -35752 -22211 -35688
rect -22147 -35752 -22131 -35688
rect -22258 -35768 -22131 -35752
rect -22258 -35832 -22211 -35768
rect -22147 -35832 -22131 -35768
rect -22258 -35848 -22131 -35832
rect -22258 -35912 -22211 -35848
rect -22147 -35912 -22131 -35848
rect -22258 -35928 -22131 -35912
rect -22258 -35992 -22211 -35928
rect -22147 -35992 -22131 -35928
rect -22258 -36008 -22131 -35992
rect -22258 -36072 -22211 -36008
rect -22147 -36072 -22131 -36008
rect -22258 -36088 -22131 -36072
rect -22258 -36152 -22211 -36088
rect -22147 -36152 -22131 -36088
rect -22258 -36168 -22131 -36152
rect -22258 -36232 -22211 -36168
rect -22147 -36232 -22131 -36168
rect -22258 -36248 -22131 -36232
rect -22258 -36312 -22211 -36248
rect -22147 -36312 -22131 -36248
rect -22258 -36328 -22131 -36312
rect -22258 -36392 -22211 -36328
rect -22147 -36392 -22131 -36328
rect -22258 -36408 -22131 -36392
rect -22258 -36472 -22211 -36408
rect -22147 -36472 -22131 -36408
rect -22258 -36488 -22131 -36472
rect -22258 -36552 -22211 -36488
rect -22147 -36552 -22131 -36488
rect -22258 -36568 -22131 -36552
rect -22258 -36632 -22211 -36568
rect -22147 -36632 -22131 -36568
rect -22258 -36648 -22131 -36632
rect -22258 -36712 -22211 -36648
rect -22147 -36712 -22131 -36648
rect -22258 -36728 -22131 -36712
rect -22258 -36792 -22211 -36728
rect -22147 -36792 -22131 -36728
rect -22258 -36808 -22131 -36792
rect -22258 -36872 -22211 -36808
rect -22147 -36872 -22131 -36808
rect -22258 -36888 -22131 -36872
rect -22258 -36952 -22211 -36888
rect -22147 -36952 -22131 -36888
rect -22258 -36968 -22131 -36952
rect -22258 -37032 -22211 -36968
rect -22147 -37032 -22131 -36968
rect -22258 -37048 -22131 -37032
rect -22258 -37112 -22211 -37048
rect -22147 -37112 -22131 -37048
rect -22258 -37128 -22131 -37112
rect -22258 -37192 -22211 -37128
rect -22147 -37192 -22131 -37128
rect -22258 -37208 -22131 -37192
rect -22258 -37272 -22211 -37208
rect -22147 -37272 -22131 -37208
rect -22258 -37288 -22131 -37272
rect -22258 -37352 -22211 -37288
rect -22147 -37352 -22131 -37288
rect -22258 -37368 -22131 -37352
rect -22258 -37432 -22211 -37368
rect -22147 -37432 -22131 -37368
rect -22258 -37448 -22131 -37432
rect -22258 -37512 -22211 -37448
rect -22147 -37512 -22131 -37448
rect -22258 -37528 -22131 -37512
rect -22258 -37592 -22211 -37528
rect -22147 -37592 -22131 -37528
rect -22258 -37608 -22131 -37592
rect -22258 -37672 -22211 -37608
rect -22147 -37672 -22131 -37608
rect -22258 -37688 -22131 -37672
rect -22258 -37752 -22211 -37688
rect -22147 -37752 -22131 -37688
rect -22258 -37768 -22131 -37752
rect -22258 -37832 -22211 -37768
rect -22147 -37832 -22131 -37768
rect -22258 -37848 -22131 -37832
rect -22258 -37912 -22211 -37848
rect -22147 -37912 -22131 -37848
rect -22258 -37928 -22131 -37912
rect -22258 -37992 -22211 -37928
rect -22147 -37992 -22131 -37928
rect -22258 -38008 -22131 -37992
rect -22258 -38072 -22211 -38008
rect -22147 -38072 -22131 -38008
rect -22258 -38088 -22131 -38072
rect -22258 -38152 -22211 -38088
rect -22147 -38152 -22131 -38088
rect -22258 -38168 -22131 -38152
rect -22258 -38232 -22211 -38168
rect -22147 -38232 -22131 -38168
rect -22258 -38248 -22131 -38232
rect -22258 -38312 -22211 -38248
rect -22147 -38312 -22131 -38248
rect -22258 -38328 -22131 -38312
rect -22258 -38392 -22211 -38328
rect -22147 -38392 -22131 -38328
rect -22258 -38408 -22131 -38392
rect -22258 -38472 -22211 -38408
rect -22147 -38472 -22131 -38408
rect -22258 -38488 -22131 -38472
rect -22258 -38552 -22211 -38488
rect -22147 -38552 -22131 -38488
rect -22258 -38568 -22131 -38552
rect -22258 -38632 -22211 -38568
rect -22147 -38632 -22131 -38568
rect -22258 -38648 -22131 -38632
rect -22258 -38712 -22211 -38648
rect -22147 -38712 -22131 -38648
rect -22258 -38728 -22131 -38712
rect -22258 -38792 -22211 -38728
rect -22147 -38792 -22131 -38728
rect -22258 -38808 -22131 -38792
rect -22258 -38872 -22211 -38808
rect -22147 -38872 -22131 -38808
rect -22258 -38888 -22131 -38872
rect -22258 -38952 -22211 -38888
rect -22147 -38952 -22131 -38888
rect -22258 -38968 -22131 -38952
rect -22258 -39032 -22211 -38968
rect -22147 -39032 -22131 -38968
rect -22258 -39048 -22131 -39032
rect -22258 -39112 -22211 -39048
rect -22147 -39112 -22131 -39048
rect -22258 -39128 -22131 -39112
rect -22258 -39192 -22211 -39128
rect -22147 -39192 -22131 -39128
rect -22258 -39208 -22131 -39192
rect -22258 -39272 -22211 -39208
rect -22147 -39272 -22131 -39208
rect -22258 -39288 -22131 -39272
rect -22258 -39352 -22211 -39288
rect -22147 -39352 -22131 -39288
rect -22258 -39368 -22131 -39352
rect -22258 -39432 -22211 -39368
rect -22147 -39432 -22131 -39368
rect -22258 -39448 -22131 -39432
rect -22258 -39512 -22211 -39448
rect -22147 -39512 -22131 -39448
rect -22258 -39528 -22131 -39512
rect -22258 -39592 -22211 -39528
rect -22147 -39592 -22131 -39528
rect -22258 -39608 -22131 -39592
rect -22258 -39672 -22211 -39608
rect -22147 -39672 -22131 -39608
rect -22258 -39688 -22131 -39672
rect -22258 -39752 -22211 -39688
rect -22147 -39752 -22131 -39688
rect -22258 -39768 -22131 -39752
rect -22258 -39832 -22211 -39768
rect -22147 -39832 -22131 -39768
rect -22258 -39848 -22131 -39832
rect -22258 -39912 -22211 -39848
rect -22147 -39912 -22131 -39848
rect -22258 -39928 -22131 -39912
rect -22258 -39992 -22211 -39928
rect -22147 -39992 -22131 -39928
rect -22258 -40008 -22131 -39992
rect -22258 -40072 -22211 -40008
rect -22147 -40072 -22131 -40008
rect -22258 -40088 -22131 -40072
rect -22258 -40152 -22211 -40088
rect -22147 -40152 -22131 -40088
rect -22258 -40168 -22131 -40152
rect -22258 -40232 -22211 -40168
rect -22147 -40232 -22131 -40168
rect -22258 -40248 -22131 -40232
rect -22258 -40312 -22211 -40248
rect -22147 -40312 -22131 -40248
rect -22258 -40328 -22131 -40312
rect -22258 -40392 -22211 -40328
rect -22147 -40392 -22131 -40328
rect -22258 -40408 -22131 -40392
rect -22258 -40472 -22211 -40408
rect -22147 -40472 -22131 -40408
rect -22258 -40488 -22131 -40472
rect -22258 -40552 -22211 -40488
rect -22147 -40552 -22131 -40488
rect -22258 -40568 -22131 -40552
rect -22258 -40632 -22211 -40568
rect -22147 -40632 -22131 -40568
rect -22258 -40648 -22131 -40632
rect -22258 -40712 -22211 -40648
rect -22147 -40712 -22131 -40648
rect -22258 -40728 -22131 -40712
rect -28577 -40808 -28450 -40792
rect -28577 -40872 -28530 -40808
rect -28466 -40872 -28450 -40808
rect -28577 -40888 -28450 -40872
rect -28577 -41012 -28473 -40888
rect -28577 -41028 -28450 -41012
rect -28577 -41092 -28530 -41028
rect -28466 -41092 -28450 -41028
rect -28577 -41108 -28450 -41092
rect -34896 -41188 -34769 -41172
rect -34896 -41252 -34849 -41188
rect -34785 -41252 -34769 -41188
rect -34896 -41268 -34769 -41252
rect -34896 -41332 -34849 -41268
rect -34785 -41332 -34769 -41268
rect -34896 -41348 -34769 -41332
rect -34896 -41412 -34849 -41348
rect -34785 -41412 -34769 -41348
rect -34896 -41428 -34769 -41412
rect -34896 -41492 -34849 -41428
rect -34785 -41492 -34769 -41428
rect -34896 -41508 -34769 -41492
rect -34896 -41572 -34849 -41508
rect -34785 -41572 -34769 -41508
rect -34896 -41588 -34769 -41572
rect -34896 -41652 -34849 -41588
rect -34785 -41652 -34769 -41588
rect -34896 -41668 -34769 -41652
rect -34896 -41732 -34849 -41668
rect -34785 -41732 -34769 -41668
rect -34896 -41748 -34769 -41732
rect -34896 -41812 -34849 -41748
rect -34785 -41812 -34769 -41748
rect -34896 -41828 -34769 -41812
rect -34896 -41892 -34849 -41828
rect -34785 -41892 -34769 -41828
rect -34896 -41908 -34769 -41892
rect -34896 -41972 -34849 -41908
rect -34785 -41972 -34769 -41908
rect -34896 -41988 -34769 -41972
rect -34896 -42052 -34849 -41988
rect -34785 -42052 -34769 -41988
rect -34896 -42068 -34769 -42052
rect -34896 -42132 -34849 -42068
rect -34785 -42132 -34769 -42068
rect -34896 -42148 -34769 -42132
rect -34896 -42212 -34849 -42148
rect -34785 -42212 -34769 -42148
rect -34896 -42228 -34769 -42212
rect -34896 -42292 -34849 -42228
rect -34785 -42292 -34769 -42228
rect -34896 -42308 -34769 -42292
rect -34896 -42372 -34849 -42308
rect -34785 -42372 -34769 -42308
rect -34896 -42388 -34769 -42372
rect -34896 -42452 -34849 -42388
rect -34785 -42452 -34769 -42388
rect -34896 -42468 -34769 -42452
rect -34896 -42532 -34849 -42468
rect -34785 -42532 -34769 -42468
rect -34896 -42548 -34769 -42532
rect -34896 -42612 -34849 -42548
rect -34785 -42612 -34769 -42548
rect -34896 -42628 -34769 -42612
rect -34896 -42692 -34849 -42628
rect -34785 -42692 -34769 -42628
rect -34896 -42708 -34769 -42692
rect -34896 -42772 -34849 -42708
rect -34785 -42772 -34769 -42708
rect -34896 -42788 -34769 -42772
rect -34896 -42852 -34849 -42788
rect -34785 -42852 -34769 -42788
rect -34896 -42868 -34769 -42852
rect -34896 -42932 -34849 -42868
rect -34785 -42932 -34769 -42868
rect -34896 -42948 -34769 -42932
rect -34896 -43012 -34849 -42948
rect -34785 -43012 -34769 -42948
rect -34896 -43028 -34769 -43012
rect -34896 -43092 -34849 -43028
rect -34785 -43092 -34769 -43028
rect -34896 -43108 -34769 -43092
rect -34896 -43172 -34849 -43108
rect -34785 -43172 -34769 -43108
rect -34896 -43188 -34769 -43172
rect -34896 -43252 -34849 -43188
rect -34785 -43252 -34769 -43188
rect -34896 -43268 -34769 -43252
rect -34896 -43332 -34849 -43268
rect -34785 -43332 -34769 -43268
rect -34896 -43348 -34769 -43332
rect -34896 -43412 -34849 -43348
rect -34785 -43412 -34769 -43348
rect -34896 -43428 -34769 -43412
rect -34896 -43492 -34849 -43428
rect -34785 -43492 -34769 -43428
rect -34896 -43508 -34769 -43492
rect -34896 -43572 -34849 -43508
rect -34785 -43572 -34769 -43508
rect -34896 -43588 -34769 -43572
rect -34896 -43652 -34849 -43588
rect -34785 -43652 -34769 -43588
rect -34896 -43668 -34769 -43652
rect -34896 -43732 -34849 -43668
rect -34785 -43732 -34769 -43668
rect -34896 -43748 -34769 -43732
rect -34896 -43812 -34849 -43748
rect -34785 -43812 -34769 -43748
rect -34896 -43828 -34769 -43812
rect -34896 -43892 -34849 -43828
rect -34785 -43892 -34769 -43828
rect -34896 -43908 -34769 -43892
rect -34896 -43972 -34849 -43908
rect -34785 -43972 -34769 -43908
rect -34896 -43988 -34769 -43972
rect -34896 -44052 -34849 -43988
rect -34785 -44052 -34769 -43988
rect -34896 -44068 -34769 -44052
rect -34896 -44132 -34849 -44068
rect -34785 -44132 -34769 -44068
rect -34896 -44148 -34769 -44132
rect -34896 -44212 -34849 -44148
rect -34785 -44212 -34769 -44148
rect -34896 -44228 -34769 -44212
rect -34896 -44292 -34849 -44228
rect -34785 -44292 -34769 -44228
rect -34896 -44308 -34769 -44292
rect -34896 -44372 -34849 -44308
rect -34785 -44372 -34769 -44308
rect -34896 -44388 -34769 -44372
rect -34896 -44452 -34849 -44388
rect -34785 -44452 -34769 -44388
rect -34896 -44468 -34769 -44452
rect -34896 -44532 -34849 -44468
rect -34785 -44532 -34769 -44468
rect -34896 -44548 -34769 -44532
rect -34896 -44612 -34849 -44548
rect -34785 -44612 -34769 -44548
rect -34896 -44628 -34769 -44612
rect -34896 -44692 -34849 -44628
rect -34785 -44692 -34769 -44628
rect -34896 -44708 -34769 -44692
rect -34896 -44772 -34849 -44708
rect -34785 -44772 -34769 -44708
rect -34896 -44788 -34769 -44772
rect -34896 -44852 -34849 -44788
rect -34785 -44852 -34769 -44788
rect -34896 -44868 -34769 -44852
rect -34896 -44932 -34849 -44868
rect -34785 -44932 -34769 -44868
rect -34896 -44948 -34769 -44932
rect -34896 -45012 -34849 -44948
rect -34785 -45012 -34769 -44948
rect -34896 -45028 -34769 -45012
rect -34896 -45092 -34849 -45028
rect -34785 -45092 -34769 -45028
rect -34896 -45108 -34769 -45092
rect -34896 -45172 -34849 -45108
rect -34785 -45172 -34769 -45108
rect -34896 -45188 -34769 -45172
rect -34896 -45252 -34849 -45188
rect -34785 -45252 -34769 -45188
rect -34896 -45268 -34769 -45252
rect -34896 -45332 -34849 -45268
rect -34785 -45332 -34769 -45268
rect -34896 -45348 -34769 -45332
rect -34896 -45412 -34849 -45348
rect -34785 -45412 -34769 -45348
rect -34896 -45428 -34769 -45412
rect -34896 -45492 -34849 -45428
rect -34785 -45492 -34769 -45428
rect -34896 -45508 -34769 -45492
rect -34896 -45572 -34849 -45508
rect -34785 -45572 -34769 -45508
rect -34896 -45588 -34769 -45572
rect -34896 -45652 -34849 -45588
rect -34785 -45652 -34769 -45588
rect -34896 -45668 -34769 -45652
rect -34896 -45732 -34849 -45668
rect -34785 -45732 -34769 -45668
rect -34896 -45748 -34769 -45732
rect -34896 -45812 -34849 -45748
rect -34785 -45812 -34769 -45748
rect -34896 -45828 -34769 -45812
rect -34896 -45892 -34849 -45828
rect -34785 -45892 -34769 -45828
rect -34896 -45908 -34769 -45892
rect -34896 -45972 -34849 -45908
rect -34785 -45972 -34769 -45908
rect -34896 -45988 -34769 -45972
rect -34896 -46052 -34849 -45988
rect -34785 -46052 -34769 -45988
rect -34896 -46068 -34769 -46052
rect -34896 -46132 -34849 -46068
rect -34785 -46132 -34769 -46068
rect -34896 -46148 -34769 -46132
rect -34896 -46212 -34849 -46148
rect -34785 -46212 -34769 -46148
rect -34896 -46228 -34769 -46212
rect -34896 -46292 -34849 -46228
rect -34785 -46292 -34769 -46228
rect -34896 -46308 -34769 -46292
rect -34896 -46372 -34849 -46308
rect -34785 -46372 -34769 -46308
rect -34896 -46388 -34769 -46372
rect -34896 -46452 -34849 -46388
rect -34785 -46452 -34769 -46388
rect -34896 -46468 -34769 -46452
rect -34896 -46532 -34849 -46468
rect -34785 -46532 -34769 -46468
rect -34896 -46548 -34769 -46532
rect -34896 -46612 -34849 -46548
rect -34785 -46612 -34769 -46548
rect -34896 -46628 -34769 -46612
rect -34896 -46692 -34849 -46628
rect -34785 -46692 -34769 -46628
rect -34896 -46708 -34769 -46692
rect -34896 -46772 -34849 -46708
rect -34785 -46772 -34769 -46708
rect -34896 -46788 -34769 -46772
rect -34896 -46852 -34849 -46788
rect -34785 -46852 -34769 -46788
rect -34896 -46868 -34769 -46852
rect -34896 -46932 -34849 -46868
rect -34785 -46932 -34769 -46868
rect -34896 -46948 -34769 -46932
rect -34896 -47012 -34849 -46948
rect -34785 -47012 -34769 -46948
rect -34896 -47028 -34769 -47012
rect -41215 -47108 -41088 -47092
rect -41215 -47172 -41168 -47108
rect -41104 -47172 -41088 -47108
rect -41215 -47188 -41088 -47172
rect -41215 -47250 -41111 -47188
rect -38016 -47250 -37912 -47061
rect -34896 -47092 -34849 -47028
rect -34785 -47092 -34769 -47028
rect -34606 -41148 -28684 -41139
rect -34606 -47052 -34597 -41148
rect -28693 -47052 -28684 -41148
rect -34606 -47061 -28684 -47052
rect -28577 -41172 -28530 -41108
rect -28466 -41172 -28450 -41108
rect -25378 -41139 -25274 -40761
rect -22258 -40792 -22211 -40728
rect -22147 -40792 -22131 -40728
rect -21968 -34848 -16046 -34839
rect -21968 -40752 -21959 -34848
rect -16055 -40752 -16046 -34848
rect -21968 -40761 -16046 -40752
rect -15939 -34872 -15892 -34808
rect -15828 -34872 -15812 -34808
rect -12740 -34839 -12636 -34461
rect -9620 -34492 -9573 -34428
rect -9509 -34492 -9493 -34428
rect -9330 -28548 -3408 -28539
rect -9330 -34452 -9321 -28548
rect -3417 -34452 -3408 -28548
rect -9330 -34461 -3408 -34452
rect -3301 -28572 -3254 -28508
rect -3190 -28572 -3174 -28508
rect -102 -28539 2 -28161
rect 3018 -28192 3065 -28128
rect 3129 -28192 3145 -28128
rect 3308 -22248 9230 -22239
rect 3308 -28152 3317 -22248
rect 9221 -28152 9230 -22248
rect 3308 -28161 9230 -28152
rect 9337 -22272 9384 -22208
rect 9448 -22272 9464 -22208
rect 12536 -22239 12640 -21861
rect 15656 -21892 15703 -21828
rect 15767 -21892 15783 -21828
rect 15946 -15948 21868 -15939
rect 15946 -21852 15955 -15948
rect 21859 -21852 21868 -15948
rect 15946 -21861 21868 -21852
rect 21975 -15972 22022 -15908
rect 22086 -15972 22102 -15908
rect 25174 -15939 25278 -15561
rect 28294 -15592 28341 -15528
rect 28405 -15592 28421 -15528
rect 28584 -9648 34506 -9639
rect 28584 -15552 28593 -9648
rect 34497 -15552 34506 -9648
rect 28584 -15561 34506 -15552
rect 34613 -9672 34660 -9608
rect 34724 -9672 34740 -9608
rect 37812 -9639 37916 -9261
rect 40932 -9292 40979 -9228
rect 41043 -9292 41059 -9228
rect 41222 -3348 47144 -3339
rect 41222 -9252 41231 -3348
rect 47135 -9252 47144 -3348
rect 41222 -9261 47144 -9252
rect 47251 -3372 47298 -3308
rect 47362 -3372 47378 -3308
rect 47251 -3388 47378 -3372
rect 47251 -3452 47298 -3388
rect 47362 -3452 47378 -3388
rect 47251 -3468 47378 -3452
rect 47251 -3532 47298 -3468
rect 47362 -3532 47378 -3468
rect 47251 -3548 47378 -3532
rect 47251 -3612 47298 -3548
rect 47362 -3612 47378 -3548
rect 47251 -3628 47378 -3612
rect 47251 -3692 47298 -3628
rect 47362 -3692 47378 -3628
rect 47251 -3708 47378 -3692
rect 47251 -3772 47298 -3708
rect 47362 -3772 47378 -3708
rect 47251 -3788 47378 -3772
rect 47251 -3852 47298 -3788
rect 47362 -3852 47378 -3788
rect 47251 -3868 47378 -3852
rect 47251 -3932 47298 -3868
rect 47362 -3932 47378 -3868
rect 47251 -3948 47378 -3932
rect 47251 -4012 47298 -3948
rect 47362 -4012 47378 -3948
rect 47251 -4028 47378 -4012
rect 47251 -4092 47298 -4028
rect 47362 -4092 47378 -4028
rect 47251 -4108 47378 -4092
rect 47251 -4172 47298 -4108
rect 47362 -4172 47378 -4108
rect 47251 -4188 47378 -4172
rect 47251 -4252 47298 -4188
rect 47362 -4252 47378 -4188
rect 47251 -4268 47378 -4252
rect 47251 -4332 47298 -4268
rect 47362 -4332 47378 -4268
rect 47251 -4348 47378 -4332
rect 47251 -4412 47298 -4348
rect 47362 -4412 47378 -4348
rect 47251 -4428 47378 -4412
rect 47251 -4492 47298 -4428
rect 47362 -4492 47378 -4428
rect 47251 -4508 47378 -4492
rect 47251 -4572 47298 -4508
rect 47362 -4572 47378 -4508
rect 47251 -4588 47378 -4572
rect 47251 -4652 47298 -4588
rect 47362 -4652 47378 -4588
rect 47251 -4668 47378 -4652
rect 47251 -4732 47298 -4668
rect 47362 -4732 47378 -4668
rect 47251 -4748 47378 -4732
rect 47251 -4812 47298 -4748
rect 47362 -4812 47378 -4748
rect 47251 -4828 47378 -4812
rect 47251 -4892 47298 -4828
rect 47362 -4892 47378 -4828
rect 47251 -4908 47378 -4892
rect 47251 -4972 47298 -4908
rect 47362 -4972 47378 -4908
rect 47251 -4988 47378 -4972
rect 47251 -5052 47298 -4988
rect 47362 -5052 47378 -4988
rect 47251 -5068 47378 -5052
rect 47251 -5132 47298 -5068
rect 47362 -5132 47378 -5068
rect 47251 -5148 47378 -5132
rect 47251 -5212 47298 -5148
rect 47362 -5212 47378 -5148
rect 47251 -5228 47378 -5212
rect 47251 -5292 47298 -5228
rect 47362 -5292 47378 -5228
rect 47251 -5308 47378 -5292
rect 47251 -5372 47298 -5308
rect 47362 -5372 47378 -5308
rect 47251 -5388 47378 -5372
rect 47251 -5452 47298 -5388
rect 47362 -5452 47378 -5388
rect 47251 -5468 47378 -5452
rect 47251 -5532 47298 -5468
rect 47362 -5532 47378 -5468
rect 47251 -5548 47378 -5532
rect 47251 -5612 47298 -5548
rect 47362 -5612 47378 -5548
rect 47251 -5628 47378 -5612
rect 47251 -5692 47298 -5628
rect 47362 -5692 47378 -5628
rect 47251 -5708 47378 -5692
rect 47251 -5772 47298 -5708
rect 47362 -5772 47378 -5708
rect 47251 -5788 47378 -5772
rect 47251 -5852 47298 -5788
rect 47362 -5852 47378 -5788
rect 47251 -5868 47378 -5852
rect 47251 -5932 47298 -5868
rect 47362 -5932 47378 -5868
rect 47251 -5948 47378 -5932
rect 47251 -6012 47298 -5948
rect 47362 -6012 47378 -5948
rect 47251 -6028 47378 -6012
rect 47251 -6092 47298 -6028
rect 47362 -6092 47378 -6028
rect 47251 -6108 47378 -6092
rect 47251 -6172 47298 -6108
rect 47362 -6172 47378 -6108
rect 47251 -6188 47378 -6172
rect 47251 -6252 47298 -6188
rect 47362 -6252 47378 -6188
rect 47251 -6268 47378 -6252
rect 47251 -6332 47298 -6268
rect 47362 -6332 47378 -6268
rect 47251 -6348 47378 -6332
rect 47251 -6412 47298 -6348
rect 47362 -6412 47378 -6348
rect 47251 -6428 47378 -6412
rect 47251 -6492 47298 -6428
rect 47362 -6492 47378 -6428
rect 47251 -6508 47378 -6492
rect 47251 -6572 47298 -6508
rect 47362 -6572 47378 -6508
rect 47251 -6588 47378 -6572
rect 47251 -6652 47298 -6588
rect 47362 -6652 47378 -6588
rect 47251 -6668 47378 -6652
rect 47251 -6732 47298 -6668
rect 47362 -6732 47378 -6668
rect 47251 -6748 47378 -6732
rect 47251 -6812 47298 -6748
rect 47362 -6812 47378 -6748
rect 47251 -6828 47378 -6812
rect 47251 -6892 47298 -6828
rect 47362 -6892 47378 -6828
rect 47251 -6908 47378 -6892
rect 47251 -6972 47298 -6908
rect 47362 -6972 47378 -6908
rect 47251 -6988 47378 -6972
rect 47251 -7052 47298 -6988
rect 47362 -7052 47378 -6988
rect 47251 -7068 47378 -7052
rect 47251 -7132 47298 -7068
rect 47362 -7132 47378 -7068
rect 47251 -7148 47378 -7132
rect 47251 -7212 47298 -7148
rect 47362 -7212 47378 -7148
rect 47251 -7228 47378 -7212
rect 47251 -7292 47298 -7228
rect 47362 -7292 47378 -7228
rect 47251 -7308 47378 -7292
rect 47251 -7372 47298 -7308
rect 47362 -7372 47378 -7308
rect 47251 -7388 47378 -7372
rect 47251 -7452 47298 -7388
rect 47362 -7452 47378 -7388
rect 47251 -7468 47378 -7452
rect 47251 -7532 47298 -7468
rect 47362 -7532 47378 -7468
rect 47251 -7548 47378 -7532
rect 47251 -7612 47298 -7548
rect 47362 -7612 47378 -7548
rect 47251 -7628 47378 -7612
rect 47251 -7692 47298 -7628
rect 47362 -7692 47378 -7628
rect 47251 -7708 47378 -7692
rect 47251 -7772 47298 -7708
rect 47362 -7772 47378 -7708
rect 47251 -7788 47378 -7772
rect 47251 -7852 47298 -7788
rect 47362 -7852 47378 -7788
rect 47251 -7868 47378 -7852
rect 47251 -7932 47298 -7868
rect 47362 -7932 47378 -7868
rect 47251 -7948 47378 -7932
rect 47251 -8012 47298 -7948
rect 47362 -8012 47378 -7948
rect 47251 -8028 47378 -8012
rect 47251 -8092 47298 -8028
rect 47362 -8092 47378 -8028
rect 47251 -8108 47378 -8092
rect 47251 -8172 47298 -8108
rect 47362 -8172 47378 -8108
rect 47251 -8188 47378 -8172
rect 47251 -8252 47298 -8188
rect 47362 -8252 47378 -8188
rect 47251 -8268 47378 -8252
rect 47251 -8332 47298 -8268
rect 47362 -8332 47378 -8268
rect 47251 -8348 47378 -8332
rect 47251 -8412 47298 -8348
rect 47362 -8412 47378 -8348
rect 47251 -8428 47378 -8412
rect 47251 -8492 47298 -8428
rect 47362 -8492 47378 -8428
rect 47251 -8508 47378 -8492
rect 47251 -8572 47298 -8508
rect 47362 -8572 47378 -8508
rect 47251 -8588 47378 -8572
rect 47251 -8652 47298 -8588
rect 47362 -8652 47378 -8588
rect 47251 -8668 47378 -8652
rect 47251 -8732 47298 -8668
rect 47362 -8732 47378 -8668
rect 47251 -8748 47378 -8732
rect 47251 -8812 47298 -8748
rect 47362 -8812 47378 -8748
rect 47251 -8828 47378 -8812
rect 47251 -8892 47298 -8828
rect 47362 -8892 47378 -8828
rect 47251 -8908 47378 -8892
rect 47251 -8972 47298 -8908
rect 47362 -8972 47378 -8908
rect 47251 -8988 47378 -8972
rect 47251 -9052 47298 -8988
rect 47362 -9052 47378 -8988
rect 47251 -9068 47378 -9052
rect 47251 -9132 47298 -9068
rect 47362 -9132 47378 -9068
rect 47251 -9148 47378 -9132
rect 47251 -9212 47298 -9148
rect 47362 -9212 47378 -9148
rect 47251 -9228 47378 -9212
rect 40932 -9308 41059 -9292
rect 40932 -9372 40979 -9308
rect 41043 -9372 41059 -9308
rect 40932 -9388 41059 -9372
rect 40932 -9512 41036 -9388
rect 40932 -9528 41059 -9512
rect 40932 -9592 40979 -9528
rect 41043 -9592 41059 -9528
rect 40932 -9608 41059 -9592
rect 34613 -9688 34740 -9672
rect 34613 -9752 34660 -9688
rect 34724 -9752 34740 -9688
rect 34613 -9768 34740 -9752
rect 34613 -9832 34660 -9768
rect 34724 -9832 34740 -9768
rect 34613 -9848 34740 -9832
rect 34613 -9912 34660 -9848
rect 34724 -9912 34740 -9848
rect 34613 -9928 34740 -9912
rect 34613 -9992 34660 -9928
rect 34724 -9992 34740 -9928
rect 34613 -10008 34740 -9992
rect 34613 -10072 34660 -10008
rect 34724 -10072 34740 -10008
rect 34613 -10088 34740 -10072
rect 34613 -10152 34660 -10088
rect 34724 -10152 34740 -10088
rect 34613 -10168 34740 -10152
rect 34613 -10232 34660 -10168
rect 34724 -10232 34740 -10168
rect 34613 -10248 34740 -10232
rect 34613 -10312 34660 -10248
rect 34724 -10312 34740 -10248
rect 34613 -10328 34740 -10312
rect 34613 -10392 34660 -10328
rect 34724 -10392 34740 -10328
rect 34613 -10408 34740 -10392
rect 34613 -10472 34660 -10408
rect 34724 -10472 34740 -10408
rect 34613 -10488 34740 -10472
rect 34613 -10552 34660 -10488
rect 34724 -10552 34740 -10488
rect 34613 -10568 34740 -10552
rect 34613 -10632 34660 -10568
rect 34724 -10632 34740 -10568
rect 34613 -10648 34740 -10632
rect 34613 -10712 34660 -10648
rect 34724 -10712 34740 -10648
rect 34613 -10728 34740 -10712
rect 34613 -10792 34660 -10728
rect 34724 -10792 34740 -10728
rect 34613 -10808 34740 -10792
rect 34613 -10872 34660 -10808
rect 34724 -10872 34740 -10808
rect 34613 -10888 34740 -10872
rect 34613 -10952 34660 -10888
rect 34724 -10952 34740 -10888
rect 34613 -10968 34740 -10952
rect 34613 -11032 34660 -10968
rect 34724 -11032 34740 -10968
rect 34613 -11048 34740 -11032
rect 34613 -11112 34660 -11048
rect 34724 -11112 34740 -11048
rect 34613 -11128 34740 -11112
rect 34613 -11192 34660 -11128
rect 34724 -11192 34740 -11128
rect 34613 -11208 34740 -11192
rect 34613 -11272 34660 -11208
rect 34724 -11272 34740 -11208
rect 34613 -11288 34740 -11272
rect 34613 -11352 34660 -11288
rect 34724 -11352 34740 -11288
rect 34613 -11368 34740 -11352
rect 34613 -11432 34660 -11368
rect 34724 -11432 34740 -11368
rect 34613 -11448 34740 -11432
rect 34613 -11512 34660 -11448
rect 34724 -11512 34740 -11448
rect 34613 -11528 34740 -11512
rect 34613 -11592 34660 -11528
rect 34724 -11592 34740 -11528
rect 34613 -11608 34740 -11592
rect 34613 -11672 34660 -11608
rect 34724 -11672 34740 -11608
rect 34613 -11688 34740 -11672
rect 34613 -11752 34660 -11688
rect 34724 -11752 34740 -11688
rect 34613 -11768 34740 -11752
rect 34613 -11832 34660 -11768
rect 34724 -11832 34740 -11768
rect 34613 -11848 34740 -11832
rect 34613 -11912 34660 -11848
rect 34724 -11912 34740 -11848
rect 34613 -11928 34740 -11912
rect 34613 -11992 34660 -11928
rect 34724 -11992 34740 -11928
rect 34613 -12008 34740 -11992
rect 34613 -12072 34660 -12008
rect 34724 -12072 34740 -12008
rect 34613 -12088 34740 -12072
rect 34613 -12152 34660 -12088
rect 34724 -12152 34740 -12088
rect 34613 -12168 34740 -12152
rect 34613 -12232 34660 -12168
rect 34724 -12232 34740 -12168
rect 34613 -12248 34740 -12232
rect 34613 -12312 34660 -12248
rect 34724 -12312 34740 -12248
rect 34613 -12328 34740 -12312
rect 34613 -12392 34660 -12328
rect 34724 -12392 34740 -12328
rect 34613 -12408 34740 -12392
rect 34613 -12472 34660 -12408
rect 34724 -12472 34740 -12408
rect 34613 -12488 34740 -12472
rect 34613 -12552 34660 -12488
rect 34724 -12552 34740 -12488
rect 34613 -12568 34740 -12552
rect 34613 -12632 34660 -12568
rect 34724 -12632 34740 -12568
rect 34613 -12648 34740 -12632
rect 34613 -12712 34660 -12648
rect 34724 -12712 34740 -12648
rect 34613 -12728 34740 -12712
rect 34613 -12792 34660 -12728
rect 34724 -12792 34740 -12728
rect 34613 -12808 34740 -12792
rect 34613 -12872 34660 -12808
rect 34724 -12872 34740 -12808
rect 34613 -12888 34740 -12872
rect 34613 -12952 34660 -12888
rect 34724 -12952 34740 -12888
rect 34613 -12968 34740 -12952
rect 34613 -13032 34660 -12968
rect 34724 -13032 34740 -12968
rect 34613 -13048 34740 -13032
rect 34613 -13112 34660 -13048
rect 34724 -13112 34740 -13048
rect 34613 -13128 34740 -13112
rect 34613 -13192 34660 -13128
rect 34724 -13192 34740 -13128
rect 34613 -13208 34740 -13192
rect 34613 -13272 34660 -13208
rect 34724 -13272 34740 -13208
rect 34613 -13288 34740 -13272
rect 34613 -13352 34660 -13288
rect 34724 -13352 34740 -13288
rect 34613 -13368 34740 -13352
rect 34613 -13432 34660 -13368
rect 34724 -13432 34740 -13368
rect 34613 -13448 34740 -13432
rect 34613 -13512 34660 -13448
rect 34724 -13512 34740 -13448
rect 34613 -13528 34740 -13512
rect 34613 -13592 34660 -13528
rect 34724 -13592 34740 -13528
rect 34613 -13608 34740 -13592
rect 34613 -13672 34660 -13608
rect 34724 -13672 34740 -13608
rect 34613 -13688 34740 -13672
rect 34613 -13752 34660 -13688
rect 34724 -13752 34740 -13688
rect 34613 -13768 34740 -13752
rect 34613 -13832 34660 -13768
rect 34724 -13832 34740 -13768
rect 34613 -13848 34740 -13832
rect 34613 -13912 34660 -13848
rect 34724 -13912 34740 -13848
rect 34613 -13928 34740 -13912
rect 34613 -13992 34660 -13928
rect 34724 -13992 34740 -13928
rect 34613 -14008 34740 -13992
rect 34613 -14072 34660 -14008
rect 34724 -14072 34740 -14008
rect 34613 -14088 34740 -14072
rect 34613 -14152 34660 -14088
rect 34724 -14152 34740 -14088
rect 34613 -14168 34740 -14152
rect 34613 -14232 34660 -14168
rect 34724 -14232 34740 -14168
rect 34613 -14248 34740 -14232
rect 34613 -14312 34660 -14248
rect 34724 -14312 34740 -14248
rect 34613 -14328 34740 -14312
rect 34613 -14392 34660 -14328
rect 34724 -14392 34740 -14328
rect 34613 -14408 34740 -14392
rect 34613 -14472 34660 -14408
rect 34724 -14472 34740 -14408
rect 34613 -14488 34740 -14472
rect 34613 -14552 34660 -14488
rect 34724 -14552 34740 -14488
rect 34613 -14568 34740 -14552
rect 34613 -14632 34660 -14568
rect 34724 -14632 34740 -14568
rect 34613 -14648 34740 -14632
rect 34613 -14712 34660 -14648
rect 34724 -14712 34740 -14648
rect 34613 -14728 34740 -14712
rect 34613 -14792 34660 -14728
rect 34724 -14792 34740 -14728
rect 34613 -14808 34740 -14792
rect 34613 -14872 34660 -14808
rect 34724 -14872 34740 -14808
rect 34613 -14888 34740 -14872
rect 34613 -14952 34660 -14888
rect 34724 -14952 34740 -14888
rect 34613 -14968 34740 -14952
rect 34613 -15032 34660 -14968
rect 34724 -15032 34740 -14968
rect 34613 -15048 34740 -15032
rect 34613 -15112 34660 -15048
rect 34724 -15112 34740 -15048
rect 34613 -15128 34740 -15112
rect 34613 -15192 34660 -15128
rect 34724 -15192 34740 -15128
rect 34613 -15208 34740 -15192
rect 34613 -15272 34660 -15208
rect 34724 -15272 34740 -15208
rect 34613 -15288 34740 -15272
rect 34613 -15352 34660 -15288
rect 34724 -15352 34740 -15288
rect 34613 -15368 34740 -15352
rect 34613 -15432 34660 -15368
rect 34724 -15432 34740 -15368
rect 34613 -15448 34740 -15432
rect 34613 -15512 34660 -15448
rect 34724 -15512 34740 -15448
rect 34613 -15528 34740 -15512
rect 28294 -15608 28421 -15592
rect 28294 -15672 28341 -15608
rect 28405 -15672 28421 -15608
rect 28294 -15688 28421 -15672
rect 28294 -15812 28398 -15688
rect 28294 -15828 28421 -15812
rect 28294 -15892 28341 -15828
rect 28405 -15892 28421 -15828
rect 28294 -15908 28421 -15892
rect 21975 -15988 22102 -15972
rect 21975 -16052 22022 -15988
rect 22086 -16052 22102 -15988
rect 21975 -16068 22102 -16052
rect 21975 -16132 22022 -16068
rect 22086 -16132 22102 -16068
rect 21975 -16148 22102 -16132
rect 21975 -16212 22022 -16148
rect 22086 -16212 22102 -16148
rect 21975 -16228 22102 -16212
rect 21975 -16292 22022 -16228
rect 22086 -16292 22102 -16228
rect 21975 -16308 22102 -16292
rect 21975 -16372 22022 -16308
rect 22086 -16372 22102 -16308
rect 21975 -16388 22102 -16372
rect 21975 -16452 22022 -16388
rect 22086 -16452 22102 -16388
rect 21975 -16468 22102 -16452
rect 21975 -16532 22022 -16468
rect 22086 -16532 22102 -16468
rect 21975 -16548 22102 -16532
rect 21975 -16612 22022 -16548
rect 22086 -16612 22102 -16548
rect 21975 -16628 22102 -16612
rect 21975 -16692 22022 -16628
rect 22086 -16692 22102 -16628
rect 21975 -16708 22102 -16692
rect 21975 -16772 22022 -16708
rect 22086 -16772 22102 -16708
rect 21975 -16788 22102 -16772
rect 21975 -16852 22022 -16788
rect 22086 -16852 22102 -16788
rect 21975 -16868 22102 -16852
rect 21975 -16932 22022 -16868
rect 22086 -16932 22102 -16868
rect 21975 -16948 22102 -16932
rect 21975 -17012 22022 -16948
rect 22086 -17012 22102 -16948
rect 21975 -17028 22102 -17012
rect 21975 -17092 22022 -17028
rect 22086 -17092 22102 -17028
rect 21975 -17108 22102 -17092
rect 21975 -17172 22022 -17108
rect 22086 -17172 22102 -17108
rect 21975 -17188 22102 -17172
rect 21975 -17252 22022 -17188
rect 22086 -17252 22102 -17188
rect 21975 -17268 22102 -17252
rect 21975 -17332 22022 -17268
rect 22086 -17332 22102 -17268
rect 21975 -17348 22102 -17332
rect 21975 -17412 22022 -17348
rect 22086 -17412 22102 -17348
rect 21975 -17428 22102 -17412
rect 21975 -17492 22022 -17428
rect 22086 -17492 22102 -17428
rect 21975 -17508 22102 -17492
rect 21975 -17572 22022 -17508
rect 22086 -17572 22102 -17508
rect 21975 -17588 22102 -17572
rect 21975 -17652 22022 -17588
rect 22086 -17652 22102 -17588
rect 21975 -17668 22102 -17652
rect 21975 -17732 22022 -17668
rect 22086 -17732 22102 -17668
rect 21975 -17748 22102 -17732
rect 21975 -17812 22022 -17748
rect 22086 -17812 22102 -17748
rect 21975 -17828 22102 -17812
rect 21975 -17892 22022 -17828
rect 22086 -17892 22102 -17828
rect 21975 -17908 22102 -17892
rect 21975 -17972 22022 -17908
rect 22086 -17972 22102 -17908
rect 21975 -17988 22102 -17972
rect 21975 -18052 22022 -17988
rect 22086 -18052 22102 -17988
rect 21975 -18068 22102 -18052
rect 21975 -18132 22022 -18068
rect 22086 -18132 22102 -18068
rect 21975 -18148 22102 -18132
rect 21975 -18212 22022 -18148
rect 22086 -18212 22102 -18148
rect 21975 -18228 22102 -18212
rect 21975 -18292 22022 -18228
rect 22086 -18292 22102 -18228
rect 21975 -18308 22102 -18292
rect 21975 -18372 22022 -18308
rect 22086 -18372 22102 -18308
rect 21975 -18388 22102 -18372
rect 21975 -18452 22022 -18388
rect 22086 -18452 22102 -18388
rect 21975 -18468 22102 -18452
rect 21975 -18532 22022 -18468
rect 22086 -18532 22102 -18468
rect 21975 -18548 22102 -18532
rect 21975 -18612 22022 -18548
rect 22086 -18612 22102 -18548
rect 21975 -18628 22102 -18612
rect 21975 -18692 22022 -18628
rect 22086 -18692 22102 -18628
rect 21975 -18708 22102 -18692
rect 21975 -18772 22022 -18708
rect 22086 -18772 22102 -18708
rect 21975 -18788 22102 -18772
rect 21975 -18852 22022 -18788
rect 22086 -18852 22102 -18788
rect 21975 -18868 22102 -18852
rect 21975 -18932 22022 -18868
rect 22086 -18932 22102 -18868
rect 21975 -18948 22102 -18932
rect 21975 -19012 22022 -18948
rect 22086 -19012 22102 -18948
rect 21975 -19028 22102 -19012
rect 21975 -19092 22022 -19028
rect 22086 -19092 22102 -19028
rect 21975 -19108 22102 -19092
rect 21975 -19172 22022 -19108
rect 22086 -19172 22102 -19108
rect 21975 -19188 22102 -19172
rect 21975 -19252 22022 -19188
rect 22086 -19252 22102 -19188
rect 21975 -19268 22102 -19252
rect 21975 -19332 22022 -19268
rect 22086 -19332 22102 -19268
rect 21975 -19348 22102 -19332
rect 21975 -19412 22022 -19348
rect 22086 -19412 22102 -19348
rect 21975 -19428 22102 -19412
rect 21975 -19492 22022 -19428
rect 22086 -19492 22102 -19428
rect 21975 -19508 22102 -19492
rect 21975 -19572 22022 -19508
rect 22086 -19572 22102 -19508
rect 21975 -19588 22102 -19572
rect 21975 -19652 22022 -19588
rect 22086 -19652 22102 -19588
rect 21975 -19668 22102 -19652
rect 21975 -19732 22022 -19668
rect 22086 -19732 22102 -19668
rect 21975 -19748 22102 -19732
rect 21975 -19812 22022 -19748
rect 22086 -19812 22102 -19748
rect 21975 -19828 22102 -19812
rect 21975 -19892 22022 -19828
rect 22086 -19892 22102 -19828
rect 21975 -19908 22102 -19892
rect 21975 -19972 22022 -19908
rect 22086 -19972 22102 -19908
rect 21975 -19988 22102 -19972
rect 21975 -20052 22022 -19988
rect 22086 -20052 22102 -19988
rect 21975 -20068 22102 -20052
rect 21975 -20132 22022 -20068
rect 22086 -20132 22102 -20068
rect 21975 -20148 22102 -20132
rect 21975 -20212 22022 -20148
rect 22086 -20212 22102 -20148
rect 21975 -20228 22102 -20212
rect 21975 -20292 22022 -20228
rect 22086 -20292 22102 -20228
rect 21975 -20308 22102 -20292
rect 21975 -20372 22022 -20308
rect 22086 -20372 22102 -20308
rect 21975 -20388 22102 -20372
rect 21975 -20452 22022 -20388
rect 22086 -20452 22102 -20388
rect 21975 -20468 22102 -20452
rect 21975 -20532 22022 -20468
rect 22086 -20532 22102 -20468
rect 21975 -20548 22102 -20532
rect 21975 -20612 22022 -20548
rect 22086 -20612 22102 -20548
rect 21975 -20628 22102 -20612
rect 21975 -20692 22022 -20628
rect 22086 -20692 22102 -20628
rect 21975 -20708 22102 -20692
rect 21975 -20772 22022 -20708
rect 22086 -20772 22102 -20708
rect 21975 -20788 22102 -20772
rect 21975 -20852 22022 -20788
rect 22086 -20852 22102 -20788
rect 21975 -20868 22102 -20852
rect 21975 -20932 22022 -20868
rect 22086 -20932 22102 -20868
rect 21975 -20948 22102 -20932
rect 21975 -21012 22022 -20948
rect 22086 -21012 22102 -20948
rect 21975 -21028 22102 -21012
rect 21975 -21092 22022 -21028
rect 22086 -21092 22102 -21028
rect 21975 -21108 22102 -21092
rect 21975 -21172 22022 -21108
rect 22086 -21172 22102 -21108
rect 21975 -21188 22102 -21172
rect 21975 -21252 22022 -21188
rect 22086 -21252 22102 -21188
rect 21975 -21268 22102 -21252
rect 21975 -21332 22022 -21268
rect 22086 -21332 22102 -21268
rect 21975 -21348 22102 -21332
rect 21975 -21412 22022 -21348
rect 22086 -21412 22102 -21348
rect 21975 -21428 22102 -21412
rect 21975 -21492 22022 -21428
rect 22086 -21492 22102 -21428
rect 21975 -21508 22102 -21492
rect 21975 -21572 22022 -21508
rect 22086 -21572 22102 -21508
rect 21975 -21588 22102 -21572
rect 21975 -21652 22022 -21588
rect 22086 -21652 22102 -21588
rect 21975 -21668 22102 -21652
rect 21975 -21732 22022 -21668
rect 22086 -21732 22102 -21668
rect 21975 -21748 22102 -21732
rect 21975 -21812 22022 -21748
rect 22086 -21812 22102 -21748
rect 21975 -21828 22102 -21812
rect 15656 -21908 15783 -21892
rect 15656 -21972 15703 -21908
rect 15767 -21972 15783 -21908
rect 15656 -21988 15783 -21972
rect 15656 -22112 15760 -21988
rect 15656 -22128 15783 -22112
rect 15656 -22192 15703 -22128
rect 15767 -22192 15783 -22128
rect 15656 -22208 15783 -22192
rect 9337 -22288 9464 -22272
rect 9337 -22352 9384 -22288
rect 9448 -22352 9464 -22288
rect 9337 -22368 9464 -22352
rect 9337 -22432 9384 -22368
rect 9448 -22432 9464 -22368
rect 9337 -22448 9464 -22432
rect 9337 -22512 9384 -22448
rect 9448 -22512 9464 -22448
rect 9337 -22528 9464 -22512
rect 9337 -22592 9384 -22528
rect 9448 -22592 9464 -22528
rect 9337 -22608 9464 -22592
rect 9337 -22672 9384 -22608
rect 9448 -22672 9464 -22608
rect 9337 -22688 9464 -22672
rect 9337 -22752 9384 -22688
rect 9448 -22752 9464 -22688
rect 9337 -22768 9464 -22752
rect 9337 -22832 9384 -22768
rect 9448 -22832 9464 -22768
rect 9337 -22848 9464 -22832
rect 9337 -22912 9384 -22848
rect 9448 -22912 9464 -22848
rect 9337 -22928 9464 -22912
rect 9337 -22992 9384 -22928
rect 9448 -22992 9464 -22928
rect 9337 -23008 9464 -22992
rect 9337 -23072 9384 -23008
rect 9448 -23072 9464 -23008
rect 9337 -23088 9464 -23072
rect 9337 -23152 9384 -23088
rect 9448 -23152 9464 -23088
rect 9337 -23168 9464 -23152
rect 9337 -23232 9384 -23168
rect 9448 -23232 9464 -23168
rect 9337 -23248 9464 -23232
rect 9337 -23312 9384 -23248
rect 9448 -23312 9464 -23248
rect 9337 -23328 9464 -23312
rect 9337 -23392 9384 -23328
rect 9448 -23392 9464 -23328
rect 9337 -23408 9464 -23392
rect 9337 -23472 9384 -23408
rect 9448 -23472 9464 -23408
rect 9337 -23488 9464 -23472
rect 9337 -23552 9384 -23488
rect 9448 -23552 9464 -23488
rect 9337 -23568 9464 -23552
rect 9337 -23632 9384 -23568
rect 9448 -23632 9464 -23568
rect 9337 -23648 9464 -23632
rect 9337 -23712 9384 -23648
rect 9448 -23712 9464 -23648
rect 9337 -23728 9464 -23712
rect 9337 -23792 9384 -23728
rect 9448 -23792 9464 -23728
rect 9337 -23808 9464 -23792
rect 9337 -23872 9384 -23808
rect 9448 -23872 9464 -23808
rect 9337 -23888 9464 -23872
rect 9337 -23952 9384 -23888
rect 9448 -23952 9464 -23888
rect 9337 -23968 9464 -23952
rect 9337 -24032 9384 -23968
rect 9448 -24032 9464 -23968
rect 9337 -24048 9464 -24032
rect 9337 -24112 9384 -24048
rect 9448 -24112 9464 -24048
rect 9337 -24128 9464 -24112
rect 9337 -24192 9384 -24128
rect 9448 -24192 9464 -24128
rect 9337 -24208 9464 -24192
rect 9337 -24272 9384 -24208
rect 9448 -24272 9464 -24208
rect 9337 -24288 9464 -24272
rect 9337 -24352 9384 -24288
rect 9448 -24352 9464 -24288
rect 9337 -24368 9464 -24352
rect 9337 -24432 9384 -24368
rect 9448 -24432 9464 -24368
rect 9337 -24448 9464 -24432
rect 9337 -24512 9384 -24448
rect 9448 -24512 9464 -24448
rect 9337 -24528 9464 -24512
rect 9337 -24592 9384 -24528
rect 9448 -24592 9464 -24528
rect 9337 -24608 9464 -24592
rect 9337 -24672 9384 -24608
rect 9448 -24672 9464 -24608
rect 9337 -24688 9464 -24672
rect 9337 -24752 9384 -24688
rect 9448 -24752 9464 -24688
rect 9337 -24768 9464 -24752
rect 9337 -24832 9384 -24768
rect 9448 -24832 9464 -24768
rect 9337 -24848 9464 -24832
rect 9337 -24912 9384 -24848
rect 9448 -24912 9464 -24848
rect 9337 -24928 9464 -24912
rect 9337 -24992 9384 -24928
rect 9448 -24992 9464 -24928
rect 9337 -25008 9464 -24992
rect 9337 -25072 9384 -25008
rect 9448 -25072 9464 -25008
rect 9337 -25088 9464 -25072
rect 9337 -25152 9384 -25088
rect 9448 -25152 9464 -25088
rect 9337 -25168 9464 -25152
rect 9337 -25232 9384 -25168
rect 9448 -25232 9464 -25168
rect 9337 -25248 9464 -25232
rect 9337 -25312 9384 -25248
rect 9448 -25312 9464 -25248
rect 9337 -25328 9464 -25312
rect 9337 -25392 9384 -25328
rect 9448 -25392 9464 -25328
rect 9337 -25408 9464 -25392
rect 9337 -25472 9384 -25408
rect 9448 -25472 9464 -25408
rect 9337 -25488 9464 -25472
rect 9337 -25552 9384 -25488
rect 9448 -25552 9464 -25488
rect 9337 -25568 9464 -25552
rect 9337 -25632 9384 -25568
rect 9448 -25632 9464 -25568
rect 9337 -25648 9464 -25632
rect 9337 -25712 9384 -25648
rect 9448 -25712 9464 -25648
rect 9337 -25728 9464 -25712
rect 9337 -25792 9384 -25728
rect 9448 -25792 9464 -25728
rect 9337 -25808 9464 -25792
rect 9337 -25872 9384 -25808
rect 9448 -25872 9464 -25808
rect 9337 -25888 9464 -25872
rect 9337 -25952 9384 -25888
rect 9448 -25952 9464 -25888
rect 9337 -25968 9464 -25952
rect 9337 -26032 9384 -25968
rect 9448 -26032 9464 -25968
rect 9337 -26048 9464 -26032
rect 9337 -26112 9384 -26048
rect 9448 -26112 9464 -26048
rect 9337 -26128 9464 -26112
rect 9337 -26192 9384 -26128
rect 9448 -26192 9464 -26128
rect 9337 -26208 9464 -26192
rect 9337 -26272 9384 -26208
rect 9448 -26272 9464 -26208
rect 9337 -26288 9464 -26272
rect 9337 -26352 9384 -26288
rect 9448 -26352 9464 -26288
rect 9337 -26368 9464 -26352
rect 9337 -26432 9384 -26368
rect 9448 -26432 9464 -26368
rect 9337 -26448 9464 -26432
rect 9337 -26512 9384 -26448
rect 9448 -26512 9464 -26448
rect 9337 -26528 9464 -26512
rect 9337 -26592 9384 -26528
rect 9448 -26592 9464 -26528
rect 9337 -26608 9464 -26592
rect 9337 -26672 9384 -26608
rect 9448 -26672 9464 -26608
rect 9337 -26688 9464 -26672
rect 9337 -26752 9384 -26688
rect 9448 -26752 9464 -26688
rect 9337 -26768 9464 -26752
rect 9337 -26832 9384 -26768
rect 9448 -26832 9464 -26768
rect 9337 -26848 9464 -26832
rect 9337 -26912 9384 -26848
rect 9448 -26912 9464 -26848
rect 9337 -26928 9464 -26912
rect 9337 -26992 9384 -26928
rect 9448 -26992 9464 -26928
rect 9337 -27008 9464 -26992
rect 9337 -27072 9384 -27008
rect 9448 -27072 9464 -27008
rect 9337 -27088 9464 -27072
rect 9337 -27152 9384 -27088
rect 9448 -27152 9464 -27088
rect 9337 -27168 9464 -27152
rect 9337 -27232 9384 -27168
rect 9448 -27232 9464 -27168
rect 9337 -27248 9464 -27232
rect 9337 -27312 9384 -27248
rect 9448 -27312 9464 -27248
rect 9337 -27328 9464 -27312
rect 9337 -27392 9384 -27328
rect 9448 -27392 9464 -27328
rect 9337 -27408 9464 -27392
rect 9337 -27472 9384 -27408
rect 9448 -27472 9464 -27408
rect 9337 -27488 9464 -27472
rect 9337 -27552 9384 -27488
rect 9448 -27552 9464 -27488
rect 9337 -27568 9464 -27552
rect 9337 -27632 9384 -27568
rect 9448 -27632 9464 -27568
rect 9337 -27648 9464 -27632
rect 9337 -27712 9384 -27648
rect 9448 -27712 9464 -27648
rect 9337 -27728 9464 -27712
rect 9337 -27792 9384 -27728
rect 9448 -27792 9464 -27728
rect 9337 -27808 9464 -27792
rect 9337 -27872 9384 -27808
rect 9448 -27872 9464 -27808
rect 9337 -27888 9464 -27872
rect 9337 -27952 9384 -27888
rect 9448 -27952 9464 -27888
rect 9337 -27968 9464 -27952
rect 9337 -28032 9384 -27968
rect 9448 -28032 9464 -27968
rect 9337 -28048 9464 -28032
rect 9337 -28112 9384 -28048
rect 9448 -28112 9464 -28048
rect 9337 -28128 9464 -28112
rect 3018 -28208 3145 -28192
rect 3018 -28272 3065 -28208
rect 3129 -28272 3145 -28208
rect 3018 -28288 3145 -28272
rect 3018 -28412 3122 -28288
rect 3018 -28428 3145 -28412
rect 3018 -28492 3065 -28428
rect 3129 -28492 3145 -28428
rect 3018 -28508 3145 -28492
rect -3301 -28588 -3174 -28572
rect -3301 -28652 -3254 -28588
rect -3190 -28652 -3174 -28588
rect -3301 -28668 -3174 -28652
rect -3301 -28732 -3254 -28668
rect -3190 -28732 -3174 -28668
rect -3301 -28748 -3174 -28732
rect -3301 -28812 -3254 -28748
rect -3190 -28812 -3174 -28748
rect -3301 -28828 -3174 -28812
rect -3301 -28892 -3254 -28828
rect -3190 -28892 -3174 -28828
rect -3301 -28908 -3174 -28892
rect -3301 -28972 -3254 -28908
rect -3190 -28972 -3174 -28908
rect -3301 -28988 -3174 -28972
rect -3301 -29052 -3254 -28988
rect -3190 -29052 -3174 -28988
rect -3301 -29068 -3174 -29052
rect -3301 -29132 -3254 -29068
rect -3190 -29132 -3174 -29068
rect -3301 -29148 -3174 -29132
rect -3301 -29212 -3254 -29148
rect -3190 -29212 -3174 -29148
rect -3301 -29228 -3174 -29212
rect -3301 -29292 -3254 -29228
rect -3190 -29292 -3174 -29228
rect -3301 -29308 -3174 -29292
rect -3301 -29372 -3254 -29308
rect -3190 -29372 -3174 -29308
rect -3301 -29388 -3174 -29372
rect -3301 -29452 -3254 -29388
rect -3190 -29452 -3174 -29388
rect -3301 -29468 -3174 -29452
rect -3301 -29532 -3254 -29468
rect -3190 -29532 -3174 -29468
rect -3301 -29548 -3174 -29532
rect -3301 -29612 -3254 -29548
rect -3190 -29612 -3174 -29548
rect -3301 -29628 -3174 -29612
rect -3301 -29692 -3254 -29628
rect -3190 -29692 -3174 -29628
rect -3301 -29708 -3174 -29692
rect -3301 -29772 -3254 -29708
rect -3190 -29772 -3174 -29708
rect -3301 -29788 -3174 -29772
rect -3301 -29852 -3254 -29788
rect -3190 -29852 -3174 -29788
rect -3301 -29868 -3174 -29852
rect -3301 -29932 -3254 -29868
rect -3190 -29932 -3174 -29868
rect -3301 -29948 -3174 -29932
rect -3301 -30012 -3254 -29948
rect -3190 -30012 -3174 -29948
rect -3301 -30028 -3174 -30012
rect -3301 -30092 -3254 -30028
rect -3190 -30092 -3174 -30028
rect -3301 -30108 -3174 -30092
rect -3301 -30172 -3254 -30108
rect -3190 -30172 -3174 -30108
rect -3301 -30188 -3174 -30172
rect -3301 -30252 -3254 -30188
rect -3190 -30252 -3174 -30188
rect -3301 -30268 -3174 -30252
rect -3301 -30332 -3254 -30268
rect -3190 -30332 -3174 -30268
rect -3301 -30348 -3174 -30332
rect -3301 -30412 -3254 -30348
rect -3190 -30412 -3174 -30348
rect -3301 -30428 -3174 -30412
rect -3301 -30492 -3254 -30428
rect -3190 -30492 -3174 -30428
rect -3301 -30508 -3174 -30492
rect -3301 -30572 -3254 -30508
rect -3190 -30572 -3174 -30508
rect -3301 -30588 -3174 -30572
rect -3301 -30652 -3254 -30588
rect -3190 -30652 -3174 -30588
rect -3301 -30668 -3174 -30652
rect -3301 -30732 -3254 -30668
rect -3190 -30732 -3174 -30668
rect -3301 -30748 -3174 -30732
rect -3301 -30812 -3254 -30748
rect -3190 -30812 -3174 -30748
rect -3301 -30828 -3174 -30812
rect -3301 -30892 -3254 -30828
rect -3190 -30892 -3174 -30828
rect -3301 -30908 -3174 -30892
rect -3301 -30972 -3254 -30908
rect -3190 -30972 -3174 -30908
rect -3301 -30988 -3174 -30972
rect -3301 -31052 -3254 -30988
rect -3190 -31052 -3174 -30988
rect -3301 -31068 -3174 -31052
rect -3301 -31132 -3254 -31068
rect -3190 -31132 -3174 -31068
rect -3301 -31148 -3174 -31132
rect -3301 -31212 -3254 -31148
rect -3190 -31212 -3174 -31148
rect -3301 -31228 -3174 -31212
rect -3301 -31292 -3254 -31228
rect -3190 -31292 -3174 -31228
rect -3301 -31308 -3174 -31292
rect -3301 -31372 -3254 -31308
rect -3190 -31372 -3174 -31308
rect -3301 -31388 -3174 -31372
rect -3301 -31452 -3254 -31388
rect -3190 -31452 -3174 -31388
rect -3301 -31468 -3174 -31452
rect -3301 -31532 -3254 -31468
rect -3190 -31532 -3174 -31468
rect -3301 -31548 -3174 -31532
rect -3301 -31612 -3254 -31548
rect -3190 -31612 -3174 -31548
rect -3301 -31628 -3174 -31612
rect -3301 -31692 -3254 -31628
rect -3190 -31692 -3174 -31628
rect -3301 -31708 -3174 -31692
rect -3301 -31772 -3254 -31708
rect -3190 -31772 -3174 -31708
rect -3301 -31788 -3174 -31772
rect -3301 -31852 -3254 -31788
rect -3190 -31852 -3174 -31788
rect -3301 -31868 -3174 -31852
rect -3301 -31932 -3254 -31868
rect -3190 -31932 -3174 -31868
rect -3301 -31948 -3174 -31932
rect -3301 -32012 -3254 -31948
rect -3190 -32012 -3174 -31948
rect -3301 -32028 -3174 -32012
rect -3301 -32092 -3254 -32028
rect -3190 -32092 -3174 -32028
rect -3301 -32108 -3174 -32092
rect -3301 -32172 -3254 -32108
rect -3190 -32172 -3174 -32108
rect -3301 -32188 -3174 -32172
rect -3301 -32252 -3254 -32188
rect -3190 -32252 -3174 -32188
rect -3301 -32268 -3174 -32252
rect -3301 -32332 -3254 -32268
rect -3190 -32332 -3174 -32268
rect -3301 -32348 -3174 -32332
rect -3301 -32412 -3254 -32348
rect -3190 -32412 -3174 -32348
rect -3301 -32428 -3174 -32412
rect -3301 -32492 -3254 -32428
rect -3190 -32492 -3174 -32428
rect -3301 -32508 -3174 -32492
rect -3301 -32572 -3254 -32508
rect -3190 -32572 -3174 -32508
rect -3301 -32588 -3174 -32572
rect -3301 -32652 -3254 -32588
rect -3190 -32652 -3174 -32588
rect -3301 -32668 -3174 -32652
rect -3301 -32732 -3254 -32668
rect -3190 -32732 -3174 -32668
rect -3301 -32748 -3174 -32732
rect -3301 -32812 -3254 -32748
rect -3190 -32812 -3174 -32748
rect -3301 -32828 -3174 -32812
rect -3301 -32892 -3254 -32828
rect -3190 -32892 -3174 -32828
rect -3301 -32908 -3174 -32892
rect -3301 -32972 -3254 -32908
rect -3190 -32972 -3174 -32908
rect -3301 -32988 -3174 -32972
rect -3301 -33052 -3254 -32988
rect -3190 -33052 -3174 -32988
rect -3301 -33068 -3174 -33052
rect -3301 -33132 -3254 -33068
rect -3190 -33132 -3174 -33068
rect -3301 -33148 -3174 -33132
rect -3301 -33212 -3254 -33148
rect -3190 -33212 -3174 -33148
rect -3301 -33228 -3174 -33212
rect -3301 -33292 -3254 -33228
rect -3190 -33292 -3174 -33228
rect -3301 -33308 -3174 -33292
rect -3301 -33372 -3254 -33308
rect -3190 -33372 -3174 -33308
rect -3301 -33388 -3174 -33372
rect -3301 -33452 -3254 -33388
rect -3190 -33452 -3174 -33388
rect -3301 -33468 -3174 -33452
rect -3301 -33532 -3254 -33468
rect -3190 -33532 -3174 -33468
rect -3301 -33548 -3174 -33532
rect -3301 -33612 -3254 -33548
rect -3190 -33612 -3174 -33548
rect -3301 -33628 -3174 -33612
rect -3301 -33692 -3254 -33628
rect -3190 -33692 -3174 -33628
rect -3301 -33708 -3174 -33692
rect -3301 -33772 -3254 -33708
rect -3190 -33772 -3174 -33708
rect -3301 -33788 -3174 -33772
rect -3301 -33852 -3254 -33788
rect -3190 -33852 -3174 -33788
rect -3301 -33868 -3174 -33852
rect -3301 -33932 -3254 -33868
rect -3190 -33932 -3174 -33868
rect -3301 -33948 -3174 -33932
rect -3301 -34012 -3254 -33948
rect -3190 -34012 -3174 -33948
rect -3301 -34028 -3174 -34012
rect -3301 -34092 -3254 -34028
rect -3190 -34092 -3174 -34028
rect -3301 -34108 -3174 -34092
rect -3301 -34172 -3254 -34108
rect -3190 -34172 -3174 -34108
rect -3301 -34188 -3174 -34172
rect -3301 -34252 -3254 -34188
rect -3190 -34252 -3174 -34188
rect -3301 -34268 -3174 -34252
rect -3301 -34332 -3254 -34268
rect -3190 -34332 -3174 -34268
rect -3301 -34348 -3174 -34332
rect -3301 -34412 -3254 -34348
rect -3190 -34412 -3174 -34348
rect -3301 -34428 -3174 -34412
rect -9620 -34508 -9493 -34492
rect -9620 -34572 -9573 -34508
rect -9509 -34572 -9493 -34508
rect -9620 -34588 -9493 -34572
rect -9620 -34712 -9516 -34588
rect -9620 -34728 -9493 -34712
rect -9620 -34792 -9573 -34728
rect -9509 -34792 -9493 -34728
rect -9620 -34808 -9493 -34792
rect -15939 -34888 -15812 -34872
rect -15939 -34952 -15892 -34888
rect -15828 -34952 -15812 -34888
rect -15939 -34968 -15812 -34952
rect -15939 -35032 -15892 -34968
rect -15828 -35032 -15812 -34968
rect -15939 -35048 -15812 -35032
rect -15939 -35112 -15892 -35048
rect -15828 -35112 -15812 -35048
rect -15939 -35128 -15812 -35112
rect -15939 -35192 -15892 -35128
rect -15828 -35192 -15812 -35128
rect -15939 -35208 -15812 -35192
rect -15939 -35272 -15892 -35208
rect -15828 -35272 -15812 -35208
rect -15939 -35288 -15812 -35272
rect -15939 -35352 -15892 -35288
rect -15828 -35352 -15812 -35288
rect -15939 -35368 -15812 -35352
rect -15939 -35432 -15892 -35368
rect -15828 -35432 -15812 -35368
rect -15939 -35448 -15812 -35432
rect -15939 -35512 -15892 -35448
rect -15828 -35512 -15812 -35448
rect -15939 -35528 -15812 -35512
rect -15939 -35592 -15892 -35528
rect -15828 -35592 -15812 -35528
rect -15939 -35608 -15812 -35592
rect -15939 -35672 -15892 -35608
rect -15828 -35672 -15812 -35608
rect -15939 -35688 -15812 -35672
rect -15939 -35752 -15892 -35688
rect -15828 -35752 -15812 -35688
rect -15939 -35768 -15812 -35752
rect -15939 -35832 -15892 -35768
rect -15828 -35832 -15812 -35768
rect -15939 -35848 -15812 -35832
rect -15939 -35912 -15892 -35848
rect -15828 -35912 -15812 -35848
rect -15939 -35928 -15812 -35912
rect -15939 -35992 -15892 -35928
rect -15828 -35992 -15812 -35928
rect -15939 -36008 -15812 -35992
rect -15939 -36072 -15892 -36008
rect -15828 -36072 -15812 -36008
rect -15939 -36088 -15812 -36072
rect -15939 -36152 -15892 -36088
rect -15828 -36152 -15812 -36088
rect -15939 -36168 -15812 -36152
rect -15939 -36232 -15892 -36168
rect -15828 -36232 -15812 -36168
rect -15939 -36248 -15812 -36232
rect -15939 -36312 -15892 -36248
rect -15828 -36312 -15812 -36248
rect -15939 -36328 -15812 -36312
rect -15939 -36392 -15892 -36328
rect -15828 -36392 -15812 -36328
rect -15939 -36408 -15812 -36392
rect -15939 -36472 -15892 -36408
rect -15828 -36472 -15812 -36408
rect -15939 -36488 -15812 -36472
rect -15939 -36552 -15892 -36488
rect -15828 -36552 -15812 -36488
rect -15939 -36568 -15812 -36552
rect -15939 -36632 -15892 -36568
rect -15828 -36632 -15812 -36568
rect -15939 -36648 -15812 -36632
rect -15939 -36712 -15892 -36648
rect -15828 -36712 -15812 -36648
rect -15939 -36728 -15812 -36712
rect -15939 -36792 -15892 -36728
rect -15828 -36792 -15812 -36728
rect -15939 -36808 -15812 -36792
rect -15939 -36872 -15892 -36808
rect -15828 -36872 -15812 -36808
rect -15939 -36888 -15812 -36872
rect -15939 -36952 -15892 -36888
rect -15828 -36952 -15812 -36888
rect -15939 -36968 -15812 -36952
rect -15939 -37032 -15892 -36968
rect -15828 -37032 -15812 -36968
rect -15939 -37048 -15812 -37032
rect -15939 -37112 -15892 -37048
rect -15828 -37112 -15812 -37048
rect -15939 -37128 -15812 -37112
rect -15939 -37192 -15892 -37128
rect -15828 -37192 -15812 -37128
rect -15939 -37208 -15812 -37192
rect -15939 -37272 -15892 -37208
rect -15828 -37272 -15812 -37208
rect -15939 -37288 -15812 -37272
rect -15939 -37352 -15892 -37288
rect -15828 -37352 -15812 -37288
rect -15939 -37368 -15812 -37352
rect -15939 -37432 -15892 -37368
rect -15828 -37432 -15812 -37368
rect -15939 -37448 -15812 -37432
rect -15939 -37512 -15892 -37448
rect -15828 -37512 -15812 -37448
rect -15939 -37528 -15812 -37512
rect -15939 -37592 -15892 -37528
rect -15828 -37592 -15812 -37528
rect -15939 -37608 -15812 -37592
rect -15939 -37672 -15892 -37608
rect -15828 -37672 -15812 -37608
rect -15939 -37688 -15812 -37672
rect -15939 -37752 -15892 -37688
rect -15828 -37752 -15812 -37688
rect -15939 -37768 -15812 -37752
rect -15939 -37832 -15892 -37768
rect -15828 -37832 -15812 -37768
rect -15939 -37848 -15812 -37832
rect -15939 -37912 -15892 -37848
rect -15828 -37912 -15812 -37848
rect -15939 -37928 -15812 -37912
rect -15939 -37992 -15892 -37928
rect -15828 -37992 -15812 -37928
rect -15939 -38008 -15812 -37992
rect -15939 -38072 -15892 -38008
rect -15828 -38072 -15812 -38008
rect -15939 -38088 -15812 -38072
rect -15939 -38152 -15892 -38088
rect -15828 -38152 -15812 -38088
rect -15939 -38168 -15812 -38152
rect -15939 -38232 -15892 -38168
rect -15828 -38232 -15812 -38168
rect -15939 -38248 -15812 -38232
rect -15939 -38312 -15892 -38248
rect -15828 -38312 -15812 -38248
rect -15939 -38328 -15812 -38312
rect -15939 -38392 -15892 -38328
rect -15828 -38392 -15812 -38328
rect -15939 -38408 -15812 -38392
rect -15939 -38472 -15892 -38408
rect -15828 -38472 -15812 -38408
rect -15939 -38488 -15812 -38472
rect -15939 -38552 -15892 -38488
rect -15828 -38552 -15812 -38488
rect -15939 -38568 -15812 -38552
rect -15939 -38632 -15892 -38568
rect -15828 -38632 -15812 -38568
rect -15939 -38648 -15812 -38632
rect -15939 -38712 -15892 -38648
rect -15828 -38712 -15812 -38648
rect -15939 -38728 -15812 -38712
rect -15939 -38792 -15892 -38728
rect -15828 -38792 -15812 -38728
rect -15939 -38808 -15812 -38792
rect -15939 -38872 -15892 -38808
rect -15828 -38872 -15812 -38808
rect -15939 -38888 -15812 -38872
rect -15939 -38952 -15892 -38888
rect -15828 -38952 -15812 -38888
rect -15939 -38968 -15812 -38952
rect -15939 -39032 -15892 -38968
rect -15828 -39032 -15812 -38968
rect -15939 -39048 -15812 -39032
rect -15939 -39112 -15892 -39048
rect -15828 -39112 -15812 -39048
rect -15939 -39128 -15812 -39112
rect -15939 -39192 -15892 -39128
rect -15828 -39192 -15812 -39128
rect -15939 -39208 -15812 -39192
rect -15939 -39272 -15892 -39208
rect -15828 -39272 -15812 -39208
rect -15939 -39288 -15812 -39272
rect -15939 -39352 -15892 -39288
rect -15828 -39352 -15812 -39288
rect -15939 -39368 -15812 -39352
rect -15939 -39432 -15892 -39368
rect -15828 -39432 -15812 -39368
rect -15939 -39448 -15812 -39432
rect -15939 -39512 -15892 -39448
rect -15828 -39512 -15812 -39448
rect -15939 -39528 -15812 -39512
rect -15939 -39592 -15892 -39528
rect -15828 -39592 -15812 -39528
rect -15939 -39608 -15812 -39592
rect -15939 -39672 -15892 -39608
rect -15828 -39672 -15812 -39608
rect -15939 -39688 -15812 -39672
rect -15939 -39752 -15892 -39688
rect -15828 -39752 -15812 -39688
rect -15939 -39768 -15812 -39752
rect -15939 -39832 -15892 -39768
rect -15828 -39832 -15812 -39768
rect -15939 -39848 -15812 -39832
rect -15939 -39912 -15892 -39848
rect -15828 -39912 -15812 -39848
rect -15939 -39928 -15812 -39912
rect -15939 -39992 -15892 -39928
rect -15828 -39992 -15812 -39928
rect -15939 -40008 -15812 -39992
rect -15939 -40072 -15892 -40008
rect -15828 -40072 -15812 -40008
rect -15939 -40088 -15812 -40072
rect -15939 -40152 -15892 -40088
rect -15828 -40152 -15812 -40088
rect -15939 -40168 -15812 -40152
rect -15939 -40232 -15892 -40168
rect -15828 -40232 -15812 -40168
rect -15939 -40248 -15812 -40232
rect -15939 -40312 -15892 -40248
rect -15828 -40312 -15812 -40248
rect -15939 -40328 -15812 -40312
rect -15939 -40392 -15892 -40328
rect -15828 -40392 -15812 -40328
rect -15939 -40408 -15812 -40392
rect -15939 -40472 -15892 -40408
rect -15828 -40472 -15812 -40408
rect -15939 -40488 -15812 -40472
rect -15939 -40552 -15892 -40488
rect -15828 -40552 -15812 -40488
rect -15939 -40568 -15812 -40552
rect -15939 -40632 -15892 -40568
rect -15828 -40632 -15812 -40568
rect -15939 -40648 -15812 -40632
rect -15939 -40712 -15892 -40648
rect -15828 -40712 -15812 -40648
rect -15939 -40728 -15812 -40712
rect -22258 -40808 -22131 -40792
rect -22258 -40872 -22211 -40808
rect -22147 -40872 -22131 -40808
rect -22258 -40888 -22131 -40872
rect -22258 -41012 -22154 -40888
rect -22258 -41028 -22131 -41012
rect -22258 -41092 -22211 -41028
rect -22147 -41092 -22131 -41028
rect -22258 -41108 -22131 -41092
rect -28577 -41188 -28450 -41172
rect -28577 -41252 -28530 -41188
rect -28466 -41252 -28450 -41188
rect -28577 -41268 -28450 -41252
rect -28577 -41332 -28530 -41268
rect -28466 -41332 -28450 -41268
rect -28577 -41348 -28450 -41332
rect -28577 -41412 -28530 -41348
rect -28466 -41412 -28450 -41348
rect -28577 -41428 -28450 -41412
rect -28577 -41492 -28530 -41428
rect -28466 -41492 -28450 -41428
rect -28577 -41508 -28450 -41492
rect -28577 -41572 -28530 -41508
rect -28466 -41572 -28450 -41508
rect -28577 -41588 -28450 -41572
rect -28577 -41652 -28530 -41588
rect -28466 -41652 -28450 -41588
rect -28577 -41668 -28450 -41652
rect -28577 -41732 -28530 -41668
rect -28466 -41732 -28450 -41668
rect -28577 -41748 -28450 -41732
rect -28577 -41812 -28530 -41748
rect -28466 -41812 -28450 -41748
rect -28577 -41828 -28450 -41812
rect -28577 -41892 -28530 -41828
rect -28466 -41892 -28450 -41828
rect -28577 -41908 -28450 -41892
rect -28577 -41972 -28530 -41908
rect -28466 -41972 -28450 -41908
rect -28577 -41988 -28450 -41972
rect -28577 -42052 -28530 -41988
rect -28466 -42052 -28450 -41988
rect -28577 -42068 -28450 -42052
rect -28577 -42132 -28530 -42068
rect -28466 -42132 -28450 -42068
rect -28577 -42148 -28450 -42132
rect -28577 -42212 -28530 -42148
rect -28466 -42212 -28450 -42148
rect -28577 -42228 -28450 -42212
rect -28577 -42292 -28530 -42228
rect -28466 -42292 -28450 -42228
rect -28577 -42308 -28450 -42292
rect -28577 -42372 -28530 -42308
rect -28466 -42372 -28450 -42308
rect -28577 -42388 -28450 -42372
rect -28577 -42452 -28530 -42388
rect -28466 -42452 -28450 -42388
rect -28577 -42468 -28450 -42452
rect -28577 -42532 -28530 -42468
rect -28466 -42532 -28450 -42468
rect -28577 -42548 -28450 -42532
rect -28577 -42612 -28530 -42548
rect -28466 -42612 -28450 -42548
rect -28577 -42628 -28450 -42612
rect -28577 -42692 -28530 -42628
rect -28466 -42692 -28450 -42628
rect -28577 -42708 -28450 -42692
rect -28577 -42772 -28530 -42708
rect -28466 -42772 -28450 -42708
rect -28577 -42788 -28450 -42772
rect -28577 -42852 -28530 -42788
rect -28466 -42852 -28450 -42788
rect -28577 -42868 -28450 -42852
rect -28577 -42932 -28530 -42868
rect -28466 -42932 -28450 -42868
rect -28577 -42948 -28450 -42932
rect -28577 -43012 -28530 -42948
rect -28466 -43012 -28450 -42948
rect -28577 -43028 -28450 -43012
rect -28577 -43092 -28530 -43028
rect -28466 -43092 -28450 -43028
rect -28577 -43108 -28450 -43092
rect -28577 -43172 -28530 -43108
rect -28466 -43172 -28450 -43108
rect -28577 -43188 -28450 -43172
rect -28577 -43252 -28530 -43188
rect -28466 -43252 -28450 -43188
rect -28577 -43268 -28450 -43252
rect -28577 -43332 -28530 -43268
rect -28466 -43332 -28450 -43268
rect -28577 -43348 -28450 -43332
rect -28577 -43412 -28530 -43348
rect -28466 -43412 -28450 -43348
rect -28577 -43428 -28450 -43412
rect -28577 -43492 -28530 -43428
rect -28466 -43492 -28450 -43428
rect -28577 -43508 -28450 -43492
rect -28577 -43572 -28530 -43508
rect -28466 -43572 -28450 -43508
rect -28577 -43588 -28450 -43572
rect -28577 -43652 -28530 -43588
rect -28466 -43652 -28450 -43588
rect -28577 -43668 -28450 -43652
rect -28577 -43732 -28530 -43668
rect -28466 -43732 -28450 -43668
rect -28577 -43748 -28450 -43732
rect -28577 -43812 -28530 -43748
rect -28466 -43812 -28450 -43748
rect -28577 -43828 -28450 -43812
rect -28577 -43892 -28530 -43828
rect -28466 -43892 -28450 -43828
rect -28577 -43908 -28450 -43892
rect -28577 -43972 -28530 -43908
rect -28466 -43972 -28450 -43908
rect -28577 -43988 -28450 -43972
rect -28577 -44052 -28530 -43988
rect -28466 -44052 -28450 -43988
rect -28577 -44068 -28450 -44052
rect -28577 -44132 -28530 -44068
rect -28466 -44132 -28450 -44068
rect -28577 -44148 -28450 -44132
rect -28577 -44212 -28530 -44148
rect -28466 -44212 -28450 -44148
rect -28577 -44228 -28450 -44212
rect -28577 -44292 -28530 -44228
rect -28466 -44292 -28450 -44228
rect -28577 -44308 -28450 -44292
rect -28577 -44372 -28530 -44308
rect -28466 -44372 -28450 -44308
rect -28577 -44388 -28450 -44372
rect -28577 -44452 -28530 -44388
rect -28466 -44452 -28450 -44388
rect -28577 -44468 -28450 -44452
rect -28577 -44532 -28530 -44468
rect -28466 -44532 -28450 -44468
rect -28577 -44548 -28450 -44532
rect -28577 -44612 -28530 -44548
rect -28466 -44612 -28450 -44548
rect -28577 -44628 -28450 -44612
rect -28577 -44692 -28530 -44628
rect -28466 -44692 -28450 -44628
rect -28577 -44708 -28450 -44692
rect -28577 -44772 -28530 -44708
rect -28466 -44772 -28450 -44708
rect -28577 -44788 -28450 -44772
rect -28577 -44852 -28530 -44788
rect -28466 -44852 -28450 -44788
rect -28577 -44868 -28450 -44852
rect -28577 -44932 -28530 -44868
rect -28466 -44932 -28450 -44868
rect -28577 -44948 -28450 -44932
rect -28577 -45012 -28530 -44948
rect -28466 -45012 -28450 -44948
rect -28577 -45028 -28450 -45012
rect -28577 -45092 -28530 -45028
rect -28466 -45092 -28450 -45028
rect -28577 -45108 -28450 -45092
rect -28577 -45172 -28530 -45108
rect -28466 -45172 -28450 -45108
rect -28577 -45188 -28450 -45172
rect -28577 -45252 -28530 -45188
rect -28466 -45252 -28450 -45188
rect -28577 -45268 -28450 -45252
rect -28577 -45332 -28530 -45268
rect -28466 -45332 -28450 -45268
rect -28577 -45348 -28450 -45332
rect -28577 -45412 -28530 -45348
rect -28466 -45412 -28450 -45348
rect -28577 -45428 -28450 -45412
rect -28577 -45492 -28530 -45428
rect -28466 -45492 -28450 -45428
rect -28577 -45508 -28450 -45492
rect -28577 -45572 -28530 -45508
rect -28466 -45572 -28450 -45508
rect -28577 -45588 -28450 -45572
rect -28577 -45652 -28530 -45588
rect -28466 -45652 -28450 -45588
rect -28577 -45668 -28450 -45652
rect -28577 -45732 -28530 -45668
rect -28466 -45732 -28450 -45668
rect -28577 -45748 -28450 -45732
rect -28577 -45812 -28530 -45748
rect -28466 -45812 -28450 -45748
rect -28577 -45828 -28450 -45812
rect -28577 -45892 -28530 -45828
rect -28466 -45892 -28450 -45828
rect -28577 -45908 -28450 -45892
rect -28577 -45972 -28530 -45908
rect -28466 -45972 -28450 -45908
rect -28577 -45988 -28450 -45972
rect -28577 -46052 -28530 -45988
rect -28466 -46052 -28450 -45988
rect -28577 -46068 -28450 -46052
rect -28577 -46132 -28530 -46068
rect -28466 -46132 -28450 -46068
rect -28577 -46148 -28450 -46132
rect -28577 -46212 -28530 -46148
rect -28466 -46212 -28450 -46148
rect -28577 -46228 -28450 -46212
rect -28577 -46292 -28530 -46228
rect -28466 -46292 -28450 -46228
rect -28577 -46308 -28450 -46292
rect -28577 -46372 -28530 -46308
rect -28466 -46372 -28450 -46308
rect -28577 -46388 -28450 -46372
rect -28577 -46452 -28530 -46388
rect -28466 -46452 -28450 -46388
rect -28577 -46468 -28450 -46452
rect -28577 -46532 -28530 -46468
rect -28466 -46532 -28450 -46468
rect -28577 -46548 -28450 -46532
rect -28577 -46612 -28530 -46548
rect -28466 -46612 -28450 -46548
rect -28577 -46628 -28450 -46612
rect -28577 -46692 -28530 -46628
rect -28466 -46692 -28450 -46628
rect -28577 -46708 -28450 -46692
rect -28577 -46772 -28530 -46708
rect -28466 -46772 -28450 -46708
rect -28577 -46788 -28450 -46772
rect -28577 -46852 -28530 -46788
rect -28466 -46852 -28450 -46788
rect -28577 -46868 -28450 -46852
rect -28577 -46932 -28530 -46868
rect -28466 -46932 -28450 -46868
rect -28577 -46948 -28450 -46932
rect -28577 -47012 -28530 -46948
rect -28466 -47012 -28450 -46948
rect -28577 -47028 -28450 -47012
rect -34896 -47108 -34769 -47092
rect -34896 -47172 -34849 -47108
rect -34785 -47172 -34769 -47108
rect -34896 -47188 -34769 -47172
rect -34896 -47250 -34792 -47188
rect -31697 -47250 -31593 -47061
rect -28577 -47092 -28530 -47028
rect -28466 -47092 -28450 -47028
rect -28287 -41148 -22365 -41139
rect -28287 -47052 -28278 -41148
rect -22374 -47052 -22365 -41148
rect -28287 -47061 -22365 -47052
rect -22258 -41172 -22211 -41108
rect -22147 -41172 -22131 -41108
rect -19059 -41139 -18955 -40761
rect -15939 -40792 -15892 -40728
rect -15828 -40792 -15812 -40728
rect -15649 -34848 -9727 -34839
rect -15649 -40752 -15640 -34848
rect -9736 -40752 -9727 -34848
rect -15649 -40761 -9727 -40752
rect -9620 -34872 -9573 -34808
rect -9509 -34872 -9493 -34808
rect -6421 -34839 -6317 -34461
rect -3301 -34492 -3254 -34428
rect -3190 -34492 -3174 -34428
rect -3011 -28548 2911 -28539
rect -3011 -34452 -3002 -28548
rect 2902 -34452 2911 -28548
rect -3011 -34461 2911 -34452
rect 3018 -28572 3065 -28508
rect 3129 -28572 3145 -28508
rect 6217 -28539 6321 -28161
rect 9337 -28192 9384 -28128
rect 9448 -28192 9464 -28128
rect 9627 -22248 15549 -22239
rect 9627 -28152 9636 -22248
rect 15540 -28152 15549 -22248
rect 9627 -28161 15549 -28152
rect 15656 -22272 15703 -22208
rect 15767 -22272 15783 -22208
rect 18855 -22239 18959 -21861
rect 21975 -21892 22022 -21828
rect 22086 -21892 22102 -21828
rect 22265 -15948 28187 -15939
rect 22265 -21852 22274 -15948
rect 28178 -21852 28187 -15948
rect 22265 -21861 28187 -21852
rect 28294 -15972 28341 -15908
rect 28405 -15972 28421 -15908
rect 31493 -15939 31597 -15561
rect 34613 -15592 34660 -15528
rect 34724 -15592 34740 -15528
rect 34903 -9648 40825 -9639
rect 34903 -15552 34912 -9648
rect 40816 -15552 40825 -9648
rect 34903 -15561 40825 -15552
rect 40932 -9672 40979 -9608
rect 41043 -9672 41059 -9608
rect 44131 -9639 44235 -9261
rect 47251 -9292 47298 -9228
rect 47362 -9292 47378 -9228
rect 47251 -9308 47378 -9292
rect 47251 -9372 47298 -9308
rect 47362 -9372 47378 -9308
rect 47251 -9388 47378 -9372
rect 47251 -9512 47355 -9388
rect 47251 -9528 47378 -9512
rect 47251 -9592 47298 -9528
rect 47362 -9592 47378 -9528
rect 47251 -9608 47378 -9592
rect 40932 -9688 41059 -9672
rect 40932 -9752 40979 -9688
rect 41043 -9752 41059 -9688
rect 40932 -9768 41059 -9752
rect 40932 -9832 40979 -9768
rect 41043 -9832 41059 -9768
rect 40932 -9848 41059 -9832
rect 40932 -9912 40979 -9848
rect 41043 -9912 41059 -9848
rect 40932 -9928 41059 -9912
rect 40932 -9992 40979 -9928
rect 41043 -9992 41059 -9928
rect 40932 -10008 41059 -9992
rect 40932 -10072 40979 -10008
rect 41043 -10072 41059 -10008
rect 40932 -10088 41059 -10072
rect 40932 -10152 40979 -10088
rect 41043 -10152 41059 -10088
rect 40932 -10168 41059 -10152
rect 40932 -10232 40979 -10168
rect 41043 -10232 41059 -10168
rect 40932 -10248 41059 -10232
rect 40932 -10312 40979 -10248
rect 41043 -10312 41059 -10248
rect 40932 -10328 41059 -10312
rect 40932 -10392 40979 -10328
rect 41043 -10392 41059 -10328
rect 40932 -10408 41059 -10392
rect 40932 -10472 40979 -10408
rect 41043 -10472 41059 -10408
rect 40932 -10488 41059 -10472
rect 40932 -10552 40979 -10488
rect 41043 -10552 41059 -10488
rect 40932 -10568 41059 -10552
rect 40932 -10632 40979 -10568
rect 41043 -10632 41059 -10568
rect 40932 -10648 41059 -10632
rect 40932 -10712 40979 -10648
rect 41043 -10712 41059 -10648
rect 40932 -10728 41059 -10712
rect 40932 -10792 40979 -10728
rect 41043 -10792 41059 -10728
rect 40932 -10808 41059 -10792
rect 40932 -10872 40979 -10808
rect 41043 -10872 41059 -10808
rect 40932 -10888 41059 -10872
rect 40932 -10952 40979 -10888
rect 41043 -10952 41059 -10888
rect 40932 -10968 41059 -10952
rect 40932 -11032 40979 -10968
rect 41043 -11032 41059 -10968
rect 40932 -11048 41059 -11032
rect 40932 -11112 40979 -11048
rect 41043 -11112 41059 -11048
rect 40932 -11128 41059 -11112
rect 40932 -11192 40979 -11128
rect 41043 -11192 41059 -11128
rect 40932 -11208 41059 -11192
rect 40932 -11272 40979 -11208
rect 41043 -11272 41059 -11208
rect 40932 -11288 41059 -11272
rect 40932 -11352 40979 -11288
rect 41043 -11352 41059 -11288
rect 40932 -11368 41059 -11352
rect 40932 -11432 40979 -11368
rect 41043 -11432 41059 -11368
rect 40932 -11448 41059 -11432
rect 40932 -11512 40979 -11448
rect 41043 -11512 41059 -11448
rect 40932 -11528 41059 -11512
rect 40932 -11592 40979 -11528
rect 41043 -11592 41059 -11528
rect 40932 -11608 41059 -11592
rect 40932 -11672 40979 -11608
rect 41043 -11672 41059 -11608
rect 40932 -11688 41059 -11672
rect 40932 -11752 40979 -11688
rect 41043 -11752 41059 -11688
rect 40932 -11768 41059 -11752
rect 40932 -11832 40979 -11768
rect 41043 -11832 41059 -11768
rect 40932 -11848 41059 -11832
rect 40932 -11912 40979 -11848
rect 41043 -11912 41059 -11848
rect 40932 -11928 41059 -11912
rect 40932 -11992 40979 -11928
rect 41043 -11992 41059 -11928
rect 40932 -12008 41059 -11992
rect 40932 -12072 40979 -12008
rect 41043 -12072 41059 -12008
rect 40932 -12088 41059 -12072
rect 40932 -12152 40979 -12088
rect 41043 -12152 41059 -12088
rect 40932 -12168 41059 -12152
rect 40932 -12232 40979 -12168
rect 41043 -12232 41059 -12168
rect 40932 -12248 41059 -12232
rect 40932 -12312 40979 -12248
rect 41043 -12312 41059 -12248
rect 40932 -12328 41059 -12312
rect 40932 -12392 40979 -12328
rect 41043 -12392 41059 -12328
rect 40932 -12408 41059 -12392
rect 40932 -12472 40979 -12408
rect 41043 -12472 41059 -12408
rect 40932 -12488 41059 -12472
rect 40932 -12552 40979 -12488
rect 41043 -12552 41059 -12488
rect 40932 -12568 41059 -12552
rect 40932 -12632 40979 -12568
rect 41043 -12632 41059 -12568
rect 40932 -12648 41059 -12632
rect 40932 -12712 40979 -12648
rect 41043 -12712 41059 -12648
rect 40932 -12728 41059 -12712
rect 40932 -12792 40979 -12728
rect 41043 -12792 41059 -12728
rect 40932 -12808 41059 -12792
rect 40932 -12872 40979 -12808
rect 41043 -12872 41059 -12808
rect 40932 -12888 41059 -12872
rect 40932 -12952 40979 -12888
rect 41043 -12952 41059 -12888
rect 40932 -12968 41059 -12952
rect 40932 -13032 40979 -12968
rect 41043 -13032 41059 -12968
rect 40932 -13048 41059 -13032
rect 40932 -13112 40979 -13048
rect 41043 -13112 41059 -13048
rect 40932 -13128 41059 -13112
rect 40932 -13192 40979 -13128
rect 41043 -13192 41059 -13128
rect 40932 -13208 41059 -13192
rect 40932 -13272 40979 -13208
rect 41043 -13272 41059 -13208
rect 40932 -13288 41059 -13272
rect 40932 -13352 40979 -13288
rect 41043 -13352 41059 -13288
rect 40932 -13368 41059 -13352
rect 40932 -13432 40979 -13368
rect 41043 -13432 41059 -13368
rect 40932 -13448 41059 -13432
rect 40932 -13512 40979 -13448
rect 41043 -13512 41059 -13448
rect 40932 -13528 41059 -13512
rect 40932 -13592 40979 -13528
rect 41043 -13592 41059 -13528
rect 40932 -13608 41059 -13592
rect 40932 -13672 40979 -13608
rect 41043 -13672 41059 -13608
rect 40932 -13688 41059 -13672
rect 40932 -13752 40979 -13688
rect 41043 -13752 41059 -13688
rect 40932 -13768 41059 -13752
rect 40932 -13832 40979 -13768
rect 41043 -13832 41059 -13768
rect 40932 -13848 41059 -13832
rect 40932 -13912 40979 -13848
rect 41043 -13912 41059 -13848
rect 40932 -13928 41059 -13912
rect 40932 -13992 40979 -13928
rect 41043 -13992 41059 -13928
rect 40932 -14008 41059 -13992
rect 40932 -14072 40979 -14008
rect 41043 -14072 41059 -14008
rect 40932 -14088 41059 -14072
rect 40932 -14152 40979 -14088
rect 41043 -14152 41059 -14088
rect 40932 -14168 41059 -14152
rect 40932 -14232 40979 -14168
rect 41043 -14232 41059 -14168
rect 40932 -14248 41059 -14232
rect 40932 -14312 40979 -14248
rect 41043 -14312 41059 -14248
rect 40932 -14328 41059 -14312
rect 40932 -14392 40979 -14328
rect 41043 -14392 41059 -14328
rect 40932 -14408 41059 -14392
rect 40932 -14472 40979 -14408
rect 41043 -14472 41059 -14408
rect 40932 -14488 41059 -14472
rect 40932 -14552 40979 -14488
rect 41043 -14552 41059 -14488
rect 40932 -14568 41059 -14552
rect 40932 -14632 40979 -14568
rect 41043 -14632 41059 -14568
rect 40932 -14648 41059 -14632
rect 40932 -14712 40979 -14648
rect 41043 -14712 41059 -14648
rect 40932 -14728 41059 -14712
rect 40932 -14792 40979 -14728
rect 41043 -14792 41059 -14728
rect 40932 -14808 41059 -14792
rect 40932 -14872 40979 -14808
rect 41043 -14872 41059 -14808
rect 40932 -14888 41059 -14872
rect 40932 -14952 40979 -14888
rect 41043 -14952 41059 -14888
rect 40932 -14968 41059 -14952
rect 40932 -15032 40979 -14968
rect 41043 -15032 41059 -14968
rect 40932 -15048 41059 -15032
rect 40932 -15112 40979 -15048
rect 41043 -15112 41059 -15048
rect 40932 -15128 41059 -15112
rect 40932 -15192 40979 -15128
rect 41043 -15192 41059 -15128
rect 40932 -15208 41059 -15192
rect 40932 -15272 40979 -15208
rect 41043 -15272 41059 -15208
rect 40932 -15288 41059 -15272
rect 40932 -15352 40979 -15288
rect 41043 -15352 41059 -15288
rect 40932 -15368 41059 -15352
rect 40932 -15432 40979 -15368
rect 41043 -15432 41059 -15368
rect 40932 -15448 41059 -15432
rect 40932 -15512 40979 -15448
rect 41043 -15512 41059 -15448
rect 40932 -15528 41059 -15512
rect 34613 -15608 34740 -15592
rect 34613 -15672 34660 -15608
rect 34724 -15672 34740 -15608
rect 34613 -15688 34740 -15672
rect 34613 -15812 34717 -15688
rect 34613 -15828 34740 -15812
rect 34613 -15892 34660 -15828
rect 34724 -15892 34740 -15828
rect 34613 -15908 34740 -15892
rect 28294 -15988 28421 -15972
rect 28294 -16052 28341 -15988
rect 28405 -16052 28421 -15988
rect 28294 -16068 28421 -16052
rect 28294 -16132 28341 -16068
rect 28405 -16132 28421 -16068
rect 28294 -16148 28421 -16132
rect 28294 -16212 28341 -16148
rect 28405 -16212 28421 -16148
rect 28294 -16228 28421 -16212
rect 28294 -16292 28341 -16228
rect 28405 -16292 28421 -16228
rect 28294 -16308 28421 -16292
rect 28294 -16372 28341 -16308
rect 28405 -16372 28421 -16308
rect 28294 -16388 28421 -16372
rect 28294 -16452 28341 -16388
rect 28405 -16452 28421 -16388
rect 28294 -16468 28421 -16452
rect 28294 -16532 28341 -16468
rect 28405 -16532 28421 -16468
rect 28294 -16548 28421 -16532
rect 28294 -16612 28341 -16548
rect 28405 -16612 28421 -16548
rect 28294 -16628 28421 -16612
rect 28294 -16692 28341 -16628
rect 28405 -16692 28421 -16628
rect 28294 -16708 28421 -16692
rect 28294 -16772 28341 -16708
rect 28405 -16772 28421 -16708
rect 28294 -16788 28421 -16772
rect 28294 -16852 28341 -16788
rect 28405 -16852 28421 -16788
rect 28294 -16868 28421 -16852
rect 28294 -16932 28341 -16868
rect 28405 -16932 28421 -16868
rect 28294 -16948 28421 -16932
rect 28294 -17012 28341 -16948
rect 28405 -17012 28421 -16948
rect 28294 -17028 28421 -17012
rect 28294 -17092 28341 -17028
rect 28405 -17092 28421 -17028
rect 28294 -17108 28421 -17092
rect 28294 -17172 28341 -17108
rect 28405 -17172 28421 -17108
rect 28294 -17188 28421 -17172
rect 28294 -17252 28341 -17188
rect 28405 -17252 28421 -17188
rect 28294 -17268 28421 -17252
rect 28294 -17332 28341 -17268
rect 28405 -17332 28421 -17268
rect 28294 -17348 28421 -17332
rect 28294 -17412 28341 -17348
rect 28405 -17412 28421 -17348
rect 28294 -17428 28421 -17412
rect 28294 -17492 28341 -17428
rect 28405 -17492 28421 -17428
rect 28294 -17508 28421 -17492
rect 28294 -17572 28341 -17508
rect 28405 -17572 28421 -17508
rect 28294 -17588 28421 -17572
rect 28294 -17652 28341 -17588
rect 28405 -17652 28421 -17588
rect 28294 -17668 28421 -17652
rect 28294 -17732 28341 -17668
rect 28405 -17732 28421 -17668
rect 28294 -17748 28421 -17732
rect 28294 -17812 28341 -17748
rect 28405 -17812 28421 -17748
rect 28294 -17828 28421 -17812
rect 28294 -17892 28341 -17828
rect 28405 -17892 28421 -17828
rect 28294 -17908 28421 -17892
rect 28294 -17972 28341 -17908
rect 28405 -17972 28421 -17908
rect 28294 -17988 28421 -17972
rect 28294 -18052 28341 -17988
rect 28405 -18052 28421 -17988
rect 28294 -18068 28421 -18052
rect 28294 -18132 28341 -18068
rect 28405 -18132 28421 -18068
rect 28294 -18148 28421 -18132
rect 28294 -18212 28341 -18148
rect 28405 -18212 28421 -18148
rect 28294 -18228 28421 -18212
rect 28294 -18292 28341 -18228
rect 28405 -18292 28421 -18228
rect 28294 -18308 28421 -18292
rect 28294 -18372 28341 -18308
rect 28405 -18372 28421 -18308
rect 28294 -18388 28421 -18372
rect 28294 -18452 28341 -18388
rect 28405 -18452 28421 -18388
rect 28294 -18468 28421 -18452
rect 28294 -18532 28341 -18468
rect 28405 -18532 28421 -18468
rect 28294 -18548 28421 -18532
rect 28294 -18612 28341 -18548
rect 28405 -18612 28421 -18548
rect 28294 -18628 28421 -18612
rect 28294 -18692 28341 -18628
rect 28405 -18692 28421 -18628
rect 28294 -18708 28421 -18692
rect 28294 -18772 28341 -18708
rect 28405 -18772 28421 -18708
rect 28294 -18788 28421 -18772
rect 28294 -18852 28341 -18788
rect 28405 -18852 28421 -18788
rect 28294 -18868 28421 -18852
rect 28294 -18932 28341 -18868
rect 28405 -18932 28421 -18868
rect 28294 -18948 28421 -18932
rect 28294 -19012 28341 -18948
rect 28405 -19012 28421 -18948
rect 28294 -19028 28421 -19012
rect 28294 -19092 28341 -19028
rect 28405 -19092 28421 -19028
rect 28294 -19108 28421 -19092
rect 28294 -19172 28341 -19108
rect 28405 -19172 28421 -19108
rect 28294 -19188 28421 -19172
rect 28294 -19252 28341 -19188
rect 28405 -19252 28421 -19188
rect 28294 -19268 28421 -19252
rect 28294 -19332 28341 -19268
rect 28405 -19332 28421 -19268
rect 28294 -19348 28421 -19332
rect 28294 -19412 28341 -19348
rect 28405 -19412 28421 -19348
rect 28294 -19428 28421 -19412
rect 28294 -19492 28341 -19428
rect 28405 -19492 28421 -19428
rect 28294 -19508 28421 -19492
rect 28294 -19572 28341 -19508
rect 28405 -19572 28421 -19508
rect 28294 -19588 28421 -19572
rect 28294 -19652 28341 -19588
rect 28405 -19652 28421 -19588
rect 28294 -19668 28421 -19652
rect 28294 -19732 28341 -19668
rect 28405 -19732 28421 -19668
rect 28294 -19748 28421 -19732
rect 28294 -19812 28341 -19748
rect 28405 -19812 28421 -19748
rect 28294 -19828 28421 -19812
rect 28294 -19892 28341 -19828
rect 28405 -19892 28421 -19828
rect 28294 -19908 28421 -19892
rect 28294 -19972 28341 -19908
rect 28405 -19972 28421 -19908
rect 28294 -19988 28421 -19972
rect 28294 -20052 28341 -19988
rect 28405 -20052 28421 -19988
rect 28294 -20068 28421 -20052
rect 28294 -20132 28341 -20068
rect 28405 -20132 28421 -20068
rect 28294 -20148 28421 -20132
rect 28294 -20212 28341 -20148
rect 28405 -20212 28421 -20148
rect 28294 -20228 28421 -20212
rect 28294 -20292 28341 -20228
rect 28405 -20292 28421 -20228
rect 28294 -20308 28421 -20292
rect 28294 -20372 28341 -20308
rect 28405 -20372 28421 -20308
rect 28294 -20388 28421 -20372
rect 28294 -20452 28341 -20388
rect 28405 -20452 28421 -20388
rect 28294 -20468 28421 -20452
rect 28294 -20532 28341 -20468
rect 28405 -20532 28421 -20468
rect 28294 -20548 28421 -20532
rect 28294 -20612 28341 -20548
rect 28405 -20612 28421 -20548
rect 28294 -20628 28421 -20612
rect 28294 -20692 28341 -20628
rect 28405 -20692 28421 -20628
rect 28294 -20708 28421 -20692
rect 28294 -20772 28341 -20708
rect 28405 -20772 28421 -20708
rect 28294 -20788 28421 -20772
rect 28294 -20852 28341 -20788
rect 28405 -20852 28421 -20788
rect 28294 -20868 28421 -20852
rect 28294 -20932 28341 -20868
rect 28405 -20932 28421 -20868
rect 28294 -20948 28421 -20932
rect 28294 -21012 28341 -20948
rect 28405 -21012 28421 -20948
rect 28294 -21028 28421 -21012
rect 28294 -21092 28341 -21028
rect 28405 -21092 28421 -21028
rect 28294 -21108 28421 -21092
rect 28294 -21172 28341 -21108
rect 28405 -21172 28421 -21108
rect 28294 -21188 28421 -21172
rect 28294 -21252 28341 -21188
rect 28405 -21252 28421 -21188
rect 28294 -21268 28421 -21252
rect 28294 -21332 28341 -21268
rect 28405 -21332 28421 -21268
rect 28294 -21348 28421 -21332
rect 28294 -21412 28341 -21348
rect 28405 -21412 28421 -21348
rect 28294 -21428 28421 -21412
rect 28294 -21492 28341 -21428
rect 28405 -21492 28421 -21428
rect 28294 -21508 28421 -21492
rect 28294 -21572 28341 -21508
rect 28405 -21572 28421 -21508
rect 28294 -21588 28421 -21572
rect 28294 -21652 28341 -21588
rect 28405 -21652 28421 -21588
rect 28294 -21668 28421 -21652
rect 28294 -21732 28341 -21668
rect 28405 -21732 28421 -21668
rect 28294 -21748 28421 -21732
rect 28294 -21812 28341 -21748
rect 28405 -21812 28421 -21748
rect 28294 -21828 28421 -21812
rect 21975 -21908 22102 -21892
rect 21975 -21972 22022 -21908
rect 22086 -21972 22102 -21908
rect 21975 -21988 22102 -21972
rect 21975 -22112 22079 -21988
rect 21975 -22128 22102 -22112
rect 21975 -22192 22022 -22128
rect 22086 -22192 22102 -22128
rect 21975 -22208 22102 -22192
rect 15656 -22288 15783 -22272
rect 15656 -22352 15703 -22288
rect 15767 -22352 15783 -22288
rect 15656 -22368 15783 -22352
rect 15656 -22432 15703 -22368
rect 15767 -22432 15783 -22368
rect 15656 -22448 15783 -22432
rect 15656 -22512 15703 -22448
rect 15767 -22512 15783 -22448
rect 15656 -22528 15783 -22512
rect 15656 -22592 15703 -22528
rect 15767 -22592 15783 -22528
rect 15656 -22608 15783 -22592
rect 15656 -22672 15703 -22608
rect 15767 -22672 15783 -22608
rect 15656 -22688 15783 -22672
rect 15656 -22752 15703 -22688
rect 15767 -22752 15783 -22688
rect 15656 -22768 15783 -22752
rect 15656 -22832 15703 -22768
rect 15767 -22832 15783 -22768
rect 15656 -22848 15783 -22832
rect 15656 -22912 15703 -22848
rect 15767 -22912 15783 -22848
rect 15656 -22928 15783 -22912
rect 15656 -22992 15703 -22928
rect 15767 -22992 15783 -22928
rect 15656 -23008 15783 -22992
rect 15656 -23072 15703 -23008
rect 15767 -23072 15783 -23008
rect 15656 -23088 15783 -23072
rect 15656 -23152 15703 -23088
rect 15767 -23152 15783 -23088
rect 15656 -23168 15783 -23152
rect 15656 -23232 15703 -23168
rect 15767 -23232 15783 -23168
rect 15656 -23248 15783 -23232
rect 15656 -23312 15703 -23248
rect 15767 -23312 15783 -23248
rect 15656 -23328 15783 -23312
rect 15656 -23392 15703 -23328
rect 15767 -23392 15783 -23328
rect 15656 -23408 15783 -23392
rect 15656 -23472 15703 -23408
rect 15767 -23472 15783 -23408
rect 15656 -23488 15783 -23472
rect 15656 -23552 15703 -23488
rect 15767 -23552 15783 -23488
rect 15656 -23568 15783 -23552
rect 15656 -23632 15703 -23568
rect 15767 -23632 15783 -23568
rect 15656 -23648 15783 -23632
rect 15656 -23712 15703 -23648
rect 15767 -23712 15783 -23648
rect 15656 -23728 15783 -23712
rect 15656 -23792 15703 -23728
rect 15767 -23792 15783 -23728
rect 15656 -23808 15783 -23792
rect 15656 -23872 15703 -23808
rect 15767 -23872 15783 -23808
rect 15656 -23888 15783 -23872
rect 15656 -23952 15703 -23888
rect 15767 -23952 15783 -23888
rect 15656 -23968 15783 -23952
rect 15656 -24032 15703 -23968
rect 15767 -24032 15783 -23968
rect 15656 -24048 15783 -24032
rect 15656 -24112 15703 -24048
rect 15767 -24112 15783 -24048
rect 15656 -24128 15783 -24112
rect 15656 -24192 15703 -24128
rect 15767 -24192 15783 -24128
rect 15656 -24208 15783 -24192
rect 15656 -24272 15703 -24208
rect 15767 -24272 15783 -24208
rect 15656 -24288 15783 -24272
rect 15656 -24352 15703 -24288
rect 15767 -24352 15783 -24288
rect 15656 -24368 15783 -24352
rect 15656 -24432 15703 -24368
rect 15767 -24432 15783 -24368
rect 15656 -24448 15783 -24432
rect 15656 -24512 15703 -24448
rect 15767 -24512 15783 -24448
rect 15656 -24528 15783 -24512
rect 15656 -24592 15703 -24528
rect 15767 -24592 15783 -24528
rect 15656 -24608 15783 -24592
rect 15656 -24672 15703 -24608
rect 15767 -24672 15783 -24608
rect 15656 -24688 15783 -24672
rect 15656 -24752 15703 -24688
rect 15767 -24752 15783 -24688
rect 15656 -24768 15783 -24752
rect 15656 -24832 15703 -24768
rect 15767 -24832 15783 -24768
rect 15656 -24848 15783 -24832
rect 15656 -24912 15703 -24848
rect 15767 -24912 15783 -24848
rect 15656 -24928 15783 -24912
rect 15656 -24992 15703 -24928
rect 15767 -24992 15783 -24928
rect 15656 -25008 15783 -24992
rect 15656 -25072 15703 -25008
rect 15767 -25072 15783 -25008
rect 15656 -25088 15783 -25072
rect 15656 -25152 15703 -25088
rect 15767 -25152 15783 -25088
rect 15656 -25168 15783 -25152
rect 15656 -25232 15703 -25168
rect 15767 -25232 15783 -25168
rect 15656 -25248 15783 -25232
rect 15656 -25312 15703 -25248
rect 15767 -25312 15783 -25248
rect 15656 -25328 15783 -25312
rect 15656 -25392 15703 -25328
rect 15767 -25392 15783 -25328
rect 15656 -25408 15783 -25392
rect 15656 -25472 15703 -25408
rect 15767 -25472 15783 -25408
rect 15656 -25488 15783 -25472
rect 15656 -25552 15703 -25488
rect 15767 -25552 15783 -25488
rect 15656 -25568 15783 -25552
rect 15656 -25632 15703 -25568
rect 15767 -25632 15783 -25568
rect 15656 -25648 15783 -25632
rect 15656 -25712 15703 -25648
rect 15767 -25712 15783 -25648
rect 15656 -25728 15783 -25712
rect 15656 -25792 15703 -25728
rect 15767 -25792 15783 -25728
rect 15656 -25808 15783 -25792
rect 15656 -25872 15703 -25808
rect 15767 -25872 15783 -25808
rect 15656 -25888 15783 -25872
rect 15656 -25952 15703 -25888
rect 15767 -25952 15783 -25888
rect 15656 -25968 15783 -25952
rect 15656 -26032 15703 -25968
rect 15767 -26032 15783 -25968
rect 15656 -26048 15783 -26032
rect 15656 -26112 15703 -26048
rect 15767 -26112 15783 -26048
rect 15656 -26128 15783 -26112
rect 15656 -26192 15703 -26128
rect 15767 -26192 15783 -26128
rect 15656 -26208 15783 -26192
rect 15656 -26272 15703 -26208
rect 15767 -26272 15783 -26208
rect 15656 -26288 15783 -26272
rect 15656 -26352 15703 -26288
rect 15767 -26352 15783 -26288
rect 15656 -26368 15783 -26352
rect 15656 -26432 15703 -26368
rect 15767 -26432 15783 -26368
rect 15656 -26448 15783 -26432
rect 15656 -26512 15703 -26448
rect 15767 -26512 15783 -26448
rect 15656 -26528 15783 -26512
rect 15656 -26592 15703 -26528
rect 15767 -26592 15783 -26528
rect 15656 -26608 15783 -26592
rect 15656 -26672 15703 -26608
rect 15767 -26672 15783 -26608
rect 15656 -26688 15783 -26672
rect 15656 -26752 15703 -26688
rect 15767 -26752 15783 -26688
rect 15656 -26768 15783 -26752
rect 15656 -26832 15703 -26768
rect 15767 -26832 15783 -26768
rect 15656 -26848 15783 -26832
rect 15656 -26912 15703 -26848
rect 15767 -26912 15783 -26848
rect 15656 -26928 15783 -26912
rect 15656 -26992 15703 -26928
rect 15767 -26992 15783 -26928
rect 15656 -27008 15783 -26992
rect 15656 -27072 15703 -27008
rect 15767 -27072 15783 -27008
rect 15656 -27088 15783 -27072
rect 15656 -27152 15703 -27088
rect 15767 -27152 15783 -27088
rect 15656 -27168 15783 -27152
rect 15656 -27232 15703 -27168
rect 15767 -27232 15783 -27168
rect 15656 -27248 15783 -27232
rect 15656 -27312 15703 -27248
rect 15767 -27312 15783 -27248
rect 15656 -27328 15783 -27312
rect 15656 -27392 15703 -27328
rect 15767 -27392 15783 -27328
rect 15656 -27408 15783 -27392
rect 15656 -27472 15703 -27408
rect 15767 -27472 15783 -27408
rect 15656 -27488 15783 -27472
rect 15656 -27552 15703 -27488
rect 15767 -27552 15783 -27488
rect 15656 -27568 15783 -27552
rect 15656 -27632 15703 -27568
rect 15767 -27632 15783 -27568
rect 15656 -27648 15783 -27632
rect 15656 -27712 15703 -27648
rect 15767 -27712 15783 -27648
rect 15656 -27728 15783 -27712
rect 15656 -27792 15703 -27728
rect 15767 -27792 15783 -27728
rect 15656 -27808 15783 -27792
rect 15656 -27872 15703 -27808
rect 15767 -27872 15783 -27808
rect 15656 -27888 15783 -27872
rect 15656 -27952 15703 -27888
rect 15767 -27952 15783 -27888
rect 15656 -27968 15783 -27952
rect 15656 -28032 15703 -27968
rect 15767 -28032 15783 -27968
rect 15656 -28048 15783 -28032
rect 15656 -28112 15703 -28048
rect 15767 -28112 15783 -28048
rect 15656 -28128 15783 -28112
rect 9337 -28208 9464 -28192
rect 9337 -28272 9384 -28208
rect 9448 -28272 9464 -28208
rect 9337 -28288 9464 -28272
rect 9337 -28412 9441 -28288
rect 9337 -28428 9464 -28412
rect 9337 -28492 9384 -28428
rect 9448 -28492 9464 -28428
rect 9337 -28508 9464 -28492
rect 3018 -28588 3145 -28572
rect 3018 -28652 3065 -28588
rect 3129 -28652 3145 -28588
rect 3018 -28668 3145 -28652
rect 3018 -28732 3065 -28668
rect 3129 -28732 3145 -28668
rect 3018 -28748 3145 -28732
rect 3018 -28812 3065 -28748
rect 3129 -28812 3145 -28748
rect 3018 -28828 3145 -28812
rect 3018 -28892 3065 -28828
rect 3129 -28892 3145 -28828
rect 3018 -28908 3145 -28892
rect 3018 -28972 3065 -28908
rect 3129 -28972 3145 -28908
rect 3018 -28988 3145 -28972
rect 3018 -29052 3065 -28988
rect 3129 -29052 3145 -28988
rect 3018 -29068 3145 -29052
rect 3018 -29132 3065 -29068
rect 3129 -29132 3145 -29068
rect 3018 -29148 3145 -29132
rect 3018 -29212 3065 -29148
rect 3129 -29212 3145 -29148
rect 3018 -29228 3145 -29212
rect 3018 -29292 3065 -29228
rect 3129 -29292 3145 -29228
rect 3018 -29308 3145 -29292
rect 3018 -29372 3065 -29308
rect 3129 -29372 3145 -29308
rect 3018 -29388 3145 -29372
rect 3018 -29452 3065 -29388
rect 3129 -29452 3145 -29388
rect 3018 -29468 3145 -29452
rect 3018 -29532 3065 -29468
rect 3129 -29532 3145 -29468
rect 3018 -29548 3145 -29532
rect 3018 -29612 3065 -29548
rect 3129 -29612 3145 -29548
rect 3018 -29628 3145 -29612
rect 3018 -29692 3065 -29628
rect 3129 -29692 3145 -29628
rect 3018 -29708 3145 -29692
rect 3018 -29772 3065 -29708
rect 3129 -29772 3145 -29708
rect 3018 -29788 3145 -29772
rect 3018 -29852 3065 -29788
rect 3129 -29852 3145 -29788
rect 3018 -29868 3145 -29852
rect 3018 -29932 3065 -29868
rect 3129 -29932 3145 -29868
rect 3018 -29948 3145 -29932
rect 3018 -30012 3065 -29948
rect 3129 -30012 3145 -29948
rect 3018 -30028 3145 -30012
rect 3018 -30092 3065 -30028
rect 3129 -30092 3145 -30028
rect 3018 -30108 3145 -30092
rect 3018 -30172 3065 -30108
rect 3129 -30172 3145 -30108
rect 3018 -30188 3145 -30172
rect 3018 -30252 3065 -30188
rect 3129 -30252 3145 -30188
rect 3018 -30268 3145 -30252
rect 3018 -30332 3065 -30268
rect 3129 -30332 3145 -30268
rect 3018 -30348 3145 -30332
rect 3018 -30412 3065 -30348
rect 3129 -30412 3145 -30348
rect 3018 -30428 3145 -30412
rect 3018 -30492 3065 -30428
rect 3129 -30492 3145 -30428
rect 3018 -30508 3145 -30492
rect 3018 -30572 3065 -30508
rect 3129 -30572 3145 -30508
rect 3018 -30588 3145 -30572
rect 3018 -30652 3065 -30588
rect 3129 -30652 3145 -30588
rect 3018 -30668 3145 -30652
rect 3018 -30732 3065 -30668
rect 3129 -30732 3145 -30668
rect 3018 -30748 3145 -30732
rect 3018 -30812 3065 -30748
rect 3129 -30812 3145 -30748
rect 3018 -30828 3145 -30812
rect 3018 -30892 3065 -30828
rect 3129 -30892 3145 -30828
rect 3018 -30908 3145 -30892
rect 3018 -30972 3065 -30908
rect 3129 -30972 3145 -30908
rect 3018 -30988 3145 -30972
rect 3018 -31052 3065 -30988
rect 3129 -31052 3145 -30988
rect 3018 -31068 3145 -31052
rect 3018 -31132 3065 -31068
rect 3129 -31132 3145 -31068
rect 3018 -31148 3145 -31132
rect 3018 -31212 3065 -31148
rect 3129 -31212 3145 -31148
rect 3018 -31228 3145 -31212
rect 3018 -31292 3065 -31228
rect 3129 -31292 3145 -31228
rect 3018 -31308 3145 -31292
rect 3018 -31372 3065 -31308
rect 3129 -31372 3145 -31308
rect 3018 -31388 3145 -31372
rect 3018 -31452 3065 -31388
rect 3129 -31452 3145 -31388
rect 3018 -31468 3145 -31452
rect 3018 -31532 3065 -31468
rect 3129 -31532 3145 -31468
rect 3018 -31548 3145 -31532
rect 3018 -31612 3065 -31548
rect 3129 -31612 3145 -31548
rect 3018 -31628 3145 -31612
rect 3018 -31692 3065 -31628
rect 3129 -31692 3145 -31628
rect 3018 -31708 3145 -31692
rect 3018 -31772 3065 -31708
rect 3129 -31772 3145 -31708
rect 3018 -31788 3145 -31772
rect 3018 -31852 3065 -31788
rect 3129 -31852 3145 -31788
rect 3018 -31868 3145 -31852
rect 3018 -31932 3065 -31868
rect 3129 -31932 3145 -31868
rect 3018 -31948 3145 -31932
rect 3018 -32012 3065 -31948
rect 3129 -32012 3145 -31948
rect 3018 -32028 3145 -32012
rect 3018 -32092 3065 -32028
rect 3129 -32092 3145 -32028
rect 3018 -32108 3145 -32092
rect 3018 -32172 3065 -32108
rect 3129 -32172 3145 -32108
rect 3018 -32188 3145 -32172
rect 3018 -32252 3065 -32188
rect 3129 -32252 3145 -32188
rect 3018 -32268 3145 -32252
rect 3018 -32332 3065 -32268
rect 3129 -32332 3145 -32268
rect 3018 -32348 3145 -32332
rect 3018 -32412 3065 -32348
rect 3129 -32412 3145 -32348
rect 3018 -32428 3145 -32412
rect 3018 -32492 3065 -32428
rect 3129 -32492 3145 -32428
rect 3018 -32508 3145 -32492
rect 3018 -32572 3065 -32508
rect 3129 -32572 3145 -32508
rect 3018 -32588 3145 -32572
rect 3018 -32652 3065 -32588
rect 3129 -32652 3145 -32588
rect 3018 -32668 3145 -32652
rect 3018 -32732 3065 -32668
rect 3129 -32732 3145 -32668
rect 3018 -32748 3145 -32732
rect 3018 -32812 3065 -32748
rect 3129 -32812 3145 -32748
rect 3018 -32828 3145 -32812
rect 3018 -32892 3065 -32828
rect 3129 -32892 3145 -32828
rect 3018 -32908 3145 -32892
rect 3018 -32972 3065 -32908
rect 3129 -32972 3145 -32908
rect 3018 -32988 3145 -32972
rect 3018 -33052 3065 -32988
rect 3129 -33052 3145 -32988
rect 3018 -33068 3145 -33052
rect 3018 -33132 3065 -33068
rect 3129 -33132 3145 -33068
rect 3018 -33148 3145 -33132
rect 3018 -33212 3065 -33148
rect 3129 -33212 3145 -33148
rect 3018 -33228 3145 -33212
rect 3018 -33292 3065 -33228
rect 3129 -33292 3145 -33228
rect 3018 -33308 3145 -33292
rect 3018 -33372 3065 -33308
rect 3129 -33372 3145 -33308
rect 3018 -33388 3145 -33372
rect 3018 -33452 3065 -33388
rect 3129 -33452 3145 -33388
rect 3018 -33468 3145 -33452
rect 3018 -33532 3065 -33468
rect 3129 -33532 3145 -33468
rect 3018 -33548 3145 -33532
rect 3018 -33612 3065 -33548
rect 3129 -33612 3145 -33548
rect 3018 -33628 3145 -33612
rect 3018 -33692 3065 -33628
rect 3129 -33692 3145 -33628
rect 3018 -33708 3145 -33692
rect 3018 -33772 3065 -33708
rect 3129 -33772 3145 -33708
rect 3018 -33788 3145 -33772
rect 3018 -33852 3065 -33788
rect 3129 -33852 3145 -33788
rect 3018 -33868 3145 -33852
rect 3018 -33932 3065 -33868
rect 3129 -33932 3145 -33868
rect 3018 -33948 3145 -33932
rect 3018 -34012 3065 -33948
rect 3129 -34012 3145 -33948
rect 3018 -34028 3145 -34012
rect 3018 -34092 3065 -34028
rect 3129 -34092 3145 -34028
rect 3018 -34108 3145 -34092
rect 3018 -34172 3065 -34108
rect 3129 -34172 3145 -34108
rect 3018 -34188 3145 -34172
rect 3018 -34252 3065 -34188
rect 3129 -34252 3145 -34188
rect 3018 -34268 3145 -34252
rect 3018 -34332 3065 -34268
rect 3129 -34332 3145 -34268
rect 3018 -34348 3145 -34332
rect 3018 -34412 3065 -34348
rect 3129 -34412 3145 -34348
rect 3018 -34428 3145 -34412
rect -3301 -34508 -3174 -34492
rect -3301 -34572 -3254 -34508
rect -3190 -34572 -3174 -34508
rect -3301 -34588 -3174 -34572
rect -3301 -34712 -3197 -34588
rect -3301 -34728 -3174 -34712
rect -3301 -34792 -3254 -34728
rect -3190 -34792 -3174 -34728
rect -3301 -34808 -3174 -34792
rect -9620 -34888 -9493 -34872
rect -9620 -34952 -9573 -34888
rect -9509 -34952 -9493 -34888
rect -9620 -34968 -9493 -34952
rect -9620 -35032 -9573 -34968
rect -9509 -35032 -9493 -34968
rect -9620 -35048 -9493 -35032
rect -9620 -35112 -9573 -35048
rect -9509 -35112 -9493 -35048
rect -9620 -35128 -9493 -35112
rect -9620 -35192 -9573 -35128
rect -9509 -35192 -9493 -35128
rect -9620 -35208 -9493 -35192
rect -9620 -35272 -9573 -35208
rect -9509 -35272 -9493 -35208
rect -9620 -35288 -9493 -35272
rect -9620 -35352 -9573 -35288
rect -9509 -35352 -9493 -35288
rect -9620 -35368 -9493 -35352
rect -9620 -35432 -9573 -35368
rect -9509 -35432 -9493 -35368
rect -9620 -35448 -9493 -35432
rect -9620 -35512 -9573 -35448
rect -9509 -35512 -9493 -35448
rect -9620 -35528 -9493 -35512
rect -9620 -35592 -9573 -35528
rect -9509 -35592 -9493 -35528
rect -9620 -35608 -9493 -35592
rect -9620 -35672 -9573 -35608
rect -9509 -35672 -9493 -35608
rect -9620 -35688 -9493 -35672
rect -9620 -35752 -9573 -35688
rect -9509 -35752 -9493 -35688
rect -9620 -35768 -9493 -35752
rect -9620 -35832 -9573 -35768
rect -9509 -35832 -9493 -35768
rect -9620 -35848 -9493 -35832
rect -9620 -35912 -9573 -35848
rect -9509 -35912 -9493 -35848
rect -9620 -35928 -9493 -35912
rect -9620 -35992 -9573 -35928
rect -9509 -35992 -9493 -35928
rect -9620 -36008 -9493 -35992
rect -9620 -36072 -9573 -36008
rect -9509 -36072 -9493 -36008
rect -9620 -36088 -9493 -36072
rect -9620 -36152 -9573 -36088
rect -9509 -36152 -9493 -36088
rect -9620 -36168 -9493 -36152
rect -9620 -36232 -9573 -36168
rect -9509 -36232 -9493 -36168
rect -9620 -36248 -9493 -36232
rect -9620 -36312 -9573 -36248
rect -9509 -36312 -9493 -36248
rect -9620 -36328 -9493 -36312
rect -9620 -36392 -9573 -36328
rect -9509 -36392 -9493 -36328
rect -9620 -36408 -9493 -36392
rect -9620 -36472 -9573 -36408
rect -9509 -36472 -9493 -36408
rect -9620 -36488 -9493 -36472
rect -9620 -36552 -9573 -36488
rect -9509 -36552 -9493 -36488
rect -9620 -36568 -9493 -36552
rect -9620 -36632 -9573 -36568
rect -9509 -36632 -9493 -36568
rect -9620 -36648 -9493 -36632
rect -9620 -36712 -9573 -36648
rect -9509 -36712 -9493 -36648
rect -9620 -36728 -9493 -36712
rect -9620 -36792 -9573 -36728
rect -9509 -36792 -9493 -36728
rect -9620 -36808 -9493 -36792
rect -9620 -36872 -9573 -36808
rect -9509 -36872 -9493 -36808
rect -9620 -36888 -9493 -36872
rect -9620 -36952 -9573 -36888
rect -9509 -36952 -9493 -36888
rect -9620 -36968 -9493 -36952
rect -9620 -37032 -9573 -36968
rect -9509 -37032 -9493 -36968
rect -9620 -37048 -9493 -37032
rect -9620 -37112 -9573 -37048
rect -9509 -37112 -9493 -37048
rect -9620 -37128 -9493 -37112
rect -9620 -37192 -9573 -37128
rect -9509 -37192 -9493 -37128
rect -9620 -37208 -9493 -37192
rect -9620 -37272 -9573 -37208
rect -9509 -37272 -9493 -37208
rect -9620 -37288 -9493 -37272
rect -9620 -37352 -9573 -37288
rect -9509 -37352 -9493 -37288
rect -9620 -37368 -9493 -37352
rect -9620 -37432 -9573 -37368
rect -9509 -37432 -9493 -37368
rect -9620 -37448 -9493 -37432
rect -9620 -37512 -9573 -37448
rect -9509 -37512 -9493 -37448
rect -9620 -37528 -9493 -37512
rect -9620 -37592 -9573 -37528
rect -9509 -37592 -9493 -37528
rect -9620 -37608 -9493 -37592
rect -9620 -37672 -9573 -37608
rect -9509 -37672 -9493 -37608
rect -9620 -37688 -9493 -37672
rect -9620 -37752 -9573 -37688
rect -9509 -37752 -9493 -37688
rect -9620 -37768 -9493 -37752
rect -9620 -37832 -9573 -37768
rect -9509 -37832 -9493 -37768
rect -9620 -37848 -9493 -37832
rect -9620 -37912 -9573 -37848
rect -9509 -37912 -9493 -37848
rect -9620 -37928 -9493 -37912
rect -9620 -37992 -9573 -37928
rect -9509 -37992 -9493 -37928
rect -9620 -38008 -9493 -37992
rect -9620 -38072 -9573 -38008
rect -9509 -38072 -9493 -38008
rect -9620 -38088 -9493 -38072
rect -9620 -38152 -9573 -38088
rect -9509 -38152 -9493 -38088
rect -9620 -38168 -9493 -38152
rect -9620 -38232 -9573 -38168
rect -9509 -38232 -9493 -38168
rect -9620 -38248 -9493 -38232
rect -9620 -38312 -9573 -38248
rect -9509 -38312 -9493 -38248
rect -9620 -38328 -9493 -38312
rect -9620 -38392 -9573 -38328
rect -9509 -38392 -9493 -38328
rect -9620 -38408 -9493 -38392
rect -9620 -38472 -9573 -38408
rect -9509 -38472 -9493 -38408
rect -9620 -38488 -9493 -38472
rect -9620 -38552 -9573 -38488
rect -9509 -38552 -9493 -38488
rect -9620 -38568 -9493 -38552
rect -9620 -38632 -9573 -38568
rect -9509 -38632 -9493 -38568
rect -9620 -38648 -9493 -38632
rect -9620 -38712 -9573 -38648
rect -9509 -38712 -9493 -38648
rect -9620 -38728 -9493 -38712
rect -9620 -38792 -9573 -38728
rect -9509 -38792 -9493 -38728
rect -9620 -38808 -9493 -38792
rect -9620 -38872 -9573 -38808
rect -9509 -38872 -9493 -38808
rect -9620 -38888 -9493 -38872
rect -9620 -38952 -9573 -38888
rect -9509 -38952 -9493 -38888
rect -9620 -38968 -9493 -38952
rect -9620 -39032 -9573 -38968
rect -9509 -39032 -9493 -38968
rect -9620 -39048 -9493 -39032
rect -9620 -39112 -9573 -39048
rect -9509 -39112 -9493 -39048
rect -9620 -39128 -9493 -39112
rect -9620 -39192 -9573 -39128
rect -9509 -39192 -9493 -39128
rect -9620 -39208 -9493 -39192
rect -9620 -39272 -9573 -39208
rect -9509 -39272 -9493 -39208
rect -9620 -39288 -9493 -39272
rect -9620 -39352 -9573 -39288
rect -9509 -39352 -9493 -39288
rect -9620 -39368 -9493 -39352
rect -9620 -39432 -9573 -39368
rect -9509 -39432 -9493 -39368
rect -9620 -39448 -9493 -39432
rect -9620 -39512 -9573 -39448
rect -9509 -39512 -9493 -39448
rect -9620 -39528 -9493 -39512
rect -9620 -39592 -9573 -39528
rect -9509 -39592 -9493 -39528
rect -9620 -39608 -9493 -39592
rect -9620 -39672 -9573 -39608
rect -9509 -39672 -9493 -39608
rect -9620 -39688 -9493 -39672
rect -9620 -39752 -9573 -39688
rect -9509 -39752 -9493 -39688
rect -9620 -39768 -9493 -39752
rect -9620 -39832 -9573 -39768
rect -9509 -39832 -9493 -39768
rect -9620 -39848 -9493 -39832
rect -9620 -39912 -9573 -39848
rect -9509 -39912 -9493 -39848
rect -9620 -39928 -9493 -39912
rect -9620 -39992 -9573 -39928
rect -9509 -39992 -9493 -39928
rect -9620 -40008 -9493 -39992
rect -9620 -40072 -9573 -40008
rect -9509 -40072 -9493 -40008
rect -9620 -40088 -9493 -40072
rect -9620 -40152 -9573 -40088
rect -9509 -40152 -9493 -40088
rect -9620 -40168 -9493 -40152
rect -9620 -40232 -9573 -40168
rect -9509 -40232 -9493 -40168
rect -9620 -40248 -9493 -40232
rect -9620 -40312 -9573 -40248
rect -9509 -40312 -9493 -40248
rect -9620 -40328 -9493 -40312
rect -9620 -40392 -9573 -40328
rect -9509 -40392 -9493 -40328
rect -9620 -40408 -9493 -40392
rect -9620 -40472 -9573 -40408
rect -9509 -40472 -9493 -40408
rect -9620 -40488 -9493 -40472
rect -9620 -40552 -9573 -40488
rect -9509 -40552 -9493 -40488
rect -9620 -40568 -9493 -40552
rect -9620 -40632 -9573 -40568
rect -9509 -40632 -9493 -40568
rect -9620 -40648 -9493 -40632
rect -9620 -40712 -9573 -40648
rect -9509 -40712 -9493 -40648
rect -9620 -40728 -9493 -40712
rect -15939 -40808 -15812 -40792
rect -15939 -40872 -15892 -40808
rect -15828 -40872 -15812 -40808
rect -15939 -40888 -15812 -40872
rect -15939 -41012 -15835 -40888
rect -15939 -41028 -15812 -41012
rect -15939 -41092 -15892 -41028
rect -15828 -41092 -15812 -41028
rect -15939 -41108 -15812 -41092
rect -22258 -41188 -22131 -41172
rect -22258 -41252 -22211 -41188
rect -22147 -41252 -22131 -41188
rect -22258 -41268 -22131 -41252
rect -22258 -41332 -22211 -41268
rect -22147 -41332 -22131 -41268
rect -22258 -41348 -22131 -41332
rect -22258 -41412 -22211 -41348
rect -22147 -41412 -22131 -41348
rect -22258 -41428 -22131 -41412
rect -22258 -41492 -22211 -41428
rect -22147 -41492 -22131 -41428
rect -22258 -41508 -22131 -41492
rect -22258 -41572 -22211 -41508
rect -22147 -41572 -22131 -41508
rect -22258 -41588 -22131 -41572
rect -22258 -41652 -22211 -41588
rect -22147 -41652 -22131 -41588
rect -22258 -41668 -22131 -41652
rect -22258 -41732 -22211 -41668
rect -22147 -41732 -22131 -41668
rect -22258 -41748 -22131 -41732
rect -22258 -41812 -22211 -41748
rect -22147 -41812 -22131 -41748
rect -22258 -41828 -22131 -41812
rect -22258 -41892 -22211 -41828
rect -22147 -41892 -22131 -41828
rect -22258 -41908 -22131 -41892
rect -22258 -41972 -22211 -41908
rect -22147 -41972 -22131 -41908
rect -22258 -41988 -22131 -41972
rect -22258 -42052 -22211 -41988
rect -22147 -42052 -22131 -41988
rect -22258 -42068 -22131 -42052
rect -22258 -42132 -22211 -42068
rect -22147 -42132 -22131 -42068
rect -22258 -42148 -22131 -42132
rect -22258 -42212 -22211 -42148
rect -22147 -42212 -22131 -42148
rect -22258 -42228 -22131 -42212
rect -22258 -42292 -22211 -42228
rect -22147 -42292 -22131 -42228
rect -22258 -42308 -22131 -42292
rect -22258 -42372 -22211 -42308
rect -22147 -42372 -22131 -42308
rect -22258 -42388 -22131 -42372
rect -22258 -42452 -22211 -42388
rect -22147 -42452 -22131 -42388
rect -22258 -42468 -22131 -42452
rect -22258 -42532 -22211 -42468
rect -22147 -42532 -22131 -42468
rect -22258 -42548 -22131 -42532
rect -22258 -42612 -22211 -42548
rect -22147 -42612 -22131 -42548
rect -22258 -42628 -22131 -42612
rect -22258 -42692 -22211 -42628
rect -22147 -42692 -22131 -42628
rect -22258 -42708 -22131 -42692
rect -22258 -42772 -22211 -42708
rect -22147 -42772 -22131 -42708
rect -22258 -42788 -22131 -42772
rect -22258 -42852 -22211 -42788
rect -22147 -42852 -22131 -42788
rect -22258 -42868 -22131 -42852
rect -22258 -42932 -22211 -42868
rect -22147 -42932 -22131 -42868
rect -22258 -42948 -22131 -42932
rect -22258 -43012 -22211 -42948
rect -22147 -43012 -22131 -42948
rect -22258 -43028 -22131 -43012
rect -22258 -43092 -22211 -43028
rect -22147 -43092 -22131 -43028
rect -22258 -43108 -22131 -43092
rect -22258 -43172 -22211 -43108
rect -22147 -43172 -22131 -43108
rect -22258 -43188 -22131 -43172
rect -22258 -43252 -22211 -43188
rect -22147 -43252 -22131 -43188
rect -22258 -43268 -22131 -43252
rect -22258 -43332 -22211 -43268
rect -22147 -43332 -22131 -43268
rect -22258 -43348 -22131 -43332
rect -22258 -43412 -22211 -43348
rect -22147 -43412 -22131 -43348
rect -22258 -43428 -22131 -43412
rect -22258 -43492 -22211 -43428
rect -22147 -43492 -22131 -43428
rect -22258 -43508 -22131 -43492
rect -22258 -43572 -22211 -43508
rect -22147 -43572 -22131 -43508
rect -22258 -43588 -22131 -43572
rect -22258 -43652 -22211 -43588
rect -22147 -43652 -22131 -43588
rect -22258 -43668 -22131 -43652
rect -22258 -43732 -22211 -43668
rect -22147 -43732 -22131 -43668
rect -22258 -43748 -22131 -43732
rect -22258 -43812 -22211 -43748
rect -22147 -43812 -22131 -43748
rect -22258 -43828 -22131 -43812
rect -22258 -43892 -22211 -43828
rect -22147 -43892 -22131 -43828
rect -22258 -43908 -22131 -43892
rect -22258 -43972 -22211 -43908
rect -22147 -43972 -22131 -43908
rect -22258 -43988 -22131 -43972
rect -22258 -44052 -22211 -43988
rect -22147 -44052 -22131 -43988
rect -22258 -44068 -22131 -44052
rect -22258 -44132 -22211 -44068
rect -22147 -44132 -22131 -44068
rect -22258 -44148 -22131 -44132
rect -22258 -44212 -22211 -44148
rect -22147 -44212 -22131 -44148
rect -22258 -44228 -22131 -44212
rect -22258 -44292 -22211 -44228
rect -22147 -44292 -22131 -44228
rect -22258 -44308 -22131 -44292
rect -22258 -44372 -22211 -44308
rect -22147 -44372 -22131 -44308
rect -22258 -44388 -22131 -44372
rect -22258 -44452 -22211 -44388
rect -22147 -44452 -22131 -44388
rect -22258 -44468 -22131 -44452
rect -22258 -44532 -22211 -44468
rect -22147 -44532 -22131 -44468
rect -22258 -44548 -22131 -44532
rect -22258 -44612 -22211 -44548
rect -22147 -44612 -22131 -44548
rect -22258 -44628 -22131 -44612
rect -22258 -44692 -22211 -44628
rect -22147 -44692 -22131 -44628
rect -22258 -44708 -22131 -44692
rect -22258 -44772 -22211 -44708
rect -22147 -44772 -22131 -44708
rect -22258 -44788 -22131 -44772
rect -22258 -44852 -22211 -44788
rect -22147 -44852 -22131 -44788
rect -22258 -44868 -22131 -44852
rect -22258 -44932 -22211 -44868
rect -22147 -44932 -22131 -44868
rect -22258 -44948 -22131 -44932
rect -22258 -45012 -22211 -44948
rect -22147 -45012 -22131 -44948
rect -22258 -45028 -22131 -45012
rect -22258 -45092 -22211 -45028
rect -22147 -45092 -22131 -45028
rect -22258 -45108 -22131 -45092
rect -22258 -45172 -22211 -45108
rect -22147 -45172 -22131 -45108
rect -22258 -45188 -22131 -45172
rect -22258 -45252 -22211 -45188
rect -22147 -45252 -22131 -45188
rect -22258 -45268 -22131 -45252
rect -22258 -45332 -22211 -45268
rect -22147 -45332 -22131 -45268
rect -22258 -45348 -22131 -45332
rect -22258 -45412 -22211 -45348
rect -22147 -45412 -22131 -45348
rect -22258 -45428 -22131 -45412
rect -22258 -45492 -22211 -45428
rect -22147 -45492 -22131 -45428
rect -22258 -45508 -22131 -45492
rect -22258 -45572 -22211 -45508
rect -22147 -45572 -22131 -45508
rect -22258 -45588 -22131 -45572
rect -22258 -45652 -22211 -45588
rect -22147 -45652 -22131 -45588
rect -22258 -45668 -22131 -45652
rect -22258 -45732 -22211 -45668
rect -22147 -45732 -22131 -45668
rect -22258 -45748 -22131 -45732
rect -22258 -45812 -22211 -45748
rect -22147 -45812 -22131 -45748
rect -22258 -45828 -22131 -45812
rect -22258 -45892 -22211 -45828
rect -22147 -45892 -22131 -45828
rect -22258 -45908 -22131 -45892
rect -22258 -45972 -22211 -45908
rect -22147 -45972 -22131 -45908
rect -22258 -45988 -22131 -45972
rect -22258 -46052 -22211 -45988
rect -22147 -46052 -22131 -45988
rect -22258 -46068 -22131 -46052
rect -22258 -46132 -22211 -46068
rect -22147 -46132 -22131 -46068
rect -22258 -46148 -22131 -46132
rect -22258 -46212 -22211 -46148
rect -22147 -46212 -22131 -46148
rect -22258 -46228 -22131 -46212
rect -22258 -46292 -22211 -46228
rect -22147 -46292 -22131 -46228
rect -22258 -46308 -22131 -46292
rect -22258 -46372 -22211 -46308
rect -22147 -46372 -22131 -46308
rect -22258 -46388 -22131 -46372
rect -22258 -46452 -22211 -46388
rect -22147 -46452 -22131 -46388
rect -22258 -46468 -22131 -46452
rect -22258 -46532 -22211 -46468
rect -22147 -46532 -22131 -46468
rect -22258 -46548 -22131 -46532
rect -22258 -46612 -22211 -46548
rect -22147 -46612 -22131 -46548
rect -22258 -46628 -22131 -46612
rect -22258 -46692 -22211 -46628
rect -22147 -46692 -22131 -46628
rect -22258 -46708 -22131 -46692
rect -22258 -46772 -22211 -46708
rect -22147 -46772 -22131 -46708
rect -22258 -46788 -22131 -46772
rect -22258 -46852 -22211 -46788
rect -22147 -46852 -22131 -46788
rect -22258 -46868 -22131 -46852
rect -22258 -46932 -22211 -46868
rect -22147 -46932 -22131 -46868
rect -22258 -46948 -22131 -46932
rect -22258 -47012 -22211 -46948
rect -22147 -47012 -22131 -46948
rect -22258 -47028 -22131 -47012
rect -28577 -47108 -28450 -47092
rect -28577 -47172 -28530 -47108
rect -28466 -47172 -28450 -47108
rect -28577 -47188 -28450 -47172
rect -28577 -47250 -28473 -47188
rect -25378 -47250 -25274 -47061
rect -22258 -47092 -22211 -47028
rect -22147 -47092 -22131 -47028
rect -21968 -41148 -16046 -41139
rect -21968 -47052 -21959 -41148
rect -16055 -47052 -16046 -41148
rect -21968 -47061 -16046 -47052
rect -15939 -41172 -15892 -41108
rect -15828 -41172 -15812 -41108
rect -12740 -41139 -12636 -40761
rect -9620 -40792 -9573 -40728
rect -9509 -40792 -9493 -40728
rect -9330 -34848 -3408 -34839
rect -9330 -40752 -9321 -34848
rect -3417 -40752 -3408 -34848
rect -9330 -40761 -3408 -40752
rect -3301 -34872 -3254 -34808
rect -3190 -34872 -3174 -34808
rect -102 -34839 2 -34461
rect 3018 -34492 3065 -34428
rect 3129 -34492 3145 -34428
rect 3308 -28548 9230 -28539
rect 3308 -34452 3317 -28548
rect 9221 -34452 9230 -28548
rect 3308 -34461 9230 -34452
rect 9337 -28572 9384 -28508
rect 9448 -28572 9464 -28508
rect 12536 -28539 12640 -28161
rect 15656 -28192 15703 -28128
rect 15767 -28192 15783 -28128
rect 15946 -22248 21868 -22239
rect 15946 -28152 15955 -22248
rect 21859 -28152 21868 -22248
rect 15946 -28161 21868 -28152
rect 21975 -22272 22022 -22208
rect 22086 -22272 22102 -22208
rect 25174 -22239 25278 -21861
rect 28294 -21892 28341 -21828
rect 28405 -21892 28421 -21828
rect 28584 -15948 34506 -15939
rect 28584 -21852 28593 -15948
rect 34497 -21852 34506 -15948
rect 28584 -21861 34506 -21852
rect 34613 -15972 34660 -15908
rect 34724 -15972 34740 -15908
rect 37812 -15939 37916 -15561
rect 40932 -15592 40979 -15528
rect 41043 -15592 41059 -15528
rect 41222 -9648 47144 -9639
rect 41222 -15552 41231 -9648
rect 47135 -15552 47144 -9648
rect 41222 -15561 47144 -15552
rect 47251 -9672 47298 -9608
rect 47362 -9672 47378 -9608
rect 47251 -9688 47378 -9672
rect 47251 -9752 47298 -9688
rect 47362 -9752 47378 -9688
rect 47251 -9768 47378 -9752
rect 47251 -9832 47298 -9768
rect 47362 -9832 47378 -9768
rect 47251 -9848 47378 -9832
rect 47251 -9912 47298 -9848
rect 47362 -9912 47378 -9848
rect 47251 -9928 47378 -9912
rect 47251 -9992 47298 -9928
rect 47362 -9992 47378 -9928
rect 47251 -10008 47378 -9992
rect 47251 -10072 47298 -10008
rect 47362 -10072 47378 -10008
rect 47251 -10088 47378 -10072
rect 47251 -10152 47298 -10088
rect 47362 -10152 47378 -10088
rect 47251 -10168 47378 -10152
rect 47251 -10232 47298 -10168
rect 47362 -10232 47378 -10168
rect 47251 -10248 47378 -10232
rect 47251 -10312 47298 -10248
rect 47362 -10312 47378 -10248
rect 47251 -10328 47378 -10312
rect 47251 -10392 47298 -10328
rect 47362 -10392 47378 -10328
rect 47251 -10408 47378 -10392
rect 47251 -10472 47298 -10408
rect 47362 -10472 47378 -10408
rect 47251 -10488 47378 -10472
rect 47251 -10552 47298 -10488
rect 47362 -10552 47378 -10488
rect 47251 -10568 47378 -10552
rect 47251 -10632 47298 -10568
rect 47362 -10632 47378 -10568
rect 47251 -10648 47378 -10632
rect 47251 -10712 47298 -10648
rect 47362 -10712 47378 -10648
rect 47251 -10728 47378 -10712
rect 47251 -10792 47298 -10728
rect 47362 -10792 47378 -10728
rect 47251 -10808 47378 -10792
rect 47251 -10872 47298 -10808
rect 47362 -10872 47378 -10808
rect 47251 -10888 47378 -10872
rect 47251 -10952 47298 -10888
rect 47362 -10952 47378 -10888
rect 47251 -10968 47378 -10952
rect 47251 -11032 47298 -10968
rect 47362 -11032 47378 -10968
rect 47251 -11048 47378 -11032
rect 47251 -11112 47298 -11048
rect 47362 -11112 47378 -11048
rect 47251 -11128 47378 -11112
rect 47251 -11192 47298 -11128
rect 47362 -11192 47378 -11128
rect 47251 -11208 47378 -11192
rect 47251 -11272 47298 -11208
rect 47362 -11272 47378 -11208
rect 47251 -11288 47378 -11272
rect 47251 -11352 47298 -11288
rect 47362 -11352 47378 -11288
rect 47251 -11368 47378 -11352
rect 47251 -11432 47298 -11368
rect 47362 -11432 47378 -11368
rect 47251 -11448 47378 -11432
rect 47251 -11512 47298 -11448
rect 47362 -11512 47378 -11448
rect 47251 -11528 47378 -11512
rect 47251 -11592 47298 -11528
rect 47362 -11592 47378 -11528
rect 47251 -11608 47378 -11592
rect 47251 -11672 47298 -11608
rect 47362 -11672 47378 -11608
rect 47251 -11688 47378 -11672
rect 47251 -11752 47298 -11688
rect 47362 -11752 47378 -11688
rect 47251 -11768 47378 -11752
rect 47251 -11832 47298 -11768
rect 47362 -11832 47378 -11768
rect 47251 -11848 47378 -11832
rect 47251 -11912 47298 -11848
rect 47362 -11912 47378 -11848
rect 47251 -11928 47378 -11912
rect 47251 -11992 47298 -11928
rect 47362 -11992 47378 -11928
rect 47251 -12008 47378 -11992
rect 47251 -12072 47298 -12008
rect 47362 -12072 47378 -12008
rect 47251 -12088 47378 -12072
rect 47251 -12152 47298 -12088
rect 47362 -12152 47378 -12088
rect 47251 -12168 47378 -12152
rect 47251 -12232 47298 -12168
rect 47362 -12232 47378 -12168
rect 47251 -12248 47378 -12232
rect 47251 -12312 47298 -12248
rect 47362 -12312 47378 -12248
rect 47251 -12328 47378 -12312
rect 47251 -12392 47298 -12328
rect 47362 -12392 47378 -12328
rect 47251 -12408 47378 -12392
rect 47251 -12472 47298 -12408
rect 47362 -12472 47378 -12408
rect 47251 -12488 47378 -12472
rect 47251 -12552 47298 -12488
rect 47362 -12552 47378 -12488
rect 47251 -12568 47378 -12552
rect 47251 -12632 47298 -12568
rect 47362 -12632 47378 -12568
rect 47251 -12648 47378 -12632
rect 47251 -12712 47298 -12648
rect 47362 -12712 47378 -12648
rect 47251 -12728 47378 -12712
rect 47251 -12792 47298 -12728
rect 47362 -12792 47378 -12728
rect 47251 -12808 47378 -12792
rect 47251 -12872 47298 -12808
rect 47362 -12872 47378 -12808
rect 47251 -12888 47378 -12872
rect 47251 -12952 47298 -12888
rect 47362 -12952 47378 -12888
rect 47251 -12968 47378 -12952
rect 47251 -13032 47298 -12968
rect 47362 -13032 47378 -12968
rect 47251 -13048 47378 -13032
rect 47251 -13112 47298 -13048
rect 47362 -13112 47378 -13048
rect 47251 -13128 47378 -13112
rect 47251 -13192 47298 -13128
rect 47362 -13192 47378 -13128
rect 47251 -13208 47378 -13192
rect 47251 -13272 47298 -13208
rect 47362 -13272 47378 -13208
rect 47251 -13288 47378 -13272
rect 47251 -13352 47298 -13288
rect 47362 -13352 47378 -13288
rect 47251 -13368 47378 -13352
rect 47251 -13432 47298 -13368
rect 47362 -13432 47378 -13368
rect 47251 -13448 47378 -13432
rect 47251 -13512 47298 -13448
rect 47362 -13512 47378 -13448
rect 47251 -13528 47378 -13512
rect 47251 -13592 47298 -13528
rect 47362 -13592 47378 -13528
rect 47251 -13608 47378 -13592
rect 47251 -13672 47298 -13608
rect 47362 -13672 47378 -13608
rect 47251 -13688 47378 -13672
rect 47251 -13752 47298 -13688
rect 47362 -13752 47378 -13688
rect 47251 -13768 47378 -13752
rect 47251 -13832 47298 -13768
rect 47362 -13832 47378 -13768
rect 47251 -13848 47378 -13832
rect 47251 -13912 47298 -13848
rect 47362 -13912 47378 -13848
rect 47251 -13928 47378 -13912
rect 47251 -13992 47298 -13928
rect 47362 -13992 47378 -13928
rect 47251 -14008 47378 -13992
rect 47251 -14072 47298 -14008
rect 47362 -14072 47378 -14008
rect 47251 -14088 47378 -14072
rect 47251 -14152 47298 -14088
rect 47362 -14152 47378 -14088
rect 47251 -14168 47378 -14152
rect 47251 -14232 47298 -14168
rect 47362 -14232 47378 -14168
rect 47251 -14248 47378 -14232
rect 47251 -14312 47298 -14248
rect 47362 -14312 47378 -14248
rect 47251 -14328 47378 -14312
rect 47251 -14392 47298 -14328
rect 47362 -14392 47378 -14328
rect 47251 -14408 47378 -14392
rect 47251 -14472 47298 -14408
rect 47362 -14472 47378 -14408
rect 47251 -14488 47378 -14472
rect 47251 -14552 47298 -14488
rect 47362 -14552 47378 -14488
rect 47251 -14568 47378 -14552
rect 47251 -14632 47298 -14568
rect 47362 -14632 47378 -14568
rect 47251 -14648 47378 -14632
rect 47251 -14712 47298 -14648
rect 47362 -14712 47378 -14648
rect 47251 -14728 47378 -14712
rect 47251 -14792 47298 -14728
rect 47362 -14792 47378 -14728
rect 47251 -14808 47378 -14792
rect 47251 -14872 47298 -14808
rect 47362 -14872 47378 -14808
rect 47251 -14888 47378 -14872
rect 47251 -14952 47298 -14888
rect 47362 -14952 47378 -14888
rect 47251 -14968 47378 -14952
rect 47251 -15032 47298 -14968
rect 47362 -15032 47378 -14968
rect 47251 -15048 47378 -15032
rect 47251 -15112 47298 -15048
rect 47362 -15112 47378 -15048
rect 47251 -15128 47378 -15112
rect 47251 -15192 47298 -15128
rect 47362 -15192 47378 -15128
rect 47251 -15208 47378 -15192
rect 47251 -15272 47298 -15208
rect 47362 -15272 47378 -15208
rect 47251 -15288 47378 -15272
rect 47251 -15352 47298 -15288
rect 47362 -15352 47378 -15288
rect 47251 -15368 47378 -15352
rect 47251 -15432 47298 -15368
rect 47362 -15432 47378 -15368
rect 47251 -15448 47378 -15432
rect 47251 -15512 47298 -15448
rect 47362 -15512 47378 -15448
rect 47251 -15528 47378 -15512
rect 40932 -15608 41059 -15592
rect 40932 -15672 40979 -15608
rect 41043 -15672 41059 -15608
rect 40932 -15688 41059 -15672
rect 40932 -15812 41036 -15688
rect 40932 -15828 41059 -15812
rect 40932 -15892 40979 -15828
rect 41043 -15892 41059 -15828
rect 40932 -15908 41059 -15892
rect 34613 -15988 34740 -15972
rect 34613 -16052 34660 -15988
rect 34724 -16052 34740 -15988
rect 34613 -16068 34740 -16052
rect 34613 -16132 34660 -16068
rect 34724 -16132 34740 -16068
rect 34613 -16148 34740 -16132
rect 34613 -16212 34660 -16148
rect 34724 -16212 34740 -16148
rect 34613 -16228 34740 -16212
rect 34613 -16292 34660 -16228
rect 34724 -16292 34740 -16228
rect 34613 -16308 34740 -16292
rect 34613 -16372 34660 -16308
rect 34724 -16372 34740 -16308
rect 34613 -16388 34740 -16372
rect 34613 -16452 34660 -16388
rect 34724 -16452 34740 -16388
rect 34613 -16468 34740 -16452
rect 34613 -16532 34660 -16468
rect 34724 -16532 34740 -16468
rect 34613 -16548 34740 -16532
rect 34613 -16612 34660 -16548
rect 34724 -16612 34740 -16548
rect 34613 -16628 34740 -16612
rect 34613 -16692 34660 -16628
rect 34724 -16692 34740 -16628
rect 34613 -16708 34740 -16692
rect 34613 -16772 34660 -16708
rect 34724 -16772 34740 -16708
rect 34613 -16788 34740 -16772
rect 34613 -16852 34660 -16788
rect 34724 -16852 34740 -16788
rect 34613 -16868 34740 -16852
rect 34613 -16932 34660 -16868
rect 34724 -16932 34740 -16868
rect 34613 -16948 34740 -16932
rect 34613 -17012 34660 -16948
rect 34724 -17012 34740 -16948
rect 34613 -17028 34740 -17012
rect 34613 -17092 34660 -17028
rect 34724 -17092 34740 -17028
rect 34613 -17108 34740 -17092
rect 34613 -17172 34660 -17108
rect 34724 -17172 34740 -17108
rect 34613 -17188 34740 -17172
rect 34613 -17252 34660 -17188
rect 34724 -17252 34740 -17188
rect 34613 -17268 34740 -17252
rect 34613 -17332 34660 -17268
rect 34724 -17332 34740 -17268
rect 34613 -17348 34740 -17332
rect 34613 -17412 34660 -17348
rect 34724 -17412 34740 -17348
rect 34613 -17428 34740 -17412
rect 34613 -17492 34660 -17428
rect 34724 -17492 34740 -17428
rect 34613 -17508 34740 -17492
rect 34613 -17572 34660 -17508
rect 34724 -17572 34740 -17508
rect 34613 -17588 34740 -17572
rect 34613 -17652 34660 -17588
rect 34724 -17652 34740 -17588
rect 34613 -17668 34740 -17652
rect 34613 -17732 34660 -17668
rect 34724 -17732 34740 -17668
rect 34613 -17748 34740 -17732
rect 34613 -17812 34660 -17748
rect 34724 -17812 34740 -17748
rect 34613 -17828 34740 -17812
rect 34613 -17892 34660 -17828
rect 34724 -17892 34740 -17828
rect 34613 -17908 34740 -17892
rect 34613 -17972 34660 -17908
rect 34724 -17972 34740 -17908
rect 34613 -17988 34740 -17972
rect 34613 -18052 34660 -17988
rect 34724 -18052 34740 -17988
rect 34613 -18068 34740 -18052
rect 34613 -18132 34660 -18068
rect 34724 -18132 34740 -18068
rect 34613 -18148 34740 -18132
rect 34613 -18212 34660 -18148
rect 34724 -18212 34740 -18148
rect 34613 -18228 34740 -18212
rect 34613 -18292 34660 -18228
rect 34724 -18292 34740 -18228
rect 34613 -18308 34740 -18292
rect 34613 -18372 34660 -18308
rect 34724 -18372 34740 -18308
rect 34613 -18388 34740 -18372
rect 34613 -18452 34660 -18388
rect 34724 -18452 34740 -18388
rect 34613 -18468 34740 -18452
rect 34613 -18532 34660 -18468
rect 34724 -18532 34740 -18468
rect 34613 -18548 34740 -18532
rect 34613 -18612 34660 -18548
rect 34724 -18612 34740 -18548
rect 34613 -18628 34740 -18612
rect 34613 -18692 34660 -18628
rect 34724 -18692 34740 -18628
rect 34613 -18708 34740 -18692
rect 34613 -18772 34660 -18708
rect 34724 -18772 34740 -18708
rect 34613 -18788 34740 -18772
rect 34613 -18852 34660 -18788
rect 34724 -18852 34740 -18788
rect 34613 -18868 34740 -18852
rect 34613 -18932 34660 -18868
rect 34724 -18932 34740 -18868
rect 34613 -18948 34740 -18932
rect 34613 -19012 34660 -18948
rect 34724 -19012 34740 -18948
rect 34613 -19028 34740 -19012
rect 34613 -19092 34660 -19028
rect 34724 -19092 34740 -19028
rect 34613 -19108 34740 -19092
rect 34613 -19172 34660 -19108
rect 34724 -19172 34740 -19108
rect 34613 -19188 34740 -19172
rect 34613 -19252 34660 -19188
rect 34724 -19252 34740 -19188
rect 34613 -19268 34740 -19252
rect 34613 -19332 34660 -19268
rect 34724 -19332 34740 -19268
rect 34613 -19348 34740 -19332
rect 34613 -19412 34660 -19348
rect 34724 -19412 34740 -19348
rect 34613 -19428 34740 -19412
rect 34613 -19492 34660 -19428
rect 34724 -19492 34740 -19428
rect 34613 -19508 34740 -19492
rect 34613 -19572 34660 -19508
rect 34724 -19572 34740 -19508
rect 34613 -19588 34740 -19572
rect 34613 -19652 34660 -19588
rect 34724 -19652 34740 -19588
rect 34613 -19668 34740 -19652
rect 34613 -19732 34660 -19668
rect 34724 -19732 34740 -19668
rect 34613 -19748 34740 -19732
rect 34613 -19812 34660 -19748
rect 34724 -19812 34740 -19748
rect 34613 -19828 34740 -19812
rect 34613 -19892 34660 -19828
rect 34724 -19892 34740 -19828
rect 34613 -19908 34740 -19892
rect 34613 -19972 34660 -19908
rect 34724 -19972 34740 -19908
rect 34613 -19988 34740 -19972
rect 34613 -20052 34660 -19988
rect 34724 -20052 34740 -19988
rect 34613 -20068 34740 -20052
rect 34613 -20132 34660 -20068
rect 34724 -20132 34740 -20068
rect 34613 -20148 34740 -20132
rect 34613 -20212 34660 -20148
rect 34724 -20212 34740 -20148
rect 34613 -20228 34740 -20212
rect 34613 -20292 34660 -20228
rect 34724 -20292 34740 -20228
rect 34613 -20308 34740 -20292
rect 34613 -20372 34660 -20308
rect 34724 -20372 34740 -20308
rect 34613 -20388 34740 -20372
rect 34613 -20452 34660 -20388
rect 34724 -20452 34740 -20388
rect 34613 -20468 34740 -20452
rect 34613 -20532 34660 -20468
rect 34724 -20532 34740 -20468
rect 34613 -20548 34740 -20532
rect 34613 -20612 34660 -20548
rect 34724 -20612 34740 -20548
rect 34613 -20628 34740 -20612
rect 34613 -20692 34660 -20628
rect 34724 -20692 34740 -20628
rect 34613 -20708 34740 -20692
rect 34613 -20772 34660 -20708
rect 34724 -20772 34740 -20708
rect 34613 -20788 34740 -20772
rect 34613 -20852 34660 -20788
rect 34724 -20852 34740 -20788
rect 34613 -20868 34740 -20852
rect 34613 -20932 34660 -20868
rect 34724 -20932 34740 -20868
rect 34613 -20948 34740 -20932
rect 34613 -21012 34660 -20948
rect 34724 -21012 34740 -20948
rect 34613 -21028 34740 -21012
rect 34613 -21092 34660 -21028
rect 34724 -21092 34740 -21028
rect 34613 -21108 34740 -21092
rect 34613 -21172 34660 -21108
rect 34724 -21172 34740 -21108
rect 34613 -21188 34740 -21172
rect 34613 -21252 34660 -21188
rect 34724 -21252 34740 -21188
rect 34613 -21268 34740 -21252
rect 34613 -21332 34660 -21268
rect 34724 -21332 34740 -21268
rect 34613 -21348 34740 -21332
rect 34613 -21412 34660 -21348
rect 34724 -21412 34740 -21348
rect 34613 -21428 34740 -21412
rect 34613 -21492 34660 -21428
rect 34724 -21492 34740 -21428
rect 34613 -21508 34740 -21492
rect 34613 -21572 34660 -21508
rect 34724 -21572 34740 -21508
rect 34613 -21588 34740 -21572
rect 34613 -21652 34660 -21588
rect 34724 -21652 34740 -21588
rect 34613 -21668 34740 -21652
rect 34613 -21732 34660 -21668
rect 34724 -21732 34740 -21668
rect 34613 -21748 34740 -21732
rect 34613 -21812 34660 -21748
rect 34724 -21812 34740 -21748
rect 34613 -21828 34740 -21812
rect 28294 -21908 28421 -21892
rect 28294 -21972 28341 -21908
rect 28405 -21972 28421 -21908
rect 28294 -21988 28421 -21972
rect 28294 -22112 28398 -21988
rect 28294 -22128 28421 -22112
rect 28294 -22192 28341 -22128
rect 28405 -22192 28421 -22128
rect 28294 -22208 28421 -22192
rect 21975 -22288 22102 -22272
rect 21975 -22352 22022 -22288
rect 22086 -22352 22102 -22288
rect 21975 -22368 22102 -22352
rect 21975 -22432 22022 -22368
rect 22086 -22432 22102 -22368
rect 21975 -22448 22102 -22432
rect 21975 -22512 22022 -22448
rect 22086 -22512 22102 -22448
rect 21975 -22528 22102 -22512
rect 21975 -22592 22022 -22528
rect 22086 -22592 22102 -22528
rect 21975 -22608 22102 -22592
rect 21975 -22672 22022 -22608
rect 22086 -22672 22102 -22608
rect 21975 -22688 22102 -22672
rect 21975 -22752 22022 -22688
rect 22086 -22752 22102 -22688
rect 21975 -22768 22102 -22752
rect 21975 -22832 22022 -22768
rect 22086 -22832 22102 -22768
rect 21975 -22848 22102 -22832
rect 21975 -22912 22022 -22848
rect 22086 -22912 22102 -22848
rect 21975 -22928 22102 -22912
rect 21975 -22992 22022 -22928
rect 22086 -22992 22102 -22928
rect 21975 -23008 22102 -22992
rect 21975 -23072 22022 -23008
rect 22086 -23072 22102 -23008
rect 21975 -23088 22102 -23072
rect 21975 -23152 22022 -23088
rect 22086 -23152 22102 -23088
rect 21975 -23168 22102 -23152
rect 21975 -23232 22022 -23168
rect 22086 -23232 22102 -23168
rect 21975 -23248 22102 -23232
rect 21975 -23312 22022 -23248
rect 22086 -23312 22102 -23248
rect 21975 -23328 22102 -23312
rect 21975 -23392 22022 -23328
rect 22086 -23392 22102 -23328
rect 21975 -23408 22102 -23392
rect 21975 -23472 22022 -23408
rect 22086 -23472 22102 -23408
rect 21975 -23488 22102 -23472
rect 21975 -23552 22022 -23488
rect 22086 -23552 22102 -23488
rect 21975 -23568 22102 -23552
rect 21975 -23632 22022 -23568
rect 22086 -23632 22102 -23568
rect 21975 -23648 22102 -23632
rect 21975 -23712 22022 -23648
rect 22086 -23712 22102 -23648
rect 21975 -23728 22102 -23712
rect 21975 -23792 22022 -23728
rect 22086 -23792 22102 -23728
rect 21975 -23808 22102 -23792
rect 21975 -23872 22022 -23808
rect 22086 -23872 22102 -23808
rect 21975 -23888 22102 -23872
rect 21975 -23952 22022 -23888
rect 22086 -23952 22102 -23888
rect 21975 -23968 22102 -23952
rect 21975 -24032 22022 -23968
rect 22086 -24032 22102 -23968
rect 21975 -24048 22102 -24032
rect 21975 -24112 22022 -24048
rect 22086 -24112 22102 -24048
rect 21975 -24128 22102 -24112
rect 21975 -24192 22022 -24128
rect 22086 -24192 22102 -24128
rect 21975 -24208 22102 -24192
rect 21975 -24272 22022 -24208
rect 22086 -24272 22102 -24208
rect 21975 -24288 22102 -24272
rect 21975 -24352 22022 -24288
rect 22086 -24352 22102 -24288
rect 21975 -24368 22102 -24352
rect 21975 -24432 22022 -24368
rect 22086 -24432 22102 -24368
rect 21975 -24448 22102 -24432
rect 21975 -24512 22022 -24448
rect 22086 -24512 22102 -24448
rect 21975 -24528 22102 -24512
rect 21975 -24592 22022 -24528
rect 22086 -24592 22102 -24528
rect 21975 -24608 22102 -24592
rect 21975 -24672 22022 -24608
rect 22086 -24672 22102 -24608
rect 21975 -24688 22102 -24672
rect 21975 -24752 22022 -24688
rect 22086 -24752 22102 -24688
rect 21975 -24768 22102 -24752
rect 21975 -24832 22022 -24768
rect 22086 -24832 22102 -24768
rect 21975 -24848 22102 -24832
rect 21975 -24912 22022 -24848
rect 22086 -24912 22102 -24848
rect 21975 -24928 22102 -24912
rect 21975 -24992 22022 -24928
rect 22086 -24992 22102 -24928
rect 21975 -25008 22102 -24992
rect 21975 -25072 22022 -25008
rect 22086 -25072 22102 -25008
rect 21975 -25088 22102 -25072
rect 21975 -25152 22022 -25088
rect 22086 -25152 22102 -25088
rect 21975 -25168 22102 -25152
rect 21975 -25232 22022 -25168
rect 22086 -25232 22102 -25168
rect 21975 -25248 22102 -25232
rect 21975 -25312 22022 -25248
rect 22086 -25312 22102 -25248
rect 21975 -25328 22102 -25312
rect 21975 -25392 22022 -25328
rect 22086 -25392 22102 -25328
rect 21975 -25408 22102 -25392
rect 21975 -25472 22022 -25408
rect 22086 -25472 22102 -25408
rect 21975 -25488 22102 -25472
rect 21975 -25552 22022 -25488
rect 22086 -25552 22102 -25488
rect 21975 -25568 22102 -25552
rect 21975 -25632 22022 -25568
rect 22086 -25632 22102 -25568
rect 21975 -25648 22102 -25632
rect 21975 -25712 22022 -25648
rect 22086 -25712 22102 -25648
rect 21975 -25728 22102 -25712
rect 21975 -25792 22022 -25728
rect 22086 -25792 22102 -25728
rect 21975 -25808 22102 -25792
rect 21975 -25872 22022 -25808
rect 22086 -25872 22102 -25808
rect 21975 -25888 22102 -25872
rect 21975 -25952 22022 -25888
rect 22086 -25952 22102 -25888
rect 21975 -25968 22102 -25952
rect 21975 -26032 22022 -25968
rect 22086 -26032 22102 -25968
rect 21975 -26048 22102 -26032
rect 21975 -26112 22022 -26048
rect 22086 -26112 22102 -26048
rect 21975 -26128 22102 -26112
rect 21975 -26192 22022 -26128
rect 22086 -26192 22102 -26128
rect 21975 -26208 22102 -26192
rect 21975 -26272 22022 -26208
rect 22086 -26272 22102 -26208
rect 21975 -26288 22102 -26272
rect 21975 -26352 22022 -26288
rect 22086 -26352 22102 -26288
rect 21975 -26368 22102 -26352
rect 21975 -26432 22022 -26368
rect 22086 -26432 22102 -26368
rect 21975 -26448 22102 -26432
rect 21975 -26512 22022 -26448
rect 22086 -26512 22102 -26448
rect 21975 -26528 22102 -26512
rect 21975 -26592 22022 -26528
rect 22086 -26592 22102 -26528
rect 21975 -26608 22102 -26592
rect 21975 -26672 22022 -26608
rect 22086 -26672 22102 -26608
rect 21975 -26688 22102 -26672
rect 21975 -26752 22022 -26688
rect 22086 -26752 22102 -26688
rect 21975 -26768 22102 -26752
rect 21975 -26832 22022 -26768
rect 22086 -26832 22102 -26768
rect 21975 -26848 22102 -26832
rect 21975 -26912 22022 -26848
rect 22086 -26912 22102 -26848
rect 21975 -26928 22102 -26912
rect 21975 -26992 22022 -26928
rect 22086 -26992 22102 -26928
rect 21975 -27008 22102 -26992
rect 21975 -27072 22022 -27008
rect 22086 -27072 22102 -27008
rect 21975 -27088 22102 -27072
rect 21975 -27152 22022 -27088
rect 22086 -27152 22102 -27088
rect 21975 -27168 22102 -27152
rect 21975 -27232 22022 -27168
rect 22086 -27232 22102 -27168
rect 21975 -27248 22102 -27232
rect 21975 -27312 22022 -27248
rect 22086 -27312 22102 -27248
rect 21975 -27328 22102 -27312
rect 21975 -27392 22022 -27328
rect 22086 -27392 22102 -27328
rect 21975 -27408 22102 -27392
rect 21975 -27472 22022 -27408
rect 22086 -27472 22102 -27408
rect 21975 -27488 22102 -27472
rect 21975 -27552 22022 -27488
rect 22086 -27552 22102 -27488
rect 21975 -27568 22102 -27552
rect 21975 -27632 22022 -27568
rect 22086 -27632 22102 -27568
rect 21975 -27648 22102 -27632
rect 21975 -27712 22022 -27648
rect 22086 -27712 22102 -27648
rect 21975 -27728 22102 -27712
rect 21975 -27792 22022 -27728
rect 22086 -27792 22102 -27728
rect 21975 -27808 22102 -27792
rect 21975 -27872 22022 -27808
rect 22086 -27872 22102 -27808
rect 21975 -27888 22102 -27872
rect 21975 -27952 22022 -27888
rect 22086 -27952 22102 -27888
rect 21975 -27968 22102 -27952
rect 21975 -28032 22022 -27968
rect 22086 -28032 22102 -27968
rect 21975 -28048 22102 -28032
rect 21975 -28112 22022 -28048
rect 22086 -28112 22102 -28048
rect 21975 -28128 22102 -28112
rect 15656 -28208 15783 -28192
rect 15656 -28272 15703 -28208
rect 15767 -28272 15783 -28208
rect 15656 -28288 15783 -28272
rect 15656 -28412 15760 -28288
rect 15656 -28428 15783 -28412
rect 15656 -28492 15703 -28428
rect 15767 -28492 15783 -28428
rect 15656 -28508 15783 -28492
rect 9337 -28588 9464 -28572
rect 9337 -28652 9384 -28588
rect 9448 -28652 9464 -28588
rect 9337 -28668 9464 -28652
rect 9337 -28732 9384 -28668
rect 9448 -28732 9464 -28668
rect 9337 -28748 9464 -28732
rect 9337 -28812 9384 -28748
rect 9448 -28812 9464 -28748
rect 9337 -28828 9464 -28812
rect 9337 -28892 9384 -28828
rect 9448 -28892 9464 -28828
rect 9337 -28908 9464 -28892
rect 9337 -28972 9384 -28908
rect 9448 -28972 9464 -28908
rect 9337 -28988 9464 -28972
rect 9337 -29052 9384 -28988
rect 9448 -29052 9464 -28988
rect 9337 -29068 9464 -29052
rect 9337 -29132 9384 -29068
rect 9448 -29132 9464 -29068
rect 9337 -29148 9464 -29132
rect 9337 -29212 9384 -29148
rect 9448 -29212 9464 -29148
rect 9337 -29228 9464 -29212
rect 9337 -29292 9384 -29228
rect 9448 -29292 9464 -29228
rect 9337 -29308 9464 -29292
rect 9337 -29372 9384 -29308
rect 9448 -29372 9464 -29308
rect 9337 -29388 9464 -29372
rect 9337 -29452 9384 -29388
rect 9448 -29452 9464 -29388
rect 9337 -29468 9464 -29452
rect 9337 -29532 9384 -29468
rect 9448 -29532 9464 -29468
rect 9337 -29548 9464 -29532
rect 9337 -29612 9384 -29548
rect 9448 -29612 9464 -29548
rect 9337 -29628 9464 -29612
rect 9337 -29692 9384 -29628
rect 9448 -29692 9464 -29628
rect 9337 -29708 9464 -29692
rect 9337 -29772 9384 -29708
rect 9448 -29772 9464 -29708
rect 9337 -29788 9464 -29772
rect 9337 -29852 9384 -29788
rect 9448 -29852 9464 -29788
rect 9337 -29868 9464 -29852
rect 9337 -29932 9384 -29868
rect 9448 -29932 9464 -29868
rect 9337 -29948 9464 -29932
rect 9337 -30012 9384 -29948
rect 9448 -30012 9464 -29948
rect 9337 -30028 9464 -30012
rect 9337 -30092 9384 -30028
rect 9448 -30092 9464 -30028
rect 9337 -30108 9464 -30092
rect 9337 -30172 9384 -30108
rect 9448 -30172 9464 -30108
rect 9337 -30188 9464 -30172
rect 9337 -30252 9384 -30188
rect 9448 -30252 9464 -30188
rect 9337 -30268 9464 -30252
rect 9337 -30332 9384 -30268
rect 9448 -30332 9464 -30268
rect 9337 -30348 9464 -30332
rect 9337 -30412 9384 -30348
rect 9448 -30412 9464 -30348
rect 9337 -30428 9464 -30412
rect 9337 -30492 9384 -30428
rect 9448 -30492 9464 -30428
rect 9337 -30508 9464 -30492
rect 9337 -30572 9384 -30508
rect 9448 -30572 9464 -30508
rect 9337 -30588 9464 -30572
rect 9337 -30652 9384 -30588
rect 9448 -30652 9464 -30588
rect 9337 -30668 9464 -30652
rect 9337 -30732 9384 -30668
rect 9448 -30732 9464 -30668
rect 9337 -30748 9464 -30732
rect 9337 -30812 9384 -30748
rect 9448 -30812 9464 -30748
rect 9337 -30828 9464 -30812
rect 9337 -30892 9384 -30828
rect 9448 -30892 9464 -30828
rect 9337 -30908 9464 -30892
rect 9337 -30972 9384 -30908
rect 9448 -30972 9464 -30908
rect 9337 -30988 9464 -30972
rect 9337 -31052 9384 -30988
rect 9448 -31052 9464 -30988
rect 9337 -31068 9464 -31052
rect 9337 -31132 9384 -31068
rect 9448 -31132 9464 -31068
rect 9337 -31148 9464 -31132
rect 9337 -31212 9384 -31148
rect 9448 -31212 9464 -31148
rect 9337 -31228 9464 -31212
rect 9337 -31292 9384 -31228
rect 9448 -31292 9464 -31228
rect 9337 -31308 9464 -31292
rect 9337 -31372 9384 -31308
rect 9448 -31372 9464 -31308
rect 9337 -31388 9464 -31372
rect 9337 -31452 9384 -31388
rect 9448 -31452 9464 -31388
rect 9337 -31468 9464 -31452
rect 9337 -31532 9384 -31468
rect 9448 -31532 9464 -31468
rect 9337 -31548 9464 -31532
rect 9337 -31612 9384 -31548
rect 9448 -31612 9464 -31548
rect 9337 -31628 9464 -31612
rect 9337 -31692 9384 -31628
rect 9448 -31692 9464 -31628
rect 9337 -31708 9464 -31692
rect 9337 -31772 9384 -31708
rect 9448 -31772 9464 -31708
rect 9337 -31788 9464 -31772
rect 9337 -31852 9384 -31788
rect 9448 -31852 9464 -31788
rect 9337 -31868 9464 -31852
rect 9337 -31932 9384 -31868
rect 9448 -31932 9464 -31868
rect 9337 -31948 9464 -31932
rect 9337 -32012 9384 -31948
rect 9448 -32012 9464 -31948
rect 9337 -32028 9464 -32012
rect 9337 -32092 9384 -32028
rect 9448 -32092 9464 -32028
rect 9337 -32108 9464 -32092
rect 9337 -32172 9384 -32108
rect 9448 -32172 9464 -32108
rect 9337 -32188 9464 -32172
rect 9337 -32252 9384 -32188
rect 9448 -32252 9464 -32188
rect 9337 -32268 9464 -32252
rect 9337 -32332 9384 -32268
rect 9448 -32332 9464 -32268
rect 9337 -32348 9464 -32332
rect 9337 -32412 9384 -32348
rect 9448 -32412 9464 -32348
rect 9337 -32428 9464 -32412
rect 9337 -32492 9384 -32428
rect 9448 -32492 9464 -32428
rect 9337 -32508 9464 -32492
rect 9337 -32572 9384 -32508
rect 9448 -32572 9464 -32508
rect 9337 -32588 9464 -32572
rect 9337 -32652 9384 -32588
rect 9448 -32652 9464 -32588
rect 9337 -32668 9464 -32652
rect 9337 -32732 9384 -32668
rect 9448 -32732 9464 -32668
rect 9337 -32748 9464 -32732
rect 9337 -32812 9384 -32748
rect 9448 -32812 9464 -32748
rect 9337 -32828 9464 -32812
rect 9337 -32892 9384 -32828
rect 9448 -32892 9464 -32828
rect 9337 -32908 9464 -32892
rect 9337 -32972 9384 -32908
rect 9448 -32972 9464 -32908
rect 9337 -32988 9464 -32972
rect 9337 -33052 9384 -32988
rect 9448 -33052 9464 -32988
rect 9337 -33068 9464 -33052
rect 9337 -33132 9384 -33068
rect 9448 -33132 9464 -33068
rect 9337 -33148 9464 -33132
rect 9337 -33212 9384 -33148
rect 9448 -33212 9464 -33148
rect 9337 -33228 9464 -33212
rect 9337 -33292 9384 -33228
rect 9448 -33292 9464 -33228
rect 9337 -33308 9464 -33292
rect 9337 -33372 9384 -33308
rect 9448 -33372 9464 -33308
rect 9337 -33388 9464 -33372
rect 9337 -33452 9384 -33388
rect 9448 -33452 9464 -33388
rect 9337 -33468 9464 -33452
rect 9337 -33532 9384 -33468
rect 9448 -33532 9464 -33468
rect 9337 -33548 9464 -33532
rect 9337 -33612 9384 -33548
rect 9448 -33612 9464 -33548
rect 9337 -33628 9464 -33612
rect 9337 -33692 9384 -33628
rect 9448 -33692 9464 -33628
rect 9337 -33708 9464 -33692
rect 9337 -33772 9384 -33708
rect 9448 -33772 9464 -33708
rect 9337 -33788 9464 -33772
rect 9337 -33852 9384 -33788
rect 9448 -33852 9464 -33788
rect 9337 -33868 9464 -33852
rect 9337 -33932 9384 -33868
rect 9448 -33932 9464 -33868
rect 9337 -33948 9464 -33932
rect 9337 -34012 9384 -33948
rect 9448 -34012 9464 -33948
rect 9337 -34028 9464 -34012
rect 9337 -34092 9384 -34028
rect 9448 -34092 9464 -34028
rect 9337 -34108 9464 -34092
rect 9337 -34172 9384 -34108
rect 9448 -34172 9464 -34108
rect 9337 -34188 9464 -34172
rect 9337 -34252 9384 -34188
rect 9448 -34252 9464 -34188
rect 9337 -34268 9464 -34252
rect 9337 -34332 9384 -34268
rect 9448 -34332 9464 -34268
rect 9337 -34348 9464 -34332
rect 9337 -34412 9384 -34348
rect 9448 -34412 9464 -34348
rect 9337 -34428 9464 -34412
rect 3018 -34508 3145 -34492
rect 3018 -34572 3065 -34508
rect 3129 -34572 3145 -34508
rect 3018 -34588 3145 -34572
rect 3018 -34712 3122 -34588
rect 3018 -34728 3145 -34712
rect 3018 -34792 3065 -34728
rect 3129 -34792 3145 -34728
rect 3018 -34808 3145 -34792
rect -3301 -34888 -3174 -34872
rect -3301 -34952 -3254 -34888
rect -3190 -34952 -3174 -34888
rect -3301 -34968 -3174 -34952
rect -3301 -35032 -3254 -34968
rect -3190 -35032 -3174 -34968
rect -3301 -35048 -3174 -35032
rect -3301 -35112 -3254 -35048
rect -3190 -35112 -3174 -35048
rect -3301 -35128 -3174 -35112
rect -3301 -35192 -3254 -35128
rect -3190 -35192 -3174 -35128
rect -3301 -35208 -3174 -35192
rect -3301 -35272 -3254 -35208
rect -3190 -35272 -3174 -35208
rect -3301 -35288 -3174 -35272
rect -3301 -35352 -3254 -35288
rect -3190 -35352 -3174 -35288
rect -3301 -35368 -3174 -35352
rect -3301 -35432 -3254 -35368
rect -3190 -35432 -3174 -35368
rect -3301 -35448 -3174 -35432
rect -3301 -35512 -3254 -35448
rect -3190 -35512 -3174 -35448
rect -3301 -35528 -3174 -35512
rect -3301 -35592 -3254 -35528
rect -3190 -35592 -3174 -35528
rect -3301 -35608 -3174 -35592
rect -3301 -35672 -3254 -35608
rect -3190 -35672 -3174 -35608
rect -3301 -35688 -3174 -35672
rect -3301 -35752 -3254 -35688
rect -3190 -35752 -3174 -35688
rect -3301 -35768 -3174 -35752
rect -3301 -35832 -3254 -35768
rect -3190 -35832 -3174 -35768
rect -3301 -35848 -3174 -35832
rect -3301 -35912 -3254 -35848
rect -3190 -35912 -3174 -35848
rect -3301 -35928 -3174 -35912
rect -3301 -35992 -3254 -35928
rect -3190 -35992 -3174 -35928
rect -3301 -36008 -3174 -35992
rect -3301 -36072 -3254 -36008
rect -3190 -36072 -3174 -36008
rect -3301 -36088 -3174 -36072
rect -3301 -36152 -3254 -36088
rect -3190 -36152 -3174 -36088
rect -3301 -36168 -3174 -36152
rect -3301 -36232 -3254 -36168
rect -3190 -36232 -3174 -36168
rect -3301 -36248 -3174 -36232
rect -3301 -36312 -3254 -36248
rect -3190 -36312 -3174 -36248
rect -3301 -36328 -3174 -36312
rect -3301 -36392 -3254 -36328
rect -3190 -36392 -3174 -36328
rect -3301 -36408 -3174 -36392
rect -3301 -36472 -3254 -36408
rect -3190 -36472 -3174 -36408
rect -3301 -36488 -3174 -36472
rect -3301 -36552 -3254 -36488
rect -3190 -36552 -3174 -36488
rect -3301 -36568 -3174 -36552
rect -3301 -36632 -3254 -36568
rect -3190 -36632 -3174 -36568
rect -3301 -36648 -3174 -36632
rect -3301 -36712 -3254 -36648
rect -3190 -36712 -3174 -36648
rect -3301 -36728 -3174 -36712
rect -3301 -36792 -3254 -36728
rect -3190 -36792 -3174 -36728
rect -3301 -36808 -3174 -36792
rect -3301 -36872 -3254 -36808
rect -3190 -36872 -3174 -36808
rect -3301 -36888 -3174 -36872
rect -3301 -36952 -3254 -36888
rect -3190 -36952 -3174 -36888
rect -3301 -36968 -3174 -36952
rect -3301 -37032 -3254 -36968
rect -3190 -37032 -3174 -36968
rect -3301 -37048 -3174 -37032
rect -3301 -37112 -3254 -37048
rect -3190 -37112 -3174 -37048
rect -3301 -37128 -3174 -37112
rect -3301 -37192 -3254 -37128
rect -3190 -37192 -3174 -37128
rect -3301 -37208 -3174 -37192
rect -3301 -37272 -3254 -37208
rect -3190 -37272 -3174 -37208
rect -3301 -37288 -3174 -37272
rect -3301 -37352 -3254 -37288
rect -3190 -37352 -3174 -37288
rect -3301 -37368 -3174 -37352
rect -3301 -37432 -3254 -37368
rect -3190 -37432 -3174 -37368
rect -3301 -37448 -3174 -37432
rect -3301 -37512 -3254 -37448
rect -3190 -37512 -3174 -37448
rect -3301 -37528 -3174 -37512
rect -3301 -37592 -3254 -37528
rect -3190 -37592 -3174 -37528
rect -3301 -37608 -3174 -37592
rect -3301 -37672 -3254 -37608
rect -3190 -37672 -3174 -37608
rect -3301 -37688 -3174 -37672
rect -3301 -37752 -3254 -37688
rect -3190 -37752 -3174 -37688
rect -3301 -37768 -3174 -37752
rect -3301 -37832 -3254 -37768
rect -3190 -37832 -3174 -37768
rect -3301 -37848 -3174 -37832
rect -3301 -37912 -3254 -37848
rect -3190 -37912 -3174 -37848
rect -3301 -37928 -3174 -37912
rect -3301 -37992 -3254 -37928
rect -3190 -37992 -3174 -37928
rect -3301 -38008 -3174 -37992
rect -3301 -38072 -3254 -38008
rect -3190 -38072 -3174 -38008
rect -3301 -38088 -3174 -38072
rect -3301 -38152 -3254 -38088
rect -3190 -38152 -3174 -38088
rect -3301 -38168 -3174 -38152
rect -3301 -38232 -3254 -38168
rect -3190 -38232 -3174 -38168
rect -3301 -38248 -3174 -38232
rect -3301 -38312 -3254 -38248
rect -3190 -38312 -3174 -38248
rect -3301 -38328 -3174 -38312
rect -3301 -38392 -3254 -38328
rect -3190 -38392 -3174 -38328
rect -3301 -38408 -3174 -38392
rect -3301 -38472 -3254 -38408
rect -3190 -38472 -3174 -38408
rect -3301 -38488 -3174 -38472
rect -3301 -38552 -3254 -38488
rect -3190 -38552 -3174 -38488
rect -3301 -38568 -3174 -38552
rect -3301 -38632 -3254 -38568
rect -3190 -38632 -3174 -38568
rect -3301 -38648 -3174 -38632
rect -3301 -38712 -3254 -38648
rect -3190 -38712 -3174 -38648
rect -3301 -38728 -3174 -38712
rect -3301 -38792 -3254 -38728
rect -3190 -38792 -3174 -38728
rect -3301 -38808 -3174 -38792
rect -3301 -38872 -3254 -38808
rect -3190 -38872 -3174 -38808
rect -3301 -38888 -3174 -38872
rect -3301 -38952 -3254 -38888
rect -3190 -38952 -3174 -38888
rect -3301 -38968 -3174 -38952
rect -3301 -39032 -3254 -38968
rect -3190 -39032 -3174 -38968
rect -3301 -39048 -3174 -39032
rect -3301 -39112 -3254 -39048
rect -3190 -39112 -3174 -39048
rect -3301 -39128 -3174 -39112
rect -3301 -39192 -3254 -39128
rect -3190 -39192 -3174 -39128
rect -3301 -39208 -3174 -39192
rect -3301 -39272 -3254 -39208
rect -3190 -39272 -3174 -39208
rect -3301 -39288 -3174 -39272
rect -3301 -39352 -3254 -39288
rect -3190 -39352 -3174 -39288
rect -3301 -39368 -3174 -39352
rect -3301 -39432 -3254 -39368
rect -3190 -39432 -3174 -39368
rect -3301 -39448 -3174 -39432
rect -3301 -39512 -3254 -39448
rect -3190 -39512 -3174 -39448
rect -3301 -39528 -3174 -39512
rect -3301 -39592 -3254 -39528
rect -3190 -39592 -3174 -39528
rect -3301 -39608 -3174 -39592
rect -3301 -39672 -3254 -39608
rect -3190 -39672 -3174 -39608
rect -3301 -39688 -3174 -39672
rect -3301 -39752 -3254 -39688
rect -3190 -39752 -3174 -39688
rect -3301 -39768 -3174 -39752
rect -3301 -39832 -3254 -39768
rect -3190 -39832 -3174 -39768
rect -3301 -39848 -3174 -39832
rect -3301 -39912 -3254 -39848
rect -3190 -39912 -3174 -39848
rect -3301 -39928 -3174 -39912
rect -3301 -39992 -3254 -39928
rect -3190 -39992 -3174 -39928
rect -3301 -40008 -3174 -39992
rect -3301 -40072 -3254 -40008
rect -3190 -40072 -3174 -40008
rect -3301 -40088 -3174 -40072
rect -3301 -40152 -3254 -40088
rect -3190 -40152 -3174 -40088
rect -3301 -40168 -3174 -40152
rect -3301 -40232 -3254 -40168
rect -3190 -40232 -3174 -40168
rect -3301 -40248 -3174 -40232
rect -3301 -40312 -3254 -40248
rect -3190 -40312 -3174 -40248
rect -3301 -40328 -3174 -40312
rect -3301 -40392 -3254 -40328
rect -3190 -40392 -3174 -40328
rect -3301 -40408 -3174 -40392
rect -3301 -40472 -3254 -40408
rect -3190 -40472 -3174 -40408
rect -3301 -40488 -3174 -40472
rect -3301 -40552 -3254 -40488
rect -3190 -40552 -3174 -40488
rect -3301 -40568 -3174 -40552
rect -3301 -40632 -3254 -40568
rect -3190 -40632 -3174 -40568
rect -3301 -40648 -3174 -40632
rect -3301 -40712 -3254 -40648
rect -3190 -40712 -3174 -40648
rect -3301 -40728 -3174 -40712
rect -9620 -40808 -9493 -40792
rect -9620 -40872 -9573 -40808
rect -9509 -40872 -9493 -40808
rect -9620 -40888 -9493 -40872
rect -9620 -41012 -9516 -40888
rect -9620 -41028 -9493 -41012
rect -9620 -41092 -9573 -41028
rect -9509 -41092 -9493 -41028
rect -9620 -41108 -9493 -41092
rect -15939 -41188 -15812 -41172
rect -15939 -41252 -15892 -41188
rect -15828 -41252 -15812 -41188
rect -15939 -41268 -15812 -41252
rect -15939 -41332 -15892 -41268
rect -15828 -41332 -15812 -41268
rect -15939 -41348 -15812 -41332
rect -15939 -41412 -15892 -41348
rect -15828 -41412 -15812 -41348
rect -15939 -41428 -15812 -41412
rect -15939 -41492 -15892 -41428
rect -15828 -41492 -15812 -41428
rect -15939 -41508 -15812 -41492
rect -15939 -41572 -15892 -41508
rect -15828 -41572 -15812 -41508
rect -15939 -41588 -15812 -41572
rect -15939 -41652 -15892 -41588
rect -15828 -41652 -15812 -41588
rect -15939 -41668 -15812 -41652
rect -15939 -41732 -15892 -41668
rect -15828 -41732 -15812 -41668
rect -15939 -41748 -15812 -41732
rect -15939 -41812 -15892 -41748
rect -15828 -41812 -15812 -41748
rect -15939 -41828 -15812 -41812
rect -15939 -41892 -15892 -41828
rect -15828 -41892 -15812 -41828
rect -15939 -41908 -15812 -41892
rect -15939 -41972 -15892 -41908
rect -15828 -41972 -15812 -41908
rect -15939 -41988 -15812 -41972
rect -15939 -42052 -15892 -41988
rect -15828 -42052 -15812 -41988
rect -15939 -42068 -15812 -42052
rect -15939 -42132 -15892 -42068
rect -15828 -42132 -15812 -42068
rect -15939 -42148 -15812 -42132
rect -15939 -42212 -15892 -42148
rect -15828 -42212 -15812 -42148
rect -15939 -42228 -15812 -42212
rect -15939 -42292 -15892 -42228
rect -15828 -42292 -15812 -42228
rect -15939 -42308 -15812 -42292
rect -15939 -42372 -15892 -42308
rect -15828 -42372 -15812 -42308
rect -15939 -42388 -15812 -42372
rect -15939 -42452 -15892 -42388
rect -15828 -42452 -15812 -42388
rect -15939 -42468 -15812 -42452
rect -15939 -42532 -15892 -42468
rect -15828 -42532 -15812 -42468
rect -15939 -42548 -15812 -42532
rect -15939 -42612 -15892 -42548
rect -15828 -42612 -15812 -42548
rect -15939 -42628 -15812 -42612
rect -15939 -42692 -15892 -42628
rect -15828 -42692 -15812 -42628
rect -15939 -42708 -15812 -42692
rect -15939 -42772 -15892 -42708
rect -15828 -42772 -15812 -42708
rect -15939 -42788 -15812 -42772
rect -15939 -42852 -15892 -42788
rect -15828 -42852 -15812 -42788
rect -15939 -42868 -15812 -42852
rect -15939 -42932 -15892 -42868
rect -15828 -42932 -15812 -42868
rect -15939 -42948 -15812 -42932
rect -15939 -43012 -15892 -42948
rect -15828 -43012 -15812 -42948
rect -15939 -43028 -15812 -43012
rect -15939 -43092 -15892 -43028
rect -15828 -43092 -15812 -43028
rect -15939 -43108 -15812 -43092
rect -15939 -43172 -15892 -43108
rect -15828 -43172 -15812 -43108
rect -15939 -43188 -15812 -43172
rect -15939 -43252 -15892 -43188
rect -15828 -43252 -15812 -43188
rect -15939 -43268 -15812 -43252
rect -15939 -43332 -15892 -43268
rect -15828 -43332 -15812 -43268
rect -15939 -43348 -15812 -43332
rect -15939 -43412 -15892 -43348
rect -15828 -43412 -15812 -43348
rect -15939 -43428 -15812 -43412
rect -15939 -43492 -15892 -43428
rect -15828 -43492 -15812 -43428
rect -15939 -43508 -15812 -43492
rect -15939 -43572 -15892 -43508
rect -15828 -43572 -15812 -43508
rect -15939 -43588 -15812 -43572
rect -15939 -43652 -15892 -43588
rect -15828 -43652 -15812 -43588
rect -15939 -43668 -15812 -43652
rect -15939 -43732 -15892 -43668
rect -15828 -43732 -15812 -43668
rect -15939 -43748 -15812 -43732
rect -15939 -43812 -15892 -43748
rect -15828 -43812 -15812 -43748
rect -15939 -43828 -15812 -43812
rect -15939 -43892 -15892 -43828
rect -15828 -43892 -15812 -43828
rect -15939 -43908 -15812 -43892
rect -15939 -43972 -15892 -43908
rect -15828 -43972 -15812 -43908
rect -15939 -43988 -15812 -43972
rect -15939 -44052 -15892 -43988
rect -15828 -44052 -15812 -43988
rect -15939 -44068 -15812 -44052
rect -15939 -44132 -15892 -44068
rect -15828 -44132 -15812 -44068
rect -15939 -44148 -15812 -44132
rect -15939 -44212 -15892 -44148
rect -15828 -44212 -15812 -44148
rect -15939 -44228 -15812 -44212
rect -15939 -44292 -15892 -44228
rect -15828 -44292 -15812 -44228
rect -15939 -44308 -15812 -44292
rect -15939 -44372 -15892 -44308
rect -15828 -44372 -15812 -44308
rect -15939 -44388 -15812 -44372
rect -15939 -44452 -15892 -44388
rect -15828 -44452 -15812 -44388
rect -15939 -44468 -15812 -44452
rect -15939 -44532 -15892 -44468
rect -15828 -44532 -15812 -44468
rect -15939 -44548 -15812 -44532
rect -15939 -44612 -15892 -44548
rect -15828 -44612 -15812 -44548
rect -15939 -44628 -15812 -44612
rect -15939 -44692 -15892 -44628
rect -15828 -44692 -15812 -44628
rect -15939 -44708 -15812 -44692
rect -15939 -44772 -15892 -44708
rect -15828 -44772 -15812 -44708
rect -15939 -44788 -15812 -44772
rect -15939 -44852 -15892 -44788
rect -15828 -44852 -15812 -44788
rect -15939 -44868 -15812 -44852
rect -15939 -44932 -15892 -44868
rect -15828 -44932 -15812 -44868
rect -15939 -44948 -15812 -44932
rect -15939 -45012 -15892 -44948
rect -15828 -45012 -15812 -44948
rect -15939 -45028 -15812 -45012
rect -15939 -45092 -15892 -45028
rect -15828 -45092 -15812 -45028
rect -15939 -45108 -15812 -45092
rect -15939 -45172 -15892 -45108
rect -15828 -45172 -15812 -45108
rect -15939 -45188 -15812 -45172
rect -15939 -45252 -15892 -45188
rect -15828 -45252 -15812 -45188
rect -15939 -45268 -15812 -45252
rect -15939 -45332 -15892 -45268
rect -15828 -45332 -15812 -45268
rect -15939 -45348 -15812 -45332
rect -15939 -45412 -15892 -45348
rect -15828 -45412 -15812 -45348
rect -15939 -45428 -15812 -45412
rect -15939 -45492 -15892 -45428
rect -15828 -45492 -15812 -45428
rect -15939 -45508 -15812 -45492
rect -15939 -45572 -15892 -45508
rect -15828 -45572 -15812 -45508
rect -15939 -45588 -15812 -45572
rect -15939 -45652 -15892 -45588
rect -15828 -45652 -15812 -45588
rect -15939 -45668 -15812 -45652
rect -15939 -45732 -15892 -45668
rect -15828 -45732 -15812 -45668
rect -15939 -45748 -15812 -45732
rect -15939 -45812 -15892 -45748
rect -15828 -45812 -15812 -45748
rect -15939 -45828 -15812 -45812
rect -15939 -45892 -15892 -45828
rect -15828 -45892 -15812 -45828
rect -15939 -45908 -15812 -45892
rect -15939 -45972 -15892 -45908
rect -15828 -45972 -15812 -45908
rect -15939 -45988 -15812 -45972
rect -15939 -46052 -15892 -45988
rect -15828 -46052 -15812 -45988
rect -15939 -46068 -15812 -46052
rect -15939 -46132 -15892 -46068
rect -15828 -46132 -15812 -46068
rect -15939 -46148 -15812 -46132
rect -15939 -46212 -15892 -46148
rect -15828 -46212 -15812 -46148
rect -15939 -46228 -15812 -46212
rect -15939 -46292 -15892 -46228
rect -15828 -46292 -15812 -46228
rect -15939 -46308 -15812 -46292
rect -15939 -46372 -15892 -46308
rect -15828 -46372 -15812 -46308
rect -15939 -46388 -15812 -46372
rect -15939 -46452 -15892 -46388
rect -15828 -46452 -15812 -46388
rect -15939 -46468 -15812 -46452
rect -15939 -46532 -15892 -46468
rect -15828 -46532 -15812 -46468
rect -15939 -46548 -15812 -46532
rect -15939 -46612 -15892 -46548
rect -15828 -46612 -15812 -46548
rect -15939 -46628 -15812 -46612
rect -15939 -46692 -15892 -46628
rect -15828 -46692 -15812 -46628
rect -15939 -46708 -15812 -46692
rect -15939 -46772 -15892 -46708
rect -15828 -46772 -15812 -46708
rect -15939 -46788 -15812 -46772
rect -15939 -46852 -15892 -46788
rect -15828 -46852 -15812 -46788
rect -15939 -46868 -15812 -46852
rect -15939 -46932 -15892 -46868
rect -15828 -46932 -15812 -46868
rect -15939 -46948 -15812 -46932
rect -15939 -47012 -15892 -46948
rect -15828 -47012 -15812 -46948
rect -15939 -47028 -15812 -47012
rect -22258 -47108 -22131 -47092
rect -22258 -47172 -22211 -47108
rect -22147 -47172 -22131 -47108
rect -22258 -47188 -22131 -47172
rect -22258 -47250 -22154 -47188
rect -19059 -47250 -18955 -47061
rect -15939 -47092 -15892 -47028
rect -15828 -47092 -15812 -47028
rect -15649 -41148 -9727 -41139
rect -15649 -47052 -15640 -41148
rect -9736 -47052 -9727 -41148
rect -15649 -47061 -9727 -47052
rect -9620 -41172 -9573 -41108
rect -9509 -41172 -9493 -41108
rect -6421 -41139 -6317 -40761
rect -3301 -40792 -3254 -40728
rect -3190 -40792 -3174 -40728
rect -3011 -34848 2911 -34839
rect -3011 -40752 -3002 -34848
rect 2902 -40752 2911 -34848
rect -3011 -40761 2911 -40752
rect 3018 -34872 3065 -34808
rect 3129 -34872 3145 -34808
rect 6217 -34839 6321 -34461
rect 9337 -34492 9384 -34428
rect 9448 -34492 9464 -34428
rect 9627 -28548 15549 -28539
rect 9627 -34452 9636 -28548
rect 15540 -34452 15549 -28548
rect 9627 -34461 15549 -34452
rect 15656 -28572 15703 -28508
rect 15767 -28572 15783 -28508
rect 18855 -28539 18959 -28161
rect 21975 -28192 22022 -28128
rect 22086 -28192 22102 -28128
rect 22265 -22248 28187 -22239
rect 22265 -28152 22274 -22248
rect 28178 -28152 28187 -22248
rect 22265 -28161 28187 -28152
rect 28294 -22272 28341 -22208
rect 28405 -22272 28421 -22208
rect 31493 -22239 31597 -21861
rect 34613 -21892 34660 -21828
rect 34724 -21892 34740 -21828
rect 34903 -15948 40825 -15939
rect 34903 -21852 34912 -15948
rect 40816 -21852 40825 -15948
rect 34903 -21861 40825 -21852
rect 40932 -15972 40979 -15908
rect 41043 -15972 41059 -15908
rect 44131 -15939 44235 -15561
rect 47251 -15592 47298 -15528
rect 47362 -15592 47378 -15528
rect 47251 -15608 47378 -15592
rect 47251 -15672 47298 -15608
rect 47362 -15672 47378 -15608
rect 47251 -15688 47378 -15672
rect 47251 -15812 47355 -15688
rect 47251 -15828 47378 -15812
rect 47251 -15892 47298 -15828
rect 47362 -15892 47378 -15828
rect 47251 -15908 47378 -15892
rect 40932 -15988 41059 -15972
rect 40932 -16052 40979 -15988
rect 41043 -16052 41059 -15988
rect 40932 -16068 41059 -16052
rect 40932 -16132 40979 -16068
rect 41043 -16132 41059 -16068
rect 40932 -16148 41059 -16132
rect 40932 -16212 40979 -16148
rect 41043 -16212 41059 -16148
rect 40932 -16228 41059 -16212
rect 40932 -16292 40979 -16228
rect 41043 -16292 41059 -16228
rect 40932 -16308 41059 -16292
rect 40932 -16372 40979 -16308
rect 41043 -16372 41059 -16308
rect 40932 -16388 41059 -16372
rect 40932 -16452 40979 -16388
rect 41043 -16452 41059 -16388
rect 40932 -16468 41059 -16452
rect 40932 -16532 40979 -16468
rect 41043 -16532 41059 -16468
rect 40932 -16548 41059 -16532
rect 40932 -16612 40979 -16548
rect 41043 -16612 41059 -16548
rect 40932 -16628 41059 -16612
rect 40932 -16692 40979 -16628
rect 41043 -16692 41059 -16628
rect 40932 -16708 41059 -16692
rect 40932 -16772 40979 -16708
rect 41043 -16772 41059 -16708
rect 40932 -16788 41059 -16772
rect 40932 -16852 40979 -16788
rect 41043 -16852 41059 -16788
rect 40932 -16868 41059 -16852
rect 40932 -16932 40979 -16868
rect 41043 -16932 41059 -16868
rect 40932 -16948 41059 -16932
rect 40932 -17012 40979 -16948
rect 41043 -17012 41059 -16948
rect 40932 -17028 41059 -17012
rect 40932 -17092 40979 -17028
rect 41043 -17092 41059 -17028
rect 40932 -17108 41059 -17092
rect 40932 -17172 40979 -17108
rect 41043 -17172 41059 -17108
rect 40932 -17188 41059 -17172
rect 40932 -17252 40979 -17188
rect 41043 -17252 41059 -17188
rect 40932 -17268 41059 -17252
rect 40932 -17332 40979 -17268
rect 41043 -17332 41059 -17268
rect 40932 -17348 41059 -17332
rect 40932 -17412 40979 -17348
rect 41043 -17412 41059 -17348
rect 40932 -17428 41059 -17412
rect 40932 -17492 40979 -17428
rect 41043 -17492 41059 -17428
rect 40932 -17508 41059 -17492
rect 40932 -17572 40979 -17508
rect 41043 -17572 41059 -17508
rect 40932 -17588 41059 -17572
rect 40932 -17652 40979 -17588
rect 41043 -17652 41059 -17588
rect 40932 -17668 41059 -17652
rect 40932 -17732 40979 -17668
rect 41043 -17732 41059 -17668
rect 40932 -17748 41059 -17732
rect 40932 -17812 40979 -17748
rect 41043 -17812 41059 -17748
rect 40932 -17828 41059 -17812
rect 40932 -17892 40979 -17828
rect 41043 -17892 41059 -17828
rect 40932 -17908 41059 -17892
rect 40932 -17972 40979 -17908
rect 41043 -17972 41059 -17908
rect 40932 -17988 41059 -17972
rect 40932 -18052 40979 -17988
rect 41043 -18052 41059 -17988
rect 40932 -18068 41059 -18052
rect 40932 -18132 40979 -18068
rect 41043 -18132 41059 -18068
rect 40932 -18148 41059 -18132
rect 40932 -18212 40979 -18148
rect 41043 -18212 41059 -18148
rect 40932 -18228 41059 -18212
rect 40932 -18292 40979 -18228
rect 41043 -18292 41059 -18228
rect 40932 -18308 41059 -18292
rect 40932 -18372 40979 -18308
rect 41043 -18372 41059 -18308
rect 40932 -18388 41059 -18372
rect 40932 -18452 40979 -18388
rect 41043 -18452 41059 -18388
rect 40932 -18468 41059 -18452
rect 40932 -18532 40979 -18468
rect 41043 -18532 41059 -18468
rect 40932 -18548 41059 -18532
rect 40932 -18612 40979 -18548
rect 41043 -18612 41059 -18548
rect 40932 -18628 41059 -18612
rect 40932 -18692 40979 -18628
rect 41043 -18692 41059 -18628
rect 40932 -18708 41059 -18692
rect 40932 -18772 40979 -18708
rect 41043 -18772 41059 -18708
rect 40932 -18788 41059 -18772
rect 40932 -18852 40979 -18788
rect 41043 -18852 41059 -18788
rect 40932 -18868 41059 -18852
rect 40932 -18932 40979 -18868
rect 41043 -18932 41059 -18868
rect 40932 -18948 41059 -18932
rect 40932 -19012 40979 -18948
rect 41043 -19012 41059 -18948
rect 40932 -19028 41059 -19012
rect 40932 -19092 40979 -19028
rect 41043 -19092 41059 -19028
rect 40932 -19108 41059 -19092
rect 40932 -19172 40979 -19108
rect 41043 -19172 41059 -19108
rect 40932 -19188 41059 -19172
rect 40932 -19252 40979 -19188
rect 41043 -19252 41059 -19188
rect 40932 -19268 41059 -19252
rect 40932 -19332 40979 -19268
rect 41043 -19332 41059 -19268
rect 40932 -19348 41059 -19332
rect 40932 -19412 40979 -19348
rect 41043 -19412 41059 -19348
rect 40932 -19428 41059 -19412
rect 40932 -19492 40979 -19428
rect 41043 -19492 41059 -19428
rect 40932 -19508 41059 -19492
rect 40932 -19572 40979 -19508
rect 41043 -19572 41059 -19508
rect 40932 -19588 41059 -19572
rect 40932 -19652 40979 -19588
rect 41043 -19652 41059 -19588
rect 40932 -19668 41059 -19652
rect 40932 -19732 40979 -19668
rect 41043 -19732 41059 -19668
rect 40932 -19748 41059 -19732
rect 40932 -19812 40979 -19748
rect 41043 -19812 41059 -19748
rect 40932 -19828 41059 -19812
rect 40932 -19892 40979 -19828
rect 41043 -19892 41059 -19828
rect 40932 -19908 41059 -19892
rect 40932 -19972 40979 -19908
rect 41043 -19972 41059 -19908
rect 40932 -19988 41059 -19972
rect 40932 -20052 40979 -19988
rect 41043 -20052 41059 -19988
rect 40932 -20068 41059 -20052
rect 40932 -20132 40979 -20068
rect 41043 -20132 41059 -20068
rect 40932 -20148 41059 -20132
rect 40932 -20212 40979 -20148
rect 41043 -20212 41059 -20148
rect 40932 -20228 41059 -20212
rect 40932 -20292 40979 -20228
rect 41043 -20292 41059 -20228
rect 40932 -20308 41059 -20292
rect 40932 -20372 40979 -20308
rect 41043 -20372 41059 -20308
rect 40932 -20388 41059 -20372
rect 40932 -20452 40979 -20388
rect 41043 -20452 41059 -20388
rect 40932 -20468 41059 -20452
rect 40932 -20532 40979 -20468
rect 41043 -20532 41059 -20468
rect 40932 -20548 41059 -20532
rect 40932 -20612 40979 -20548
rect 41043 -20612 41059 -20548
rect 40932 -20628 41059 -20612
rect 40932 -20692 40979 -20628
rect 41043 -20692 41059 -20628
rect 40932 -20708 41059 -20692
rect 40932 -20772 40979 -20708
rect 41043 -20772 41059 -20708
rect 40932 -20788 41059 -20772
rect 40932 -20852 40979 -20788
rect 41043 -20852 41059 -20788
rect 40932 -20868 41059 -20852
rect 40932 -20932 40979 -20868
rect 41043 -20932 41059 -20868
rect 40932 -20948 41059 -20932
rect 40932 -21012 40979 -20948
rect 41043 -21012 41059 -20948
rect 40932 -21028 41059 -21012
rect 40932 -21092 40979 -21028
rect 41043 -21092 41059 -21028
rect 40932 -21108 41059 -21092
rect 40932 -21172 40979 -21108
rect 41043 -21172 41059 -21108
rect 40932 -21188 41059 -21172
rect 40932 -21252 40979 -21188
rect 41043 -21252 41059 -21188
rect 40932 -21268 41059 -21252
rect 40932 -21332 40979 -21268
rect 41043 -21332 41059 -21268
rect 40932 -21348 41059 -21332
rect 40932 -21412 40979 -21348
rect 41043 -21412 41059 -21348
rect 40932 -21428 41059 -21412
rect 40932 -21492 40979 -21428
rect 41043 -21492 41059 -21428
rect 40932 -21508 41059 -21492
rect 40932 -21572 40979 -21508
rect 41043 -21572 41059 -21508
rect 40932 -21588 41059 -21572
rect 40932 -21652 40979 -21588
rect 41043 -21652 41059 -21588
rect 40932 -21668 41059 -21652
rect 40932 -21732 40979 -21668
rect 41043 -21732 41059 -21668
rect 40932 -21748 41059 -21732
rect 40932 -21812 40979 -21748
rect 41043 -21812 41059 -21748
rect 40932 -21828 41059 -21812
rect 34613 -21908 34740 -21892
rect 34613 -21972 34660 -21908
rect 34724 -21972 34740 -21908
rect 34613 -21988 34740 -21972
rect 34613 -22112 34717 -21988
rect 34613 -22128 34740 -22112
rect 34613 -22192 34660 -22128
rect 34724 -22192 34740 -22128
rect 34613 -22208 34740 -22192
rect 28294 -22288 28421 -22272
rect 28294 -22352 28341 -22288
rect 28405 -22352 28421 -22288
rect 28294 -22368 28421 -22352
rect 28294 -22432 28341 -22368
rect 28405 -22432 28421 -22368
rect 28294 -22448 28421 -22432
rect 28294 -22512 28341 -22448
rect 28405 -22512 28421 -22448
rect 28294 -22528 28421 -22512
rect 28294 -22592 28341 -22528
rect 28405 -22592 28421 -22528
rect 28294 -22608 28421 -22592
rect 28294 -22672 28341 -22608
rect 28405 -22672 28421 -22608
rect 28294 -22688 28421 -22672
rect 28294 -22752 28341 -22688
rect 28405 -22752 28421 -22688
rect 28294 -22768 28421 -22752
rect 28294 -22832 28341 -22768
rect 28405 -22832 28421 -22768
rect 28294 -22848 28421 -22832
rect 28294 -22912 28341 -22848
rect 28405 -22912 28421 -22848
rect 28294 -22928 28421 -22912
rect 28294 -22992 28341 -22928
rect 28405 -22992 28421 -22928
rect 28294 -23008 28421 -22992
rect 28294 -23072 28341 -23008
rect 28405 -23072 28421 -23008
rect 28294 -23088 28421 -23072
rect 28294 -23152 28341 -23088
rect 28405 -23152 28421 -23088
rect 28294 -23168 28421 -23152
rect 28294 -23232 28341 -23168
rect 28405 -23232 28421 -23168
rect 28294 -23248 28421 -23232
rect 28294 -23312 28341 -23248
rect 28405 -23312 28421 -23248
rect 28294 -23328 28421 -23312
rect 28294 -23392 28341 -23328
rect 28405 -23392 28421 -23328
rect 28294 -23408 28421 -23392
rect 28294 -23472 28341 -23408
rect 28405 -23472 28421 -23408
rect 28294 -23488 28421 -23472
rect 28294 -23552 28341 -23488
rect 28405 -23552 28421 -23488
rect 28294 -23568 28421 -23552
rect 28294 -23632 28341 -23568
rect 28405 -23632 28421 -23568
rect 28294 -23648 28421 -23632
rect 28294 -23712 28341 -23648
rect 28405 -23712 28421 -23648
rect 28294 -23728 28421 -23712
rect 28294 -23792 28341 -23728
rect 28405 -23792 28421 -23728
rect 28294 -23808 28421 -23792
rect 28294 -23872 28341 -23808
rect 28405 -23872 28421 -23808
rect 28294 -23888 28421 -23872
rect 28294 -23952 28341 -23888
rect 28405 -23952 28421 -23888
rect 28294 -23968 28421 -23952
rect 28294 -24032 28341 -23968
rect 28405 -24032 28421 -23968
rect 28294 -24048 28421 -24032
rect 28294 -24112 28341 -24048
rect 28405 -24112 28421 -24048
rect 28294 -24128 28421 -24112
rect 28294 -24192 28341 -24128
rect 28405 -24192 28421 -24128
rect 28294 -24208 28421 -24192
rect 28294 -24272 28341 -24208
rect 28405 -24272 28421 -24208
rect 28294 -24288 28421 -24272
rect 28294 -24352 28341 -24288
rect 28405 -24352 28421 -24288
rect 28294 -24368 28421 -24352
rect 28294 -24432 28341 -24368
rect 28405 -24432 28421 -24368
rect 28294 -24448 28421 -24432
rect 28294 -24512 28341 -24448
rect 28405 -24512 28421 -24448
rect 28294 -24528 28421 -24512
rect 28294 -24592 28341 -24528
rect 28405 -24592 28421 -24528
rect 28294 -24608 28421 -24592
rect 28294 -24672 28341 -24608
rect 28405 -24672 28421 -24608
rect 28294 -24688 28421 -24672
rect 28294 -24752 28341 -24688
rect 28405 -24752 28421 -24688
rect 28294 -24768 28421 -24752
rect 28294 -24832 28341 -24768
rect 28405 -24832 28421 -24768
rect 28294 -24848 28421 -24832
rect 28294 -24912 28341 -24848
rect 28405 -24912 28421 -24848
rect 28294 -24928 28421 -24912
rect 28294 -24992 28341 -24928
rect 28405 -24992 28421 -24928
rect 28294 -25008 28421 -24992
rect 28294 -25072 28341 -25008
rect 28405 -25072 28421 -25008
rect 28294 -25088 28421 -25072
rect 28294 -25152 28341 -25088
rect 28405 -25152 28421 -25088
rect 28294 -25168 28421 -25152
rect 28294 -25232 28341 -25168
rect 28405 -25232 28421 -25168
rect 28294 -25248 28421 -25232
rect 28294 -25312 28341 -25248
rect 28405 -25312 28421 -25248
rect 28294 -25328 28421 -25312
rect 28294 -25392 28341 -25328
rect 28405 -25392 28421 -25328
rect 28294 -25408 28421 -25392
rect 28294 -25472 28341 -25408
rect 28405 -25472 28421 -25408
rect 28294 -25488 28421 -25472
rect 28294 -25552 28341 -25488
rect 28405 -25552 28421 -25488
rect 28294 -25568 28421 -25552
rect 28294 -25632 28341 -25568
rect 28405 -25632 28421 -25568
rect 28294 -25648 28421 -25632
rect 28294 -25712 28341 -25648
rect 28405 -25712 28421 -25648
rect 28294 -25728 28421 -25712
rect 28294 -25792 28341 -25728
rect 28405 -25792 28421 -25728
rect 28294 -25808 28421 -25792
rect 28294 -25872 28341 -25808
rect 28405 -25872 28421 -25808
rect 28294 -25888 28421 -25872
rect 28294 -25952 28341 -25888
rect 28405 -25952 28421 -25888
rect 28294 -25968 28421 -25952
rect 28294 -26032 28341 -25968
rect 28405 -26032 28421 -25968
rect 28294 -26048 28421 -26032
rect 28294 -26112 28341 -26048
rect 28405 -26112 28421 -26048
rect 28294 -26128 28421 -26112
rect 28294 -26192 28341 -26128
rect 28405 -26192 28421 -26128
rect 28294 -26208 28421 -26192
rect 28294 -26272 28341 -26208
rect 28405 -26272 28421 -26208
rect 28294 -26288 28421 -26272
rect 28294 -26352 28341 -26288
rect 28405 -26352 28421 -26288
rect 28294 -26368 28421 -26352
rect 28294 -26432 28341 -26368
rect 28405 -26432 28421 -26368
rect 28294 -26448 28421 -26432
rect 28294 -26512 28341 -26448
rect 28405 -26512 28421 -26448
rect 28294 -26528 28421 -26512
rect 28294 -26592 28341 -26528
rect 28405 -26592 28421 -26528
rect 28294 -26608 28421 -26592
rect 28294 -26672 28341 -26608
rect 28405 -26672 28421 -26608
rect 28294 -26688 28421 -26672
rect 28294 -26752 28341 -26688
rect 28405 -26752 28421 -26688
rect 28294 -26768 28421 -26752
rect 28294 -26832 28341 -26768
rect 28405 -26832 28421 -26768
rect 28294 -26848 28421 -26832
rect 28294 -26912 28341 -26848
rect 28405 -26912 28421 -26848
rect 28294 -26928 28421 -26912
rect 28294 -26992 28341 -26928
rect 28405 -26992 28421 -26928
rect 28294 -27008 28421 -26992
rect 28294 -27072 28341 -27008
rect 28405 -27072 28421 -27008
rect 28294 -27088 28421 -27072
rect 28294 -27152 28341 -27088
rect 28405 -27152 28421 -27088
rect 28294 -27168 28421 -27152
rect 28294 -27232 28341 -27168
rect 28405 -27232 28421 -27168
rect 28294 -27248 28421 -27232
rect 28294 -27312 28341 -27248
rect 28405 -27312 28421 -27248
rect 28294 -27328 28421 -27312
rect 28294 -27392 28341 -27328
rect 28405 -27392 28421 -27328
rect 28294 -27408 28421 -27392
rect 28294 -27472 28341 -27408
rect 28405 -27472 28421 -27408
rect 28294 -27488 28421 -27472
rect 28294 -27552 28341 -27488
rect 28405 -27552 28421 -27488
rect 28294 -27568 28421 -27552
rect 28294 -27632 28341 -27568
rect 28405 -27632 28421 -27568
rect 28294 -27648 28421 -27632
rect 28294 -27712 28341 -27648
rect 28405 -27712 28421 -27648
rect 28294 -27728 28421 -27712
rect 28294 -27792 28341 -27728
rect 28405 -27792 28421 -27728
rect 28294 -27808 28421 -27792
rect 28294 -27872 28341 -27808
rect 28405 -27872 28421 -27808
rect 28294 -27888 28421 -27872
rect 28294 -27952 28341 -27888
rect 28405 -27952 28421 -27888
rect 28294 -27968 28421 -27952
rect 28294 -28032 28341 -27968
rect 28405 -28032 28421 -27968
rect 28294 -28048 28421 -28032
rect 28294 -28112 28341 -28048
rect 28405 -28112 28421 -28048
rect 28294 -28128 28421 -28112
rect 21975 -28208 22102 -28192
rect 21975 -28272 22022 -28208
rect 22086 -28272 22102 -28208
rect 21975 -28288 22102 -28272
rect 21975 -28412 22079 -28288
rect 21975 -28428 22102 -28412
rect 21975 -28492 22022 -28428
rect 22086 -28492 22102 -28428
rect 21975 -28508 22102 -28492
rect 15656 -28588 15783 -28572
rect 15656 -28652 15703 -28588
rect 15767 -28652 15783 -28588
rect 15656 -28668 15783 -28652
rect 15656 -28732 15703 -28668
rect 15767 -28732 15783 -28668
rect 15656 -28748 15783 -28732
rect 15656 -28812 15703 -28748
rect 15767 -28812 15783 -28748
rect 15656 -28828 15783 -28812
rect 15656 -28892 15703 -28828
rect 15767 -28892 15783 -28828
rect 15656 -28908 15783 -28892
rect 15656 -28972 15703 -28908
rect 15767 -28972 15783 -28908
rect 15656 -28988 15783 -28972
rect 15656 -29052 15703 -28988
rect 15767 -29052 15783 -28988
rect 15656 -29068 15783 -29052
rect 15656 -29132 15703 -29068
rect 15767 -29132 15783 -29068
rect 15656 -29148 15783 -29132
rect 15656 -29212 15703 -29148
rect 15767 -29212 15783 -29148
rect 15656 -29228 15783 -29212
rect 15656 -29292 15703 -29228
rect 15767 -29292 15783 -29228
rect 15656 -29308 15783 -29292
rect 15656 -29372 15703 -29308
rect 15767 -29372 15783 -29308
rect 15656 -29388 15783 -29372
rect 15656 -29452 15703 -29388
rect 15767 -29452 15783 -29388
rect 15656 -29468 15783 -29452
rect 15656 -29532 15703 -29468
rect 15767 -29532 15783 -29468
rect 15656 -29548 15783 -29532
rect 15656 -29612 15703 -29548
rect 15767 -29612 15783 -29548
rect 15656 -29628 15783 -29612
rect 15656 -29692 15703 -29628
rect 15767 -29692 15783 -29628
rect 15656 -29708 15783 -29692
rect 15656 -29772 15703 -29708
rect 15767 -29772 15783 -29708
rect 15656 -29788 15783 -29772
rect 15656 -29852 15703 -29788
rect 15767 -29852 15783 -29788
rect 15656 -29868 15783 -29852
rect 15656 -29932 15703 -29868
rect 15767 -29932 15783 -29868
rect 15656 -29948 15783 -29932
rect 15656 -30012 15703 -29948
rect 15767 -30012 15783 -29948
rect 15656 -30028 15783 -30012
rect 15656 -30092 15703 -30028
rect 15767 -30092 15783 -30028
rect 15656 -30108 15783 -30092
rect 15656 -30172 15703 -30108
rect 15767 -30172 15783 -30108
rect 15656 -30188 15783 -30172
rect 15656 -30252 15703 -30188
rect 15767 -30252 15783 -30188
rect 15656 -30268 15783 -30252
rect 15656 -30332 15703 -30268
rect 15767 -30332 15783 -30268
rect 15656 -30348 15783 -30332
rect 15656 -30412 15703 -30348
rect 15767 -30412 15783 -30348
rect 15656 -30428 15783 -30412
rect 15656 -30492 15703 -30428
rect 15767 -30492 15783 -30428
rect 15656 -30508 15783 -30492
rect 15656 -30572 15703 -30508
rect 15767 -30572 15783 -30508
rect 15656 -30588 15783 -30572
rect 15656 -30652 15703 -30588
rect 15767 -30652 15783 -30588
rect 15656 -30668 15783 -30652
rect 15656 -30732 15703 -30668
rect 15767 -30732 15783 -30668
rect 15656 -30748 15783 -30732
rect 15656 -30812 15703 -30748
rect 15767 -30812 15783 -30748
rect 15656 -30828 15783 -30812
rect 15656 -30892 15703 -30828
rect 15767 -30892 15783 -30828
rect 15656 -30908 15783 -30892
rect 15656 -30972 15703 -30908
rect 15767 -30972 15783 -30908
rect 15656 -30988 15783 -30972
rect 15656 -31052 15703 -30988
rect 15767 -31052 15783 -30988
rect 15656 -31068 15783 -31052
rect 15656 -31132 15703 -31068
rect 15767 -31132 15783 -31068
rect 15656 -31148 15783 -31132
rect 15656 -31212 15703 -31148
rect 15767 -31212 15783 -31148
rect 15656 -31228 15783 -31212
rect 15656 -31292 15703 -31228
rect 15767 -31292 15783 -31228
rect 15656 -31308 15783 -31292
rect 15656 -31372 15703 -31308
rect 15767 -31372 15783 -31308
rect 15656 -31388 15783 -31372
rect 15656 -31452 15703 -31388
rect 15767 -31452 15783 -31388
rect 15656 -31468 15783 -31452
rect 15656 -31532 15703 -31468
rect 15767 -31532 15783 -31468
rect 15656 -31548 15783 -31532
rect 15656 -31612 15703 -31548
rect 15767 -31612 15783 -31548
rect 15656 -31628 15783 -31612
rect 15656 -31692 15703 -31628
rect 15767 -31692 15783 -31628
rect 15656 -31708 15783 -31692
rect 15656 -31772 15703 -31708
rect 15767 -31772 15783 -31708
rect 15656 -31788 15783 -31772
rect 15656 -31852 15703 -31788
rect 15767 -31852 15783 -31788
rect 15656 -31868 15783 -31852
rect 15656 -31932 15703 -31868
rect 15767 -31932 15783 -31868
rect 15656 -31948 15783 -31932
rect 15656 -32012 15703 -31948
rect 15767 -32012 15783 -31948
rect 15656 -32028 15783 -32012
rect 15656 -32092 15703 -32028
rect 15767 -32092 15783 -32028
rect 15656 -32108 15783 -32092
rect 15656 -32172 15703 -32108
rect 15767 -32172 15783 -32108
rect 15656 -32188 15783 -32172
rect 15656 -32252 15703 -32188
rect 15767 -32252 15783 -32188
rect 15656 -32268 15783 -32252
rect 15656 -32332 15703 -32268
rect 15767 -32332 15783 -32268
rect 15656 -32348 15783 -32332
rect 15656 -32412 15703 -32348
rect 15767 -32412 15783 -32348
rect 15656 -32428 15783 -32412
rect 15656 -32492 15703 -32428
rect 15767 -32492 15783 -32428
rect 15656 -32508 15783 -32492
rect 15656 -32572 15703 -32508
rect 15767 -32572 15783 -32508
rect 15656 -32588 15783 -32572
rect 15656 -32652 15703 -32588
rect 15767 -32652 15783 -32588
rect 15656 -32668 15783 -32652
rect 15656 -32732 15703 -32668
rect 15767 -32732 15783 -32668
rect 15656 -32748 15783 -32732
rect 15656 -32812 15703 -32748
rect 15767 -32812 15783 -32748
rect 15656 -32828 15783 -32812
rect 15656 -32892 15703 -32828
rect 15767 -32892 15783 -32828
rect 15656 -32908 15783 -32892
rect 15656 -32972 15703 -32908
rect 15767 -32972 15783 -32908
rect 15656 -32988 15783 -32972
rect 15656 -33052 15703 -32988
rect 15767 -33052 15783 -32988
rect 15656 -33068 15783 -33052
rect 15656 -33132 15703 -33068
rect 15767 -33132 15783 -33068
rect 15656 -33148 15783 -33132
rect 15656 -33212 15703 -33148
rect 15767 -33212 15783 -33148
rect 15656 -33228 15783 -33212
rect 15656 -33292 15703 -33228
rect 15767 -33292 15783 -33228
rect 15656 -33308 15783 -33292
rect 15656 -33372 15703 -33308
rect 15767 -33372 15783 -33308
rect 15656 -33388 15783 -33372
rect 15656 -33452 15703 -33388
rect 15767 -33452 15783 -33388
rect 15656 -33468 15783 -33452
rect 15656 -33532 15703 -33468
rect 15767 -33532 15783 -33468
rect 15656 -33548 15783 -33532
rect 15656 -33612 15703 -33548
rect 15767 -33612 15783 -33548
rect 15656 -33628 15783 -33612
rect 15656 -33692 15703 -33628
rect 15767 -33692 15783 -33628
rect 15656 -33708 15783 -33692
rect 15656 -33772 15703 -33708
rect 15767 -33772 15783 -33708
rect 15656 -33788 15783 -33772
rect 15656 -33852 15703 -33788
rect 15767 -33852 15783 -33788
rect 15656 -33868 15783 -33852
rect 15656 -33932 15703 -33868
rect 15767 -33932 15783 -33868
rect 15656 -33948 15783 -33932
rect 15656 -34012 15703 -33948
rect 15767 -34012 15783 -33948
rect 15656 -34028 15783 -34012
rect 15656 -34092 15703 -34028
rect 15767 -34092 15783 -34028
rect 15656 -34108 15783 -34092
rect 15656 -34172 15703 -34108
rect 15767 -34172 15783 -34108
rect 15656 -34188 15783 -34172
rect 15656 -34252 15703 -34188
rect 15767 -34252 15783 -34188
rect 15656 -34268 15783 -34252
rect 15656 -34332 15703 -34268
rect 15767 -34332 15783 -34268
rect 15656 -34348 15783 -34332
rect 15656 -34412 15703 -34348
rect 15767 -34412 15783 -34348
rect 15656 -34428 15783 -34412
rect 9337 -34508 9464 -34492
rect 9337 -34572 9384 -34508
rect 9448 -34572 9464 -34508
rect 9337 -34588 9464 -34572
rect 9337 -34712 9441 -34588
rect 9337 -34728 9464 -34712
rect 9337 -34792 9384 -34728
rect 9448 -34792 9464 -34728
rect 9337 -34808 9464 -34792
rect 3018 -34888 3145 -34872
rect 3018 -34952 3065 -34888
rect 3129 -34952 3145 -34888
rect 3018 -34968 3145 -34952
rect 3018 -35032 3065 -34968
rect 3129 -35032 3145 -34968
rect 3018 -35048 3145 -35032
rect 3018 -35112 3065 -35048
rect 3129 -35112 3145 -35048
rect 3018 -35128 3145 -35112
rect 3018 -35192 3065 -35128
rect 3129 -35192 3145 -35128
rect 3018 -35208 3145 -35192
rect 3018 -35272 3065 -35208
rect 3129 -35272 3145 -35208
rect 3018 -35288 3145 -35272
rect 3018 -35352 3065 -35288
rect 3129 -35352 3145 -35288
rect 3018 -35368 3145 -35352
rect 3018 -35432 3065 -35368
rect 3129 -35432 3145 -35368
rect 3018 -35448 3145 -35432
rect 3018 -35512 3065 -35448
rect 3129 -35512 3145 -35448
rect 3018 -35528 3145 -35512
rect 3018 -35592 3065 -35528
rect 3129 -35592 3145 -35528
rect 3018 -35608 3145 -35592
rect 3018 -35672 3065 -35608
rect 3129 -35672 3145 -35608
rect 3018 -35688 3145 -35672
rect 3018 -35752 3065 -35688
rect 3129 -35752 3145 -35688
rect 3018 -35768 3145 -35752
rect 3018 -35832 3065 -35768
rect 3129 -35832 3145 -35768
rect 3018 -35848 3145 -35832
rect 3018 -35912 3065 -35848
rect 3129 -35912 3145 -35848
rect 3018 -35928 3145 -35912
rect 3018 -35992 3065 -35928
rect 3129 -35992 3145 -35928
rect 3018 -36008 3145 -35992
rect 3018 -36072 3065 -36008
rect 3129 -36072 3145 -36008
rect 3018 -36088 3145 -36072
rect 3018 -36152 3065 -36088
rect 3129 -36152 3145 -36088
rect 3018 -36168 3145 -36152
rect 3018 -36232 3065 -36168
rect 3129 -36232 3145 -36168
rect 3018 -36248 3145 -36232
rect 3018 -36312 3065 -36248
rect 3129 -36312 3145 -36248
rect 3018 -36328 3145 -36312
rect 3018 -36392 3065 -36328
rect 3129 -36392 3145 -36328
rect 3018 -36408 3145 -36392
rect 3018 -36472 3065 -36408
rect 3129 -36472 3145 -36408
rect 3018 -36488 3145 -36472
rect 3018 -36552 3065 -36488
rect 3129 -36552 3145 -36488
rect 3018 -36568 3145 -36552
rect 3018 -36632 3065 -36568
rect 3129 -36632 3145 -36568
rect 3018 -36648 3145 -36632
rect 3018 -36712 3065 -36648
rect 3129 -36712 3145 -36648
rect 3018 -36728 3145 -36712
rect 3018 -36792 3065 -36728
rect 3129 -36792 3145 -36728
rect 3018 -36808 3145 -36792
rect 3018 -36872 3065 -36808
rect 3129 -36872 3145 -36808
rect 3018 -36888 3145 -36872
rect 3018 -36952 3065 -36888
rect 3129 -36952 3145 -36888
rect 3018 -36968 3145 -36952
rect 3018 -37032 3065 -36968
rect 3129 -37032 3145 -36968
rect 3018 -37048 3145 -37032
rect 3018 -37112 3065 -37048
rect 3129 -37112 3145 -37048
rect 3018 -37128 3145 -37112
rect 3018 -37192 3065 -37128
rect 3129 -37192 3145 -37128
rect 3018 -37208 3145 -37192
rect 3018 -37272 3065 -37208
rect 3129 -37272 3145 -37208
rect 3018 -37288 3145 -37272
rect 3018 -37352 3065 -37288
rect 3129 -37352 3145 -37288
rect 3018 -37368 3145 -37352
rect 3018 -37432 3065 -37368
rect 3129 -37432 3145 -37368
rect 3018 -37448 3145 -37432
rect 3018 -37512 3065 -37448
rect 3129 -37512 3145 -37448
rect 3018 -37528 3145 -37512
rect 3018 -37592 3065 -37528
rect 3129 -37592 3145 -37528
rect 3018 -37608 3145 -37592
rect 3018 -37672 3065 -37608
rect 3129 -37672 3145 -37608
rect 3018 -37688 3145 -37672
rect 3018 -37752 3065 -37688
rect 3129 -37752 3145 -37688
rect 3018 -37768 3145 -37752
rect 3018 -37832 3065 -37768
rect 3129 -37832 3145 -37768
rect 3018 -37848 3145 -37832
rect 3018 -37912 3065 -37848
rect 3129 -37912 3145 -37848
rect 3018 -37928 3145 -37912
rect 3018 -37992 3065 -37928
rect 3129 -37992 3145 -37928
rect 3018 -38008 3145 -37992
rect 3018 -38072 3065 -38008
rect 3129 -38072 3145 -38008
rect 3018 -38088 3145 -38072
rect 3018 -38152 3065 -38088
rect 3129 -38152 3145 -38088
rect 3018 -38168 3145 -38152
rect 3018 -38232 3065 -38168
rect 3129 -38232 3145 -38168
rect 3018 -38248 3145 -38232
rect 3018 -38312 3065 -38248
rect 3129 -38312 3145 -38248
rect 3018 -38328 3145 -38312
rect 3018 -38392 3065 -38328
rect 3129 -38392 3145 -38328
rect 3018 -38408 3145 -38392
rect 3018 -38472 3065 -38408
rect 3129 -38472 3145 -38408
rect 3018 -38488 3145 -38472
rect 3018 -38552 3065 -38488
rect 3129 -38552 3145 -38488
rect 3018 -38568 3145 -38552
rect 3018 -38632 3065 -38568
rect 3129 -38632 3145 -38568
rect 3018 -38648 3145 -38632
rect 3018 -38712 3065 -38648
rect 3129 -38712 3145 -38648
rect 3018 -38728 3145 -38712
rect 3018 -38792 3065 -38728
rect 3129 -38792 3145 -38728
rect 3018 -38808 3145 -38792
rect 3018 -38872 3065 -38808
rect 3129 -38872 3145 -38808
rect 3018 -38888 3145 -38872
rect 3018 -38952 3065 -38888
rect 3129 -38952 3145 -38888
rect 3018 -38968 3145 -38952
rect 3018 -39032 3065 -38968
rect 3129 -39032 3145 -38968
rect 3018 -39048 3145 -39032
rect 3018 -39112 3065 -39048
rect 3129 -39112 3145 -39048
rect 3018 -39128 3145 -39112
rect 3018 -39192 3065 -39128
rect 3129 -39192 3145 -39128
rect 3018 -39208 3145 -39192
rect 3018 -39272 3065 -39208
rect 3129 -39272 3145 -39208
rect 3018 -39288 3145 -39272
rect 3018 -39352 3065 -39288
rect 3129 -39352 3145 -39288
rect 3018 -39368 3145 -39352
rect 3018 -39432 3065 -39368
rect 3129 -39432 3145 -39368
rect 3018 -39448 3145 -39432
rect 3018 -39512 3065 -39448
rect 3129 -39512 3145 -39448
rect 3018 -39528 3145 -39512
rect 3018 -39592 3065 -39528
rect 3129 -39592 3145 -39528
rect 3018 -39608 3145 -39592
rect 3018 -39672 3065 -39608
rect 3129 -39672 3145 -39608
rect 3018 -39688 3145 -39672
rect 3018 -39752 3065 -39688
rect 3129 -39752 3145 -39688
rect 3018 -39768 3145 -39752
rect 3018 -39832 3065 -39768
rect 3129 -39832 3145 -39768
rect 3018 -39848 3145 -39832
rect 3018 -39912 3065 -39848
rect 3129 -39912 3145 -39848
rect 3018 -39928 3145 -39912
rect 3018 -39992 3065 -39928
rect 3129 -39992 3145 -39928
rect 3018 -40008 3145 -39992
rect 3018 -40072 3065 -40008
rect 3129 -40072 3145 -40008
rect 3018 -40088 3145 -40072
rect 3018 -40152 3065 -40088
rect 3129 -40152 3145 -40088
rect 3018 -40168 3145 -40152
rect 3018 -40232 3065 -40168
rect 3129 -40232 3145 -40168
rect 3018 -40248 3145 -40232
rect 3018 -40312 3065 -40248
rect 3129 -40312 3145 -40248
rect 3018 -40328 3145 -40312
rect 3018 -40392 3065 -40328
rect 3129 -40392 3145 -40328
rect 3018 -40408 3145 -40392
rect 3018 -40472 3065 -40408
rect 3129 -40472 3145 -40408
rect 3018 -40488 3145 -40472
rect 3018 -40552 3065 -40488
rect 3129 -40552 3145 -40488
rect 3018 -40568 3145 -40552
rect 3018 -40632 3065 -40568
rect 3129 -40632 3145 -40568
rect 3018 -40648 3145 -40632
rect 3018 -40712 3065 -40648
rect 3129 -40712 3145 -40648
rect 3018 -40728 3145 -40712
rect -3301 -40808 -3174 -40792
rect -3301 -40872 -3254 -40808
rect -3190 -40872 -3174 -40808
rect -3301 -40888 -3174 -40872
rect -3301 -41012 -3197 -40888
rect -3301 -41028 -3174 -41012
rect -3301 -41092 -3254 -41028
rect -3190 -41092 -3174 -41028
rect -3301 -41108 -3174 -41092
rect -9620 -41188 -9493 -41172
rect -9620 -41252 -9573 -41188
rect -9509 -41252 -9493 -41188
rect -9620 -41268 -9493 -41252
rect -9620 -41332 -9573 -41268
rect -9509 -41332 -9493 -41268
rect -9620 -41348 -9493 -41332
rect -9620 -41412 -9573 -41348
rect -9509 -41412 -9493 -41348
rect -9620 -41428 -9493 -41412
rect -9620 -41492 -9573 -41428
rect -9509 -41492 -9493 -41428
rect -9620 -41508 -9493 -41492
rect -9620 -41572 -9573 -41508
rect -9509 -41572 -9493 -41508
rect -9620 -41588 -9493 -41572
rect -9620 -41652 -9573 -41588
rect -9509 -41652 -9493 -41588
rect -9620 -41668 -9493 -41652
rect -9620 -41732 -9573 -41668
rect -9509 -41732 -9493 -41668
rect -9620 -41748 -9493 -41732
rect -9620 -41812 -9573 -41748
rect -9509 -41812 -9493 -41748
rect -9620 -41828 -9493 -41812
rect -9620 -41892 -9573 -41828
rect -9509 -41892 -9493 -41828
rect -9620 -41908 -9493 -41892
rect -9620 -41972 -9573 -41908
rect -9509 -41972 -9493 -41908
rect -9620 -41988 -9493 -41972
rect -9620 -42052 -9573 -41988
rect -9509 -42052 -9493 -41988
rect -9620 -42068 -9493 -42052
rect -9620 -42132 -9573 -42068
rect -9509 -42132 -9493 -42068
rect -9620 -42148 -9493 -42132
rect -9620 -42212 -9573 -42148
rect -9509 -42212 -9493 -42148
rect -9620 -42228 -9493 -42212
rect -9620 -42292 -9573 -42228
rect -9509 -42292 -9493 -42228
rect -9620 -42308 -9493 -42292
rect -9620 -42372 -9573 -42308
rect -9509 -42372 -9493 -42308
rect -9620 -42388 -9493 -42372
rect -9620 -42452 -9573 -42388
rect -9509 -42452 -9493 -42388
rect -9620 -42468 -9493 -42452
rect -9620 -42532 -9573 -42468
rect -9509 -42532 -9493 -42468
rect -9620 -42548 -9493 -42532
rect -9620 -42612 -9573 -42548
rect -9509 -42612 -9493 -42548
rect -9620 -42628 -9493 -42612
rect -9620 -42692 -9573 -42628
rect -9509 -42692 -9493 -42628
rect -9620 -42708 -9493 -42692
rect -9620 -42772 -9573 -42708
rect -9509 -42772 -9493 -42708
rect -9620 -42788 -9493 -42772
rect -9620 -42852 -9573 -42788
rect -9509 -42852 -9493 -42788
rect -9620 -42868 -9493 -42852
rect -9620 -42932 -9573 -42868
rect -9509 -42932 -9493 -42868
rect -9620 -42948 -9493 -42932
rect -9620 -43012 -9573 -42948
rect -9509 -43012 -9493 -42948
rect -9620 -43028 -9493 -43012
rect -9620 -43092 -9573 -43028
rect -9509 -43092 -9493 -43028
rect -9620 -43108 -9493 -43092
rect -9620 -43172 -9573 -43108
rect -9509 -43172 -9493 -43108
rect -9620 -43188 -9493 -43172
rect -9620 -43252 -9573 -43188
rect -9509 -43252 -9493 -43188
rect -9620 -43268 -9493 -43252
rect -9620 -43332 -9573 -43268
rect -9509 -43332 -9493 -43268
rect -9620 -43348 -9493 -43332
rect -9620 -43412 -9573 -43348
rect -9509 -43412 -9493 -43348
rect -9620 -43428 -9493 -43412
rect -9620 -43492 -9573 -43428
rect -9509 -43492 -9493 -43428
rect -9620 -43508 -9493 -43492
rect -9620 -43572 -9573 -43508
rect -9509 -43572 -9493 -43508
rect -9620 -43588 -9493 -43572
rect -9620 -43652 -9573 -43588
rect -9509 -43652 -9493 -43588
rect -9620 -43668 -9493 -43652
rect -9620 -43732 -9573 -43668
rect -9509 -43732 -9493 -43668
rect -9620 -43748 -9493 -43732
rect -9620 -43812 -9573 -43748
rect -9509 -43812 -9493 -43748
rect -9620 -43828 -9493 -43812
rect -9620 -43892 -9573 -43828
rect -9509 -43892 -9493 -43828
rect -9620 -43908 -9493 -43892
rect -9620 -43972 -9573 -43908
rect -9509 -43972 -9493 -43908
rect -9620 -43988 -9493 -43972
rect -9620 -44052 -9573 -43988
rect -9509 -44052 -9493 -43988
rect -9620 -44068 -9493 -44052
rect -9620 -44132 -9573 -44068
rect -9509 -44132 -9493 -44068
rect -9620 -44148 -9493 -44132
rect -9620 -44212 -9573 -44148
rect -9509 -44212 -9493 -44148
rect -9620 -44228 -9493 -44212
rect -9620 -44292 -9573 -44228
rect -9509 -44292 -9493 -44228
rect -9620 -44308 -9493 -44292
rect -9620 -44372 -9573 -44308
rect -9509 -44372 -9493 -44308
rect -9620 -44388 -9493 -44372
rect -9620 -44452 -9573 -44388
rect -9509 -44452 -9493 -44388
rect -9620 -44468 -9493 -44452
rect -9620 -44532 -9573 -44468
rect -9509 -44532 -9493 -44468
rect -9620 -44548 -9493 -44532
rect -9620 -44612 -9573 -44548
rect -9509 -44612 -9493 -44548
rect -9620 -44628 -9493 -44612
rect -9620 -44692 -9573 -44628
rect -9509 -44692 -9493 -44628
rect -9620 -44708 -9493 -44692
rect -9620 -44772 -9573 -44708
rect -9509 -44772 -9493 -44708
rect -9620 -44788 -9493 -44772
rect -9620 -44852 -9573 -44788
rect -9509 -44852 -9493 -44788
rect -9620 -44868 -9493 -44852
rect -9620 -44932 -9573 -44868
rect -9509 -44932 -9493 -44868
rect -9620 -44948 -9493 -44932
rect -9620 -45012 -9573 -44948
rect -9509 -45012 -9493 -44948
rect -9620 -45028 -9493 -45012
rect -9620 -45092 -9573 -45028
rect -9509 -45092 -9493 -45028
rect -9620 -45108 -9493 -45092
rect -9620 -45172 -9573 -45108
rect -9509 -45172 -9493 -45108
rect -9620 -45188 -9493 -45172
rect -9620 -45252 -9573 -45188
rect -9509 -45252 -9493 -45188
rect -9620 -45268 -9493 -45252
rect -9620 -45332 -9573 -45268
rect -9509 -45332 -9493 -45268
rect -9620 -45348 -9493 -45332
rect -9620 -45412 -9573 -45348
rect -9509 -45412 -9493 -45348
rect -9620 -45428 -9493 -45412
rect -9620 -45492 -9573 -45428
rect -9509 -45492 -9493 -45428
rect -9620 -45508 -9493 -45492
rect -9620 -45572 -9573 -45508
rect -9509 -45572 -9493 -45508
rect -9620 -45588 -9493 -45572
rect -9620 -45652 -9573 -45588
rect -9509 -45652 -9493 -45588
rect -9620 -45668 -9493 -45652
rect -9620 -45732 -9573 -45668
rect -9509 -45732 -9493 -45668
rect -9620 -45748 -9493 -45732
rect -9620 -45812 -9573 -45748
rect -9509 -45812 -9493 -45748
rect -9620 -45828 -9493 -45812
rect -9620 -45892 -9573 -45828
rect -9509 -45892 -9493 -45828
rect -9620 -45908 -9493 -45892
rect -9620 -45972 -9573 -45908
rect -9509 -45972 -9493 -45908
rect -9620 -45988 -9493 -45972
rect -9620 -46052 -9573 -45988
rect -9509 -46052 -9493 -45988
rect -9620 -46068 -9493 -46052
rect -9620 -46132 -9573 -46068
rect -9509 -46132 -9493 -46068
rect -9620 -46148 -9493 -46132
rect -9620 -46212 -9573 -46148
rect -9509 -46212 -9493 -46148
rect -9620 -46228 -9493 -46212
rect -9620 -46292 -9573 -46228
rect -9509 -46292 -9493 -46228
rect -9620 -46308 -9493 -46292
rect -9620 -46372 -9573 -46308
rect -9509 -46372 -9493 -46308
rect -9620 -46388 -9493 -46372
rect -9620 -46452 -9573 -46388
rect -9509 -46452 -9493 -46388
rect -9620 -46468 -9493 -46452
rect -9620 -46532 -9573 -46468
rect -9509 -46532 -9493 -46468
rect -9620 -46548 -9493 -46532
rect -9620 -46612 -9573 -46548
rect -9509 -46612 -9493 -46548
rect -9620 -46628 -9493 -46612
rect -9620 -46692 -9573 -46628
rect -9509 -46692 -9493 -46628
rect -9620 -46708 -9493 -46692
rect -9620 -46772 -9573 -46708
rect -9509 -46772 -9493 -46708
rect -9620 -46788 -9493 -46772
rect -9620 -46852 -9573 -46788
rect -9509 -46852 -9493 -46788
rect -9620 -46868 -9493 -46852
rect -9620 -46932 -9573 -46868
rect -9509 -46932 -9493 -46868
rect -9620 -46948 -9493 -46932
rect -9620 -47012 -9573 -46948
rect -9509 -47012 -9493 -46948
rect -9620 -47028 -9493 -47012
rect -15939 -47108 -15812 -47092
rect -15939 -47172 -15892 -47108
rect -15828 -47172 -15812 -47108
rect -15939 -47188 -15812 -47172
rect -15939 -47250 -15835 -47188
rect -12740 -47250 -12636 -47061
rect -9620 -47092 -9573 -47028
rect -9509 -47092 -9493 -47028
rect -9330 -41148 -3408 -41139
rect -9330 -47052 -9321 -41148
rect -3417 -47052 -3408 -41148
rect -9330 -47061 -3408 -47052
rect -3301 -41172 -3254 -41108
rect -3190 -41172 -3174 -41108
rect -102 -41139 2 -40761
rect 3018 -40792 3065 -40728
rect 3129 -40792 3145 -40728
rect 3308 -34848 9230 -34839
rect 3308 -40752 3317 -34848
rect 9221 -40752 9230 -34848
rect 3308 -40761 9230 -40752
rect 9337 -34872 9384 -34808
rect 9448 -34872 9464 -34808
rect 12536 -34839 12640 -34461
rect 15656 -34492 15703 -34428
rect 15767 -34492 15783 -34428
rect 15946 -28548 21868 -28539
rect 15946 -34452 15955 -28548
rect 21859 -34452 21868 -28548
rect 15946 -34461 21868 -34452
rect 21975 -28572 22022 -28508
rect 22086 -28572 22102 -28508
rect 25174 -28539 25278 -28161
rect 28294 -28192 28341 -28128
rect 28405 -28192 28421 -28128
rect 28584 -22248 34506 -22239
rect 28584 -28152 28593 -22248
rect 34497 -28152 34506 -22248
rect 28584 -28161 34506 -28152
rect 34613 -22272 34660 -22208
rect 34724 -22272 34740 -22208
rect 37812 -22239 37916 -21861
rect 40932 -21892 40979 -21828
rect 41043 -21892 41059 -21828
rect 41222 -15948 47144 -15939
rect 41222 -21852 41231 -15948
rect 47135 -21852 47144 -15948
rect 41222 -21861 47144 -21852
rect 47251 -15972 47298 -15908
rect 47362 -15972 47378 -15908
rect 47251 -15988 47378 -15972
rect 47251 -16052 47298 -15988
rect 47362 -16052 47378 -15988
rect 47251 -16068 47378 -16052
rect 47251 -16132 47298 -16068
rect 47362 -16132 47378 -16068
rect 47251 -16148 47378 -16132
rect 47251 -16212 47298 -16148
rect 47362 -16212 47378 -16148
rect 47251 -16228 47378 -16212
rect 47251 -16292 47298 -16228
rect 47362 -16292 47378 -16228
rect 47251 -16308 47378 -16292
rect 47251 -16372 47298 -16308
rect 47362 -16372 47378 -16308
rect 47251 -16388 47378 -16372
rect 47251 -16452 47298 -16388
rect 47362 -16452 47378 -16388
rect 47251 -16468 47378 -16452
rect 47251 -16532 47298 -16468
rect 47362 -16532 47378 -16468
rect 47251 -16548 47378 -16532
rect 47251 -16612 47298 -16548
rect 47362 -16612 47378 -16548
rect 47251 -16628 47378 -16612
rect 47251 -16692 47298 -16628
rect 47362 -16692 47378 -16628
rect 47251 -16708 47378 -16692
rect 47251 -16772 47298 -16708
rect 47362 -16772 47378 -16708
rect 47251 -16788 47378 -16772
rect 47251 -16852 47298 -16788
rect 47362 -16852 47378 -16788
rect 47251 -16868 47378 -16852
rect 47251 -16932 47298 -16868
rect 47362 -16932 47378 -16868
rect 47251 -16948 47378 -16932
rect 47251 -17012 47298 -16948
rect 47362 -17012 47378 -16948
rect 47251 -17028 47378 -17012
rect 47251 -17092 47298 -17028
rect 47362 -17092 47378 -17028
rect 47251 -17108 47378 -17092
rect 47251 -17172 47298 -17108
rect 47362 -17172 47378 -17108
rect 47251 -17188 47378 -17172
rect 47251 -17252 47298 -17188
rect 47362 -17252 47378 -17188
rect 47251 -17268 47378 -17252
rect 47251 -17332 47298 -17268
rect 47362 -17332 47378 -17268
rect 47251 -17348 47378 -17332
rect 47251 -17412 47298 -17348
rect 47362 -17412 47378 -17348
rect 47251 -17428 47378 -17412
rect 47251 -17492 47298 -17428
rect 47362 -17492 47378 -17428
rect 47251 -17508 47378 -17492
rect 47251 -17572 47298 -17508
rect 47362 -17572 47378 -17508
rect 47251 -17588 47378 -17572
rect 47251 -17652 47298 -17588
rect 47362 -17652 47378 -17588
rect 47251 -17668 47378 -17652
rect 47251 -17732 47298 -17668
rect 47362 -17732 47378 -17668
rect 47251 -17748 47378 -17732
rect 47251 -17812 47298 -17748
rect 47362 -17812 47378 -17748
rect 47251 -17828 47378 -17812
rect 47251 -17892 47298 -17828
rect 47362 -17892 47378 -17828
rect 47251 -17908 47378 -17892
rect 47251 -17972 47298 -17908
rect 47362 -17972 47378 -17908
rect 47251 -17988 47378 -17972
rect 47251 -18052 47298 -17988
rect 47362 -18052 47378 -17988
rect 47251 -18068 47378 -18052
rect 47251 -18132 47298 -18068
rect 47362 -18132 47378 -18068
rect 47251 -18148 47378 -18132
rect 47251 -18212 47298 -18148
rect 47362 -18212 47378 -18148
rect 47251 -18228 47378 -18212
rect 47251 -18292 47298 -18228
rect 47362 -18292 47378 -18228
rect 47251 -18308 47378 -18292
rect 47251 -18372 47298 -18308
rect 47362 -18372 47378 -18308
rect 47251 -18388 47378 -18372
rect 47251 -18452 47298 -18388
rect 47362 -18452 47378 -18388
rect 47251 -18468 47378 -18452
rect 47251 -18532 47298 -18468
rect 47362 -18532 47378 -18468
rect 47251 -18548 47378 -18532
rect 47251 -18612 47298 -18548
rect 47362 -18612 47378 -18548
rect 47251 -18628 47378 -18612
rect 47251 -18692 47298 -18628
rect 47362 -18692 47378 -18628
rect 47251 -18708 47378 -18692
rect 47251 -18772 47298 -18708
rect 47362 -18772 47378 -18708
rect 47251 -18788 47378 -18772
rect 47251 -18852 47298 -18788
rect 47362 -18852 47378 -18788
rect 47251 -18868 47378 -18852
rect 47251 -18932 47298 -18868
rect 47362 -18932 47378 -18868
rect 47251 -18948 47378 -18932
rect 47251 -19012 47298 -18948
rect 47362 -19012 47378 -18948
rect 47251 -19028 47378 -19012
rect 47251 -19092 47298 -19028
rect 47362 -19092 47378 -19028
rect 47251 -19108 47378 -19092
rect 47251 -19172 47298 -19108
rect 47362 -19172 47378 -19108
rect 47251 -19188 47378 -19172
rect 47251 -19252 47298 -19188
rect 47362 -19252 47378 -19188
rect 47251 -19268 47378 -19252
rect 47251 -19332 47298 -19268
rect 47362 -19332 47378 -19268
rect 47251 -19348 47378 -19332
rect 47251 -19412 47298 -19348
rect 47362 -19412 47378 -19348
rect 47251 -19428 47378 -19412
rect 47251 -19492 47298 -19428
rect 47362 -19492 47378 -19428
rect 47251 -19508 47378 -19492
rect 47251 -19572 47298 -19508
rect 47362 -19572 47378 -19508
rect 47251 -19588 47378 -19572
rect 47251 -19652 47298 -19588
rect 47362 -19652 47378 -19588
rect 47251 -19668 47378 -19652
rect 47251 -19732 47298 -19668
rect 47362 -19732 47378 -19668
rect 47251 -19748 47378 -19732
rect 47251 -19812 47298 -19748
rect 47362 -19812 47378 -19748
rect 47251 -19828 47378 -19812
rect 47251 -19892 47298 -19828
rect 47362 -19892 47378 -19828
rect 47251 -19908 47378 -19892
rect 47251 -19972 47298 -19908
rect 47362 -19972 47378 -19908
rect 47251 -19988 47378 -19972
rect 47251 -20052 47298 -19988
rect 47362 -20052 47378 -19988
rect 47251 -20068 47378 -20052
rect 47251 -20132 47298 -20068
rect 47362 -20132 47378 -20068
rect 47251 -20148 47378 -20132
rect 47251 -20212 47298 -20148
rect 47362 -20212 47378 -20148
rect 47251 -20228 47378 -20212
rect 47251 -20292 47298 -20228
rect 47362 -20292 47378 -20228
rect 47251 -20308 47378 -20292
rect 47251 -20372 47298 -20308
rect 47362 -20372 47378 -20308
rect 47251 -20388 47378 -20372
rect 47251 -20452 47298 -20388
rect 47362 -20452 47378 -20388
rect 47251 -20468 47378 -20452
rect 47251 -20532 47298 -20468
rect 47362 -20532 47378 -20468
rect 47251 -20548 47378 -20532
rect 47251 -20612 47298 -20548
rect 47362 -20612 47378 -20548
rect 47251 -20628 47378 -20612
rect 47251 -20692 47298 -20628
rect 47362 -20692 47378 -20628
rect 47251 -20708 47378 -20692
rect 47251 -20772 47298 -20708
rect 47362 -20772 47378 -20708
rect 47251 -20788 47378 -20772
rect 47251 -20852 47298 -20788
rect 47362 -20852 47378 -20788
rect 47251 -20868 47378 -20852
rect 47251 -20932 47298 -20868
rect 47362 -20932 47378 -20868
rect 47251 -20948 47378 -20932
rect 47251 -21012 47298 -20948
rect 47362 -21012 47378 -20948
rect 47251 -21028 47378 -21012
rect 47251 -21092 47298 -21028
rect 47362 -21092 47378 -21028
rect 47251 -21108 47378 -21092
rect 47251 -21172 47298 -21108
rect 47362 -21172 47378 -21108
rect 47251 -21188 47378 -21172
rect 47251 -21252 47298 -21188
rect 47362 -21252 47378 -21188
rect 47251 -21268 47378 -21252
rect 47251 -21332 47298 -21268
rect 47362 -21332 47378 -21268
rect 47251 -21348 47378 -21332
rect 47251 -21412 47298 -21348
rect 47362 -21412 47378 -21348
rect 47251 -21428 47378 -21412
rect 47251 -21492 47298 -21428
rect 47362 -21492 47378 -21428
rect 47251 -21508 47378 -21492
rect 47251 -21572 47298 -21508
rect 47362 -21572 47378 -21508
rect 47251 -21588 47378 -21572
rect 47251 -21652 47298 -21588
rect 47362 -21652 47378 -21588
rect 47251 -21668 47378 -21652
rect 47251 -21732 47298 -21668
rect 47362 -21732 47378 -21668
rect 47251 -21748 47378 -21732
rect 47251 -21812 47298 -21748
rect 47362 -21812 47378 -21748
rect 47251 -21828 47378 -21812
rect 40932 -21908 41059 -21892
rect 40932 -21972 40979 -21908
rect 41043 -21972 41059 -21908
rect 40932 -21988 41059 -21972
rect 40932 -22112 41036 -21988
rect 40932 -22128 41059 -22112
rect 40932 -22192 40979 -22128
rect 41043 -22192 41059 -22128
rect 40932 -22208 41059 -22192
rect 34613 -22288 34740 -22272
rect 34613 -22352 34660 -22288
rect 34724 -22352 34740 -22288
rect 34613 -22368 34740 -22352
rect 34613 -22432 34660 -22368
rect 34724 -22432 34740 -22368
rect 34613 -22448 34740 -22432
rect 34613 -22512 34660 -22448
rect 34724 -22512 34740 -22448
rect 34613 -22528 34740 -22512
rect 34613 -22592 34660 -22528
rect 34724 -22592 34740 -22528
rect 34613 -22608 34740 -22592
rect 34613 -22672 34660 -22608
rect 34724 -22672 34740 -22608
rect 34613 -22688 34740 -22672
rect 34613 -22752 34660 -22688
rect 34724 -22752 34740 -22688
rect 34613 -22768 34740 -22752
rect 34613 -22832 34660 -22768
rect 34724 -22832 34740 -22768
rect 34613 -22848 34740 -22832
rect 34613 -22912 34660 -22848
rect 34724 -22912 34740 -22848
rect 34613 -22928 34740 -22912
rect 34613 -22992 34660 -22928
rect 34724 -22992 34740 -22928
rect 34613 -23008 34740 -22992
rect 34613 -23072 34660 -23008
rect 34724 -23072 34740 -23008
rect 34613 -23088 34740 -23072
rect 34613 -23152 34660 -23088
rect 34724 -23152 34740 -23088
rect 34613 -23168 34740 -23152
rect 34613 -23232 34660 -23168
rect 34724 -23232 34740 -23168
rect 34613 -23248 34740 -23232
rect 34613 -23312 34660 -23248
rect 34724 -23312 34740 -23248
rect 34613 -23328 34740 -23312
rect 34613 -23392 34660 -23328
rect 34724 -23392 34740 -23328
rect 34613 -23408 34740 -23392
rect 34613 -23472 34660 -23408
rect 34724 -23472 34740 -23408
rect 34613 -23488 34740 -23472
rect 34613 -23552 34660 -23488
rect 34724 -23552 34740 -23488
rect 34613 -23568 34740 -23552
rect 34613 -23632 34660 -23568
rect 34724 -23632 34740 -23568
rect 34613 -23648 34740 -23632
rect 34613 -23712 34660 -23648
rect 34724 -23712 34740 -23648
rect 34613 -23728 34740 -23712
rect 34613 -23792 34660 -23728
rect 34724 -23792 34740 -23728
rect 34613 -23808 34740 -23792
rect 34613 -23872 34660 -23808
rect 34724 -23872 34740 -23808
rect 34613 -23888 34740 -23872
rect 34613 -23952 34660 -23888
rect 34724 -23952 34740 -23888
rect 34613 -23968 34740 -23952
rect 34613 -24032 34660 -23968
rect 34724 -24032 34740 -23968
rect 34613 -24048 34740 -24032
rect 34613 -24112 34660 -24048
rect 34724 -24112 34740 -24048
rect 34613 -24128 34740 -24112
rect 34613 -24192 34660 -24128
rect 34724 -24192 34740 -24128
rect 34613 -24208 34740 -24192
rect 34613 -24272 34660 -24208
rect 34724 -24272 34740 -24208
rect 34613 -24288 34740 -24272
rect 34613 -24352 34660 -24288
rect 34724 -24352 34740 -24288
rect 34613 -24368 34740 -24352
rect 34613 -24432 34660 -24368
rect 34724 -24432 34740 -24368
rect 34613 -24448 34740 -24432
rect 34613 -24512 34660 -24448
rect 34724 -24512 34740 -24448
rect 34613 -24528 34740 -24512
rect 34613 -24592 34660 -24528
rect 34724 -24592 34740 -24528
rect 34613 -24608 34740 -24592
rect 34613 -24672 34660 -24608
rect 34724 -24672 34740 -24608
rect 34613 -24688 34740 -24672
rect 34613 -24752 34660 -24688
rect 34724 -24752 34740 -24688
rect 34613 -24768 34740 -24752
rect 34613 -24832 34660 -24768
rect 34724 -24832 34740 -24768
rect 34613 -24848 34740 -24832
rect 34613 -24912 34660 -24848
rect 34724 -24912 34740 -24848
rect 34613 -24928 34740 -24912
rect 34613 -24992 34660 -24928
rect 34724 -24992 34740 -24928
rect 34613 -25008 34740 -24992
rect 34613 -25072 34660 -25008
rect 34724 -25072 34740 -25008
rect 34613 -25088 34740 -25072
rect 34613 -25152 34660 -25088
rect 34724 -25152 34740 -25088
rect 34613 -25168 34740 -25152
rect 34613 -25232 34660 -25168
rect 34724 -25232 34740 -25168
rect 34613 -25248 34740 -25232
rect 34613 -25312 34660 -25248
rect 34724 -25312 34740 -25248
rect 34613 -25328 34740 -25312
rect 34613 -25392 34660 -25328
rect 34724 -25392 34740 -25328
rect 34613 -25408 34740 -25392
rect 34613 -25472 34660 -25408
rect 34724 -25472 34740 -25408
rect 34613 -25488 34740 -25472
rect 34613 -25552 34660 -25488
rect 34724 -25552 34740 -25488
rect 34613 -25568 34740 -25552
rect 34613 -25632 34660 -25568
rect 34724 -25632 34740 -25568
rect 34613 -25648 34740 -25632
rect 34613 -25712 34660 -25648
rect 34724 -25712 34740 -25648
rect 34613 -25728 34740 -25712
rect 34613 -25792 34660 -25728
rect 34724 -25792 34740 -25728
rect 34613 -25808 34740 -25792
rect 34613 -25872 34660 -25808
rect 34724 -25872 34740 -25808
rect 34613 -25888 34740 -25872
rect 34613 -25952 34660 -25888
rect 34724 -25952 34740 -25888
rect 34613 -25968 34740 -25952
rect 34613 -26032 34660 -25968
rect 34724 -26032 34740 -25968
rect 34613 -26048 34740 -26032
rect 34613 -26112 34660 -26048
rect 34724 -26112 34740 -26048
rect 34613 -26128 34740 -26112
rect 34613 -26192 34660 -26128
rect 34724 -26192 34740 -26128
rect 34613 -26208 34740 -26192
rect 34613 -26272 34660 -26208
rect 34724 -26272 34740 -26208
rect 34613 -26288 34740 -26272
rect 34613 -26352 34660 -26288
rect 34724 -26352 34740 -26288
rect 34613 -26368 34740 -26352
rect 34613 -26432 34660 -26368
rect 34724 -26432 34740 -26368
rect 34613 -26448 34740 -26432
rect 34613 -26512 34660 -26448
rect 34724 -26512 34740 -26448
rect 34613 -26528 34740 -26512
rect 34613 -26592 34660 -26528
rect 34724 -26592 34740 -26528
rect 34613 -26608 34740 -26592
rect 34613 -26672 34660 -26608
rect 34724 -26672 34740 -26608
rect 34613 -26688 34740 -26672
rect 34613 -26752 34660 -26688
rect 34724 -26752 34740 -26688
rect 34613 -26768 34740 -26752
rect 34613 -26832 34660 -26768
rect 34724 -26832 34740 -26768
rect 34613 -26848 34740 -26832
rect 34613 -26912 34660 -26848
rect 34724 -26912 34740 -26848
rect 34613 -26928 34740 -26912
rect 34613 -26992 34660 -26928
rect 34724 -26992 34740 -26928
rect 34613 -27008 34740 -26992
rect 34613 -27072 34660 -27008
rect 34724 -27072 34740 -27008
rect 34613 -27088 34740 -27072
rect 34613 -27152 34660 -27088
rect 34724 -27152 34740 -27088
rect 34613 -27168 34740 -27152
rect 34613 -27232 34660 -27168
rect 34724 -27232 34740 -27168
rect 34613 -27248 34740 -27232
rect 34613 -27312 34660 -27248
rect 34724 -27312 34740 -27248
rect 34613 -27328 34740 -27312
rect 34613 -27392 34660 -27328
rect 34724 -27392 34740 -27328
rect 34613 -27408 34740 -27392
rect 34613 -27472 34660 -27408
rect 34724 -27472 34740 -27408
rect 34613 -27488 34740 -27472
rect 34613 -27552 34660 -27488
rect 34724 -27552 34740 -27488
rect 34613 -27568 34740 -27552
rect 34613 -27632 34660 -27568
rect 34724 -27632 34740 -27568
rect 34613 -27648 34740 -27632
rect 34613 -27712 34660 -27648
rect 34724 -27712 34740 -27648
rect 34613 -27728 34740 -27712
rect 34613 -27792 34660 -27728
rect 34724 -27792 34740 -27728
rect 34613 -27808 34740 -27792
rect 34613 -27872 34660 -27808
rect 34724 -27872 34740 -27808
rect 34613 -27888 34740 -27872
rect 34613 -27952 34660 -27888
rect 34724 -27952 34740 -27888
rect 34613 -27968 34740 -27952
rect 34613 -28032 34660 -27968
rect 34724 -28032 34740 -27968
rect 34613 -28048 34740 -28032
rect 34613 -28112 34660 -28048
rect 34724 -28112 34740 -28048
rect 34613 -28128 34740 -28112
rect 28294 -28208 28421 -28192
rect 28294 -28272 28341 -28208
rect 28405 -28272 28421 -28208
rect 28294 -28288 28421 -28272
rect 28294 -28412 28398 -28288
rect 28294 -28428 28421 -28412
rect 28294 -28492 28341 -28428
rect 28405 -28492 28421 -28428
rect 28294 -28508 28421 -28492
rect 21975 -28588 22102 -28572
rect 21975 -28652 22022 -28588
rect 22086 -28652 22102 -28588
rect 21975 -28668 22102 -28652
rect 21975 -28732 22022 -28668
rect 22086 -28732 22102 -28668
rect 21975 -28748 22102 -28732
rect 21975 -28812 22022 -28748
rect 22086 -28812 22102 -28748
rect 21975 -28828 22102 -28812
rect 21975 -28892 22022 -28828
rect 22086 -28892 22102 -28828
rect 21975 -28908 22102 -28892
rect 21975 -28972 22022 -28908
rect 22086 -28972 22102 -28908
rect 21975 -28988 22102 -28972
rect 21975 -29052 22022 -28988
rect 22086 -29052 22102 -28988
rect 21975 -29068 22102 -29052
rect 21975 -29132 22022 -29068
rect 22086 -29132 22102 -29068
rect 21975 -29148 22102 -29132
rect 21975 -29212 22022 -29148
rect 22086 -29212 22102 -29148
rect 21975 -29228 22102 -29212
rect 21975 -29292 22022 -29228
rect 22086 -29292 22102 -29228
rect 21975 -29308 22102 -29292
rect 21975 -29372 22022 -29308
rect 22086 -29372 22102 -29308
rect 21975 -29388 22102 -29372
rect 21975 -29452 22022 -29388
rect 22086 -29452 22102 -29388
rect 21975 -29468 22102 -29452
rect 21975 -29532 22022 -29468
rect 22086 -29532 22102 -29468
rect 21975 -29548 22102 -29532
rect 21975 -29612 22022 -29548
rect 22086 -29612 22102 -29548
rect 21975 -29628 22102 -29612
rect 21975 -29692 22022 -29628
rect 22086 -29692 22102 -29628
rect 21975 -29708 22102 -29692
rect 21975 -29772 22022 -29708
rect 22086 -29772 22102 -29708
rect 21975 -29788 22102 -29772
rect 21975 -29852 22022 -29788
rect 22086 -29852 22102 -29788
rect 21975 -29868 22102 -29852
rect 21975 -29932 22022 -29868
rect 22086 -29932 22102 -29868
rect 21975 -29948 22102 -29932
rect 21975 -30012 22022 -29948
rect 22086 -30012 22102 -29948
rect 21975 -30028 22102 -30012
rect 21975 -30092 22022 -30028
rect 22086 -30092 22102 -30028
rect 21975 -30108 22102 -30092
rect 21975 -30172 22022 -30108
rect 22086 -30172 22102 -30108
rect 21975 -30188 22102 -30172
rect 21975 -30252 22022 -30188
rect 22086 -30252 22102 -30188
rect 21975 -30268 22102 -30252
rect 21975 -30332 22022 -30268
rect 22086 -30332 22102 -30268
rect 21975 -30348 22102 -30332
rect 21975 -30412 22022 -30348
rect 22086 -30412 22102 -30348
rect 21975 -30428 22102 -30412
rect 21975 -30492 22022 -30428
rect 22086 -30492 22102 -30428
rect 21975 -30508 22102 -30492
rect 21975 -30572 22022 -30508
rect 22086 -30572 22102 -30508
rect 21975 -30588 22102 -30572
rect 21975 -30652 22022 -30588
rect 22086 -30652 22102 -30588
rect 21975 -30668 22102 -30652
rect 21975 -30732 22022 -30668
rect 22086 -30732 22102 -30668
rect 21975 -30748 22102 -30732
rect 21975 -30812 22022 -30748
rect 22086 -30812 22102 -30748
rect 21975 -30828 22102 -30812
rect 21975 -30892 22022 -30828
rect 22086 -30892 22102 -30828
rect 21975 -30908 22102 -30892
rect 21975 -30972 22022 -30908
rect 22086 -30972 22102 -30908
rect 21975 -30988 22102 -30972
rect 21975 -31052 22022 -30988
rect 22086 -31052 22102 -30988
rect 21975 -31068 22102 -31052
rect 21975 -31132 22022 -31068
rect 22086 -31132 22102 -31068
rect 21975 -31148 22102 -31132
rect 21975 -31212 22022 -31148
rect 22086 -31212 22102 -31148
rect 21975 -31228 22102 -31212
rect 21975 -31292 22022 -31228
rect 22086 -31292 22102 -31228
rect 21975 -31308 22102 -31292
rect 21975 -31372 22022 -31308
rect 22086 -31372 22102 -31308
rect 21975 -31388 22102 -31372
rect 21975 -31452 22022 -31388
rect 22086 -31452 22102 -31388
rect 21975 -31468 22102 -31452
rect 21975 -31532 22022 -31468
rect 22086 -31532 22102 -31468
rect 21975 -31548 22102 -31532
rect 21975 -31612 22022 -31548
rect 22086 -31612 22102 -31548
rect 21975 -31628 22102 -31612
rect 21975 -31692 22022 -31628
rect 22086 -31692 22102 -31628
rect 21975 -31708 22102 -31692
rect 21975 -31772 22022 -31708
rect 22086 -31772 22102 -31708
rect 21975 -31788 22102 -31772
rect 21975 -31852 22022 -31788
rect 22086 -31852 22102 -31788
rect 21975 -31868 22102 -31852
rect 21975 -31932 22022 -31868
rect 22086 -31932 22102 -31868
rect 21975 -31948 22102 -31932
rect 21975 -32012 22022 -31948
rect 22086 -32012 22102 -31948
rect 21975 -32028 22102 -32012
rect 21975 -32092 22022 -32028
rect 22086 -32092 22102 -32028
rect 21975 -32108 22102 -32092
rect 21975 -32172 22022 -32108
rect 22086 -32172 22102 -32108
rect 21975 -32188 22102 -32172
rect 21975 -32252 22022 -32188
rect 22086 -32252 22102 -32188
rect 21975 -32268 22102 -32252
rect 21975 -32332 22022 -32268
rect 22086 -32332 22102 -32268
rect 21975 -32348 22102 -32332
rect 21975 -32412 22022 -32348
rect 22086 -32412 22102 -32348
rect 21975 -32428 22102 -32412
rect 21975 -32492 22022 -32428
rect 22086 -32492 22102 -32428
rect 21975 -32508 22102 -32492
rect 21975 -32572 22022 -32508
rect 22086 -32572 22102 -32508
rect 21975 -32588 22102 -32572
rect 21975 -32652 22022 -32588
rect 22086 -32652 22102 -32588
rect 21975 -32668 22102 -32652
rect 21975 -32732 22022 -32668
rect 22086 -32732 22102 -32668
rect 21975 -32748 22102 -32732
rect 21975 -32812 22022 -32748
rect 22086 -32812 22102 -32748
rect 21975 -32828 22102 -32812
rect 21975 -32892 22022 -32828
rect 22086 -32892 22102 -32828
rect 21975 -32908 22102 -32892
rect 21975 -32972 22022 -32908
rect 22086 -32972 22102 -32908
rect 21975 -32988 22102 -32972
rect 21975 -33052 22022 -32988
rect 22086 -33052 22102 -32988
rect 21975 -33068 22102 -33052
rect 21975 -33132 22022 -33068
rect 22086 -33132 22102 -33068
rect 21975 -33148 22102 -33132
rect 21975 -33212 22022 -33148
rect 22086 -33212 22102 -33148
rect 21975 -33228 22102 -33212
rect 21975 -33292 22022 -33228
rect 22086 -33292 22102 -33228
rect 21975 -33308 22102 -33292
rect 21975 -33372 22022 -33308
rect 22086 -33372 22102 -33308
rect 21975 -33388 22102 -33372
rect 21975 -33452 22022 -33388
rect 22086 -33452 22102 -33388
rect 21975 -33468 22102 -33452
rect 21975 -33532 22022 -33468
rect 22086 -33532 22102 -33468
rect 21975 -33548 22102 -33532
rect 21975 -33612 22022 -33548
rect 22086 -33612 22102 -33548
rect 21975 -33628 22102 -33612
rect 21975 -33692 22022 -33628
rect 22086 -33692 22102 -33628
rect 21975 -33708 22102 -33692
rect 21975 -33772 22022 -33708
rect 22086 -33772 22102 -33708
rect 21975 -33788 22102 -33772
rect 21975 -33852 22022 -33788
rect 22086 -33852 22102 -33788
rect 21975 -33868 22102 -33852
rect 21975 -33932 22022 -33868
rect 22086 -33932 22102 -33868
rect 21975 -33948 22102 -33932
rect 21975 -34012 22022 -33948
rect 22086 -34012 22102 -33948
rect 21975 -34028 22102 -34012
rect 21975 -34092 22022 -34028
rect 22086 -34092 22102 -34028
rect 21975 -34108 22102 -34092
rect 21975 -34172 22022 -34108
rect 22086 -34172 22102 -34108
rect 21975 -34188 22102 -34172
rect 21975 -34252 22022 -34188
rect 22086 -34252 22102 -34188
rect 21975 -34268 22102 -34252
rect 21975 -34332 22022 -34268
rect 22086 -34332 22102 -34268
rect 21975 -34348 22102 -34332
rect 21975 -34412 22022 -34348
rect 22086 -34412 22102 -34348
rect 21975 -34428 22102 -34412
rect 15656 -34508 15783 -34492
rect 15656 -34572 15703 -34508
rect 15767 -34572 15783 -34508
rect 15656 -34588 15783 -34572
rect 15656 -34712 15760 -34588
rect 15656 -34728 15783 -34712
rect 15656 -34792 15703 -34728
rect 15767 -34792 15783 -34728
rect 15656 -34808 15783 -34792
rect 9337 -34888 9464 -34872
rect 9337 -34952 9384 -34888
rect 9448 -34952 9464 -34888
rect 9337 -34968 9464 -34952
rect 9337 -35032 9384 -34968
rect 9448 -35032 9464 -34968
rect 9337 -35048 9464 -35032
rect 9337 -35112 9384 -35048
rect 9448 -35112 9464 -35048
rect 9337 -35128 9464 -35112
rect 9337 -35192 9384 -35128
rect 9448 -35192 9464 -35128
rect 9337 -35208 9464 -35192
rect 9337 -35272 9384 -35208
rect 9448 -35272 9464 -35208
rect 9337 -35288 9464 -35272
rect 9337 -35352 9384 -35288
rect 9448 -35352 9464 -35288
rect 9337 -35368 9464 -35352
rect 9337 -35432 9384 -35368
rect 9448 -35432 9464 -35368
rect 9337 -35448 9464 -35432
rect 9337 -35512 9384 -35448
rect 9448 -35512 9464 -35448
rect 9337 -35528 9464 -35512
rect 9337 -35592 9384 -35528
rect 9448 -35592 9464 -35528
rect 9337 -35608 9464 -35592
rect 9337 -35672 9384 -35608
rect 9448 -35672 9464 -35608
rect 9337 -35688 9464 -35672
rect 9337 -35752 9384 -35688
rect 9448 -35752 9464 -35688
rect 9337 -35768 9464 -35752
rect 9337 -35832 9384 -35768
rect 9448 -35832 9464 -35768
rect 9337 -35848 9464 -35832
rect 9337 -35912 9384 -35848
rect 9448 -35912 9464 -35848
rect 9337 -35928 9464 -35912
rect 9337 -35992 9384 -35928
rect 9448 -35992 9464 -35928
rect 9337 -36008 9464 -35992
rect 9337 -36072 9384 -36008
rect 9448 -36072 9464 -36008
rect 9337 -36088 9464 -36072
rect 9337 -36152 9384 -36088
rect 9448 -36152 9464 -36088
rect 9337 -36168 9464 -36152
rect 9337 -36232 9384 -36168
rect 9448 -36232 9464 -36168
rect 9337 -36248 9464 -36232
rect 9337 -36312 9384 -36248
rect 9448 -36312 9464 -36248
rect 9337 -36328 9464 -36312
rect 9337 -36392 9384 -36328
rect 9448 -36392 9464 -36328
rect 9337 -36408 9464 -36392
rect 9337 -36472 9384 -36408
rect 9448 -36472 9464 -36408
rect 9337 -36488 9464 -36472
rect 9337 -36552 9384 -36488
rect 9448 -36552 9464 -36488
rect 9337 -36568 9464 -36552
rect 9337 -36632 9384 -36568
rect 9448 -36632 9464 -36568
rect 9337 -36648 9464 -36632
rect 9337 -36712 9384 -36648
rect 9448 -36712 9464 -36648
rect 9337 -36728 9464 -36712
rect 9337 -36792 9384 -36728
rect 9448 -36792 9464 -36728
rect 9337 -36808 9464 -36792
rect 9337 -36872 9384 -36808
rect 9448 -36872 9464 -36808
rect 9337 -36888 9464 -36872
rect 9337 -36952 9384 -36888
rect 9448 -36952 9464 -36888
rect 9337 -36968 9464 -36952
rect 9337 -37032 9384 -36968
rect 9448 -37032 9464 -36968
rect 9337 -37048 9464 -37032
rect 9337 -37112 9384 -37048
rect 9448 -37112 9464 -37048
rect 9337 -37128 9464 -37112
rect 9337 -37192 9384 -37128
rect 9448 -37192 9464 -37128
rect 9337 -37208 9464 -37192
rect 9337 -37272 9384 -37208
rect 9448 -37272 9464 -37208
rect 9337 -37288 9464 -37272
rect 9337 -37352 9384 -37288
rect 9448 -37352 9464 -37288
rect 9337 -37368 9464 -37352
rect 9337 -37432 9384 -37368
rect 9448 -37432 9464 -37368
rect 9337 -37448 9464 -37432
rect 9337 -37512 9384 -37448
rect 9448 -37512 9464 -37448
rect 9337 -37528 9464 -37512
rect 9337 -37592 9384 -37528
rect 9448 -37592 9464 -37528
rect 9337 -37608 9464 -37592
rect 9337 -37672 9384 -37608
rect 9448 -37672 9464 -37608
rect 9337 -37688 9464 -37672
rect 9337 -37752 9384 -37688
rect 9448 -37752 9464 -37688
rect 9337 -37768 9464 -37752
rect 9337 -37832 9384 -37768
rect 9448 -37832 9464 -37768
rect 9337 -37848 9464 -37832
rect 9337 -37912 9384 -37848
rect 9448 -37912 9464 -37848
rect 9337 -37928 9464 -37912
rect 9337 -37992 9384 -37928
rect 9448 -37992 9464 -37928
rect 9337 -38008 9464 -37992
rect 9337 -38072 9384 -38008
rect 9448 -38072 9464 -38008
rect 9337 -38088 9464 -38072
rect 9337 -38152 9384 -38088
rect 9448 -38152 9464 -38088
rect 9337 -38168 9464 -38152
rect 9337 -38232 9384 -38168
rect 9448 -38232 9464 -38168
rect 9337 -38248 9464 -38232
rect 9337 -38312 9384 -38248
rect 9448 -38312 9464 -38248
rect 9337 -38328 9464 -38312
rect 9337 -38392 9384 -38328
rect 9448 -38392 9464 -38328
rect 9337 -38408 9464 -38392
rect 9337 -38472 9384 -38408
rect 9448 -38472 9464 -38408
rect 9337 -38488 9464 -38472
rect 9337 -38552 9384 -38488
rect 9448 -38552 9464 -38488
rect 9337 -38568 9464 -38552
rect 9337 -38632 9384 -38568
rect 9448 -38632 9464 -38568
rect 9337 -38648 9464 -38632
rect 9337 -38712 9384 -38648
rect 9448 -38712 9464 -38648
rect 9337 -38728 9464 -38712
rect 9337 -38792 9384 -38728
rect 9448 -38792 9464 -38728
rect 9337 -38808 9464 -38792
rect 9337 -38872 9384 -38808
rect 9448 -38872 9464 -38808
rect 9337 -38888 9464 -38872
rect 9337 -38952 9384 -38888
rect 9448 -38952 9464 -38888
rect 9337 -38968 9464 -38952
rect 9337 -39032 9384 -38968
rect 9448 -39032 9464 -38968
rect 9337 -39048 9464 -39032
rect 9337 -39112 9384 -39048
rect 9448 -39112 9464 -39048
rect 9337 -39128 9464 -39112
rect 9337 -39192 9384 -39128
rect 9448 -39192 9464 -39128
rect 9337 -39208 9464 -39192
rect 9337 -39272 9384 -39208
rect 9448 -39272 9464 -39208
rect 9337 -39288 9464 -39272
rect 9337 -39352 9384 -39288
rect 9448 -39352 9464 -39288
rect 9337 -39368 9464 -39352
rect 9337 -39432 9384 -39368
rect 9448 -39432 9464 -39368
rect 9337 -39448 9464 -39432
rect 9337 -39512 9384 -39448
rect 9448 -39512 9464 -39448
rect 9337 -39528 9464 -39512
rect 9337 -39592 9384 -39528
rect 9448 -39592 9464 -39528
rect 9337 -39608 9464 -39592
rect 9337 -39672 9384 -39608
rect 9448 -39672 9464 -39608
rect 9337 -39688 9464 -39672
rect 9337 -39752 9384 -39688
rect 9448 -39752 9464 -39688
rect 9337 -39768 9464 -39752
rect 9337 -39832 9384 -39768
rect 9448 -39832 9464 -39768
rect 9337 -39848 9464 -39832
rect 9337 -39912 9384 -39848
rect 9448 -39912 9464 -39848
rect 9337 -39928 9464 -39912
rect 9337 -39992 9384 -39928
rect 9448 -39992 9464 -39928
rect 9337 -40008 9464 -39992
rect 9337 -40072 9384 -40008
rect 9448 -40072 9464 -40008
rect 9337 -40088 9464 -40072
rect 9337 -40152 9384 -40088
rect 9448 -40152 9464 -40088
rect 9337 -40168 9464 -40152
rect 9337 -40232 9384 -40168
rect 9448 -40232 9464 -40168
rect 9337 -40248 9464 -40232
rect 9337 -40312 9384 -40248
rect 9448 -40312 9464 -40248
rect 9337 -40328 9464 -40312
rect 9337 -40392 9384 -40328
rect 9448 -40392 9464 -40328
rect 9337 -40408 9464 -40392
rect 9337 -40472 9384 -40408
rect 9448 -40472 9464 -40408
rect 9337 -40488 9464 -40472
rect 9337 -40552 9384 -40488
rect 9448 -40552 9464 -40488
rect 9337 -40568 9464 -40552
rect 9337 -40632 9384 -40568
rect 9448 -40632 9464 -40568
rect 9337 -40648 9464 -40632
rect 9337 -40712 9384 -40648
rect 9448 -40712 9464 -40648
rect 9337 -40728 9464 -40712
rect 3018 -40808 3145 -40792
rect 3018 -40872 3065 -40808
rect 3129 -40872 3145 -40808
rect 3018 -40888 3145 -40872
rect 3018 -41012 3122 -40888
rect 3018 -41028 3145 -41012
rect 3018 -41092 3065 -41028
rect 3129 -41092 3145 -41028
rect 3018 -41108 3145 -41092
rect -3301 -41188 -3174 -41172
rect -3301 -41252 -3254 -41188
rect -3190 -41252 -3174 -41188
rect -3301 -41268 -3174 -41252
rect -3301 -41332 -3254 -41268
rect -3190 -41332 -3174 -41268
rect -3301 -41348 -3174 -41332
rect -3301 -41412 -3254 -41348
rect -3190 -41412 -3174 -41348
rect -3301 -41428 -3174 -41412
rect -3301 -41492 -3254 -41428
rect -3190 -41492 -3174 -41428
rect -3301 -41508 -3174 -41492
rect -3301 -41572 -3254 -41508
rect -3190 -41572 -3174 -41508
rect -3301 -41588 -3174 -41572
rect -3301 -41652 -3254 -41588
rect -3190 -41652 -3174 -41588
rect -3301 -41668 -3174 -41652
rect -3301 -41732 -3254 -41668
rect -3190 -41732 -3174 -41668
rect -3301 -41748 -3174 -41732
rect -3301 -41812 -3254 -41748
rect -3190 -41812 -3174 -41748
rect -3301 -41828 -3174 -41812
rect -3301 -41892 -3254 -41828
rect -3190 -41892 -3174 -41828
rect -3301 -41908 -3174 -41892
rect -3301 -41972 -3254 -41908
rect -3190 -41972 -3174 -41908
rect -3301 -41988 -3174 -41972
rect -3301 -42052 -3254 -41988
rect -3190 -42052 -3174 -41988
rect -3301 -42068 -3174 -42052
rect -3301 -42132 -3254 -42068
rect -3190 -42132 -3174 -42068
rect -3301 -42148 -3174 -42132
rect -3301 -42212 -3254 -42148
rect -3190 -42212 -3174 -42148
rect -3301 -42228 -3174 -42212
rect -3301 -42292 -3254 -42228
rect -3190 -42292 -3174 -42228
rect -3301 -42308 -3174 -42292
rect -3301 -42372 -3254 -42308
rect -3190 -42372 -3174 -42308
rect -3301 -42388 -3174 -42372
rect -3301 -42452 -3254 -42388
rect -3190 -42452 -3174 -42388
rect -3301 -42468 -3174 -42452
rect -3301 -42532 -3254 -42468
rect -3190 -42532 -3174 -42468
rect -3301 -42548 -3174 -42532
rect -3301 -42612 -3254 -42548
rect -3190 -42612 -3174 -42548
rect -3301 -42628 -3174 -42612
rect -3301 -42692 -3254 -42628
rect -3190 -42692 -3174 -42628
rect -3301 -42708 -3174 -42692
rect -3301 -42772 -3254 -42708
rect -3190 -42772 -3174 -42708
rect -3301 -42788 -3174 -42772
rect -3301 -42852 -3254 -42788
rect -3190 -42852 -3174 -42788
rect -3301 -42868 -3174 -42852
rect -3301 -42932 -3254 -42868
rect -3190 -42932 -3174 -42868
rect -3301 -42948 -3174 -42932
rect -3301 -43012 -3254 -42948
rect -3190 -43012 -3174 -42948
rect -3301 -43028 -3174 -43012
rect -3301 -43092 -3254 -43028
rect -3190 -43092 -3174 -43028
rect -3301 -43108 -3174 -43092
rect -3301 -43172 -3254 -43108
rect -3190 -43172 -3174 -43108
rect -3301 -43188 -3174 -43172
rect -3301 -43252 -3254 -43188
rect -3190 -43252 -3174 -43188
rect -3301 -43268 -3174 -43252
rect -3301 -43332 -3254 -43268
rect -3190 -43332 -3174 -43268
rect -3301 -43348 -3174 -43332
rect -3301 -43412 -3254 -43348
rect -3190 -43412 -3174 -43348
rect -3301 -43428 -3174 -43412
rect -3301 -43492 -3254 -43428
rect -3190 -43492 -3174 -43428
rect -3301 -43508 -3174 -43492
rect -3301 -43572 -3254 -43508
rect -3190 -43572 -3174 -43508
rect -3301 -43588 -3174 -43572
rect -3301 -43652 -3254 -43588
rect -3190 -43652 -3174 -43588
rect -3301 -43668 -3174 -43652
rect -3301 -43732 -3254 -43668
rect -3190 -43732 -3174 -43668
rect -3301 -43748 -3174 -43732
rect -3301 -43812 -3254 -43748
rect -3190 -43812 -3174 -43748
rect -3301 -43828 -3174 -43812
rect -3301 -43892 -3254 -43828
rect -3190 -43892 -3174 -43828
rect -3301 -43908 -3174 -43892
rect -3301 -43972 -3254 -43908
rect -3190 -43972 -3174 -43908
rect -3301 -43988 -3174 -43972
rect -3301 -44052 -3254 -43988
rect -3190 -44052 -3174 -43988
rect -3301 -44068 -3174 -44052
rect -3301 -44132 -3254 -44068
rect -3190 -44132 -3174 -44068
rect -3301 -44148 -3174 -44132
rect -3301 -44212 -3254 -44148
rect -3190 -44212 -3174 -44148
rect -3301 -44228 -3174 -44212
rect -3301 -44292 -3254 -44228
rect -3190 -44292 -3174 -44228
rect -3301 -44308 -3174 -44292
rect -3301 -44372 -3254 -44308
rect -3190 -44372 -3174 -44308
rect -3301 -44388 -3174 -44372
rect -3301 -44452 -3254 -44388
rect -3190 -44452 -3174 -44388
rect -3301 -44468 -3174 -44452
rect -3301 -44532 -3254 -44468
rect -3190 -44532 -3174 -44468
rect -3301 -44548 -3174 -44532
rect -3301 -44612 -3254 -44548
rect -3190 -44612 -3174 -44548
rect -3301 -44628 -3174 -44612
rect -3301 -44692 -3254 -44628
rect -3190 -44692 -3174 -44628
rect -3301 -44708 -3174 -44692
rect -3301 -44772 -3254 -44708
rect -3190 -44772 -3174 -44708
rect -3301 -44788 -3174 -44772
rect -3301 -44852 -3254 -44788
rect -3190 -44852 -3174 -44788
rect -3301 -44868 -3174 -44852
rect -3301 -44932 -3254 -44868
rect -3190 -44932 -3174 -44868
rect -3301 -44948 -3174 -44932
rect -3301 -45012 -3254 -44948
rect -3190 -45012 -3174 -44948
rect -3301 -45028 -3174 -45012
rect -3301 -45092 -3254 -45028
rect -3190 -45092 -3174 -45028
rect -3301 -45108 -3174 -45092
rect -3301 -45172 -3254 -45108
rect -3190 -45172 -3174 -45108
rect -3301 -45188 -3174 -45172
rect -3301 -45252 -3254 -45188
rect -3190 -45252 -3174 -45188
rect -3301 -45268 -3174 -45252
rect -3301 -45332 -3254 -45268
rect -3190 -45332 -3174 -45268
rect -3301 -45348 -3174 -45332
rect -3301 -45412 -3254 -45348
rect -3190 -45412 -3174 -45348
rect -3301 -45428 -3174 -45412
rect -3301 -45492 -3254 -45428
rect -3190 -45492 -3174 -45428
rect -3301 -45508 -3174 -45492
rect -3301 -45572 -3254 -45508
rect -3190 -45572 -3174 -45508
rect -3301 -45588 -3174 -45572
rect -3301 -45652 -3254 -45588
rect -3190 -45652 -3174 -45588
rect -3301 -45668 -3174 -45652
rect -3301 -45732 -3254 -45668
rect -3190 -45732 -3174 -45668
rect -3301 -45748 -3174 -45732
rect -3301 -45812 -3254 -45748
rect -3190 -45812 -3174 -45748
rect -3301 -45828 -3174 -45812
rect -3301 -45892 -3254 -45828
rect -3190 -45892 -3174 -45828
rect -3301 -45908 -3174 -45892
rect -3301 -45972 -3254 -45908
rect -3190 -45972 -3174 -45908
rect -3301 -45988 -3174 -45972
rect -3301 -46052 -3254 -45988
rect -3190 -46052 -3174 -45988
rect -3301 -46068 -3174 -46052
rect -3301 -46132 -3254 -46068
rect -3190 -46132 -3174 -46068
rect -3301 -46148 -3174 -46132
rect -3301 -46212 -3254 -46148
rect -3190 -46212 -3174 -46148
rect -3301 -46228 -3174 -46212
rect -3301 -46292 -3254 -46228
rect -3190 -46292 -3174 -46228
rect -3301 -46308 -3174 -46292
rect -3301 -46372 -3254 -46308
rect -3190 -46372 -3174 -46308
rect -3301 -46388 -3174 -46372
rect -3301 -46452 -3254 -46388
rect -3190 -46452 -3174 -46388
rect -3301 -46468 -3174 -46452
rect -3301 -46532 -3254 -46468
rect -3190 -46532 -3174 -46468
rect -3301 -46548 -3174 -46532
rect -3301 -46612 -3254 -46548
rect -3190 -46612 -3174 -46548
rect -3301 -46628 -3174 -46612
rect -3301 -46692 -3254 -46628
rect -3190 -46692 -3174 -46628
rect -3301 -46708 -3174 -46692
rect -3301 -46772 -3254 -46708
rect -3190 -46772 -3174 -46708
rect -3301 -46788 -3174 -46772
rect -3301 -46852 -3254 -46788
rect -3190 -46852 -3174 -46788
rect -3301 -46868 -3174 -46852
rect -3301 -46932 -3254 -46868
rect -3190 -46932 -3174 -46868
rect -3301 -46948 -3174 -46932
rect -3301 -47012 -3254 -46948
rect -3190 -47012 -3174 -46948
rect -3301 -47028 -3174 -47012
rect -9620 -47108 -9493 -47092
rect -9620 -47172 -9573 -47108
rect -9509 -47172 -9493 -47108
rect -9620 -47188 -9493 -47172
rect -9620 -47250 -9516 -47188
rect -6421 -47250 -6317 -47061
rect -3301 -47092 -3254 -47028
rect -3190 -47092 -3174 -47028
rect -3011 -41148 2911 -41139
rect -3011 -47052 -3002 -41148
rect 2902 -47052 2911 -41148
rect -3011 -47061 2911 -47052
rect 3018 -41172 3065 -41108
rect 3129 -41172 3145 -41108
rect 6217 -41139 6321 -40761
rect 9337 -40792 9384 -40728
rect 9448 -40792 9464 -40728
rect 9627 -34848 15549 -34839
rect 9627 -40752 9636 -34848
rect 15540 -40752 15549 -34848
rect 9627 -40761 15549 -40752
rect 15656 -34872 15703 -34808
rect 15767 -34872 15783 -34808
rect 18855 -34839 18959 -34461
rect 21975 -34492 22022 -34428
rect 22086 -34492 22102 -34428
rect 22265 -28548 28187 -28539
rect 22265 -34452 22274 -28548
rect 28178 -34452 28187 -28548
rect 22265 -34461 28187 -34452
rect 28294 -28572 28341 -28508
rect 28405 -28572 28421 -28508
rect 31493 -28539 31597 -28161
rect 34613 -28192 34660 -28128
rect 34724 -28192 34740 -28128
rect 34903 -22248 40825 -22239
rect 34903 -28152 34912 -22248
rect 40816 -28152 40825 -22248
rect 34903 -28161 40825 -28152
rect 40932 -22272 40979 -22208
rect 41043 -22272 41059 -22208
rect 44131 -22239 44235 -21861
rect 47251 -21892 47298 -21828
rect 47362 -21892 47378 -21828
rect 47251 -21908 47378 -21892
rect 47251 -21972 47298 -21908
rect 47362 -21972 47378 -21908
rect 47251 -21988 47378 -21972
rect 47251 -22112 47355 -21988
rect 47251 -22128 47378 -22112
rect 47251 -22192 47298 -22128
rect 47362 -22192 47378 -22128
rect 47251 -22208 47378 -22192
rect 40932 -22288 41059 -22272
rect 40932 -22352 40979 -22288
rect 41043 -22352 41059 -22288
rect 40932 -22368 41059 -22352
rect 40932 -22432 40979 -22368
rect 41043 -22432 41059 -22368
rect 40932 -22448 41059 -22432
rect 40932 -22512 40979 -22448
rect 41043 -22512 41059 -22448
rect 40932 -22528 41059 -22512
rect 40932 -22592 40979 -22528
rect 41043 -22592 41059 -22528
rect 40932 -22608 41059 -22592
rect 40932 -22672 40979 -22608
rect 41043 -22672 41059 -22608
rect 40932 -22688 41059 -22672
rect 40932 -22752 40979 -22688
rect 41043 -22752 41059 -22688
rect 40932 -22768 41059 -22752
rect 40932 -22832 40979 -22768
rect 41043 -22832 41059 -22768
rect 40932 -22848 41059 -22832
rect 40932 -22912 40979 -22848
rect 41043 -22912 41059 -22848
rect 40932 -22928 41059 -22912
rect 40932 -22992 40979 -22928
rect 41043 -22992 41059 -22928
rect 40932 -23008 41059 -22992
rect 40932 -23072 40979 -23008
rect 41043 -23072 41059 -23008
rect 40932 -23088 41059 -23072
rect 40932 -23152 40979 -23088
rect 41043 -23152 41059 -23088
rect 40932 -23168 41059 -23152
rect 40932 -23232 40979 -23168
rect 41043 -23232 41059 -23168
rect 40932 -23248 41059 -23232
rect 40932 -23312 40979 -23248
rect 41043 -23312 41059 -23248
rect 40932 -23328 41059 -23312
rect 40932 -23392 40979 -23328
rect 41043 -23392 41059 -23328
rect 40932 -23408 41059 -23392
rect 40932 -23472 40979 -23408
rect 41043 -23472 41059 -23408
rect 40932 -23488 41059 -23472
rect 40932 -23552 40979 -23488
rect 41043 -23552 41059 -23488
rect 40932 -23568 41059 -23552
rect 40932 -23632 40979 -23568
rect 41043 -23632 41059 -23568
rect 40932 -23648 41059 -23632
rect 40932 -23712 40979 -23648
rect 41043 -23712 41059 -23648
rect 40932 -23728 41059 -23712
rect 40932 -23792 40979 -23728
rect 41043 -23792 41059 -23728
rect 40932 -23808 41059 -23792
rect 40932 -23872 40979 -23808
rect 41043 -23872 41059 -23808
rect 40932 -23888 41059 -23872
rect 40932 -23952 40979 -23888
rect 41043 -23952 41059 -23888
rect 40932 -23968 41059 -23952
rect 40932 -24032 40979 -23968
rect 41043 -24032 41059 -23968
rect 40932 -24048 41059 -24032
rect 40932 -24112 40979 -24048
rect 41043 -24112 41059 -24048
rect 40932 -24128 41059 -24112
rect 40932 -24192 40979 -24128
rect 41043 -24192 41059 -24128
rect 40932 -24208 41059 -24192
rect 40932 -24272 40979 -24208
rect 41043 -24272 41059 -24208
rect 40932 -24288 41059 -24272
rect 40932 -24352 40979 -24288
rect 41043 -24352 41059 -24288
rect 40932 -24368 41059 -24352
rect 40932 -24432 40979 -24368
rect 41043 -24432 41059 -24368
rect 40932 -24448 41059 -24432
rect 40932 -24512 40979 -24448
rect 41043 -24512 41059 -24448
rect 40932 -24528 41059 -24512
rect 40932 -24592 40979 -24528
rect 41043 -24592 41059 -24528
rect 40932 -24608 41059 -24592
rect 40932 -24672 40979 -24608
rect 41043 -24672 41059 -24608
rect 40932 -24688 41059 -24672
rect 40932 -24752 40979 -24688
rect 41043 -24752 41059 -24688
rect 40932 -24768 41059 -24752
rect 40932 -24832 40979 -24768
rect 41043 -24832 41059 -24768
rect 40932 -24848 41059 -24832
rect 40932 -24912 40979 -24848
rect 41043 -24912 41059 -24848
rect 40932 -24928 41059 -24912
rect 40932 -24992 40979 -24928
rect 41043 -24992 41059 -24928
rect 40932 -25008 41059 -24992
rect 40932 -25072 40979 -25008
rect 41043 -25072 41059 -25008
rect 40932 -25088 41059 -25072
rect 40932 -25152 40979 -25088
rect 41043 -25152 41059 -25088
rect 40932 -25168 41059 -25152
rect 40932 -25232 40979 -25168
rect 41043 -25232 41059 -25168
rect 40932 -25248 41059 -25232
rect 40932 -25312 40979 -25248
rect 41043 -25312 41059 -25248
rect 40932 -25328 41059 -25312
rect 40932 -25392 40979 -25328
rect 41043 -25392 41059 -25328
rect 40932 -25408 41059 -25392
rect 40932 -25472 40979 -25408
rect 41043 -25472 41059 -25408
rect 40932 -25488 41059 -25472
rect 40932 -25552 40979 -25488
rect 41043 -25552 41059 -25488
rect 40932 -25568 41059 -25552
rect 40932 -25632 40979 -25568
rect 41043 -25632 41059 -25568
rect 40932 -25648 41059 -25632
rect 40932 -25712 40979 -25648
rect 41043 -25712 41059 -25648
rect 40932 -25728 41059 -25712
rect 40932 -25792 40979 -25728
rect 41043 -25792 41059 -25728
rect 40932 -25808 41059 -25792
rect 40932 -25872 40979 -25808
rect 41043 -25872 41059 -25808
rect 40932 -25888 41059 -25872
rect 40932 -25952 40979 -25888
rect 41043 -25952 41059 -25888
rect 40932 -25968 41059 -25952
rect 40932 -26032 40979 -25968
rect 41043 -26032 41059 -25968
rect 40932 -26048 41059 -26032
rect 40932 -26112 40979 -26048
rect 41043 -26112 41059 -26048
rect 40932 -26128 41059 -26112
rect 40932 -26192 40979 -26128
rect 41043 -26192 41059 -26128
rect 40932 -26208 41059 -26192
rect 40932 -26272 40979 -26208
rect 41043 -26272 41059 -26208
rect 40932 -26288 41059 -26272
rect 40932 -26352 40979 -26288
rect 41043 -26352 41059 -26288
rect 40932 -26368 41059 -26352
rect 40932 -26432 40979 -26368
rect 41043 -26432 41059 -26368
rect 40932 -26448 41059 -26432
rect 40932 -26512 40979 -26448
rect 41043 -26512 41059 -26448
rect 40932 -26528 41059 -26512
rect 40932 -26592 40979 -26528
rect 41043 -26592 41059 -26528
rect 40932 -26608 41059 -26592
rect 40932 -26672 40979 -26608
rect 41043 -26672 41059 -26608
rect 40932 -26688 41059 -26672
rect 40932 -26752 40979 -26688
rect 41043 -26752 41059 -26688
rect 40932 -26768 41059 -26752
rect 40932 -26832 40979 -26768
rect 41043 -26832 41059 -26768
rect 40932 -26848 41059 -26832
rect 40932 -26912 40979 -26848
rect 41043 -26912 41059 -26848
rect 40932 -26928 41059 -26912
rect 40932 -26992 40979 -26928
rect 41043 -26992 41059 -26928
rect 40932 -27008 41059 -26992
rect 40932 -27072 40979 -27008
rect 41043 -27072 41059 -27008
rect 40932 -27088 41059 -27072
rect 40932 -27152 40979 -27088
rect 41043 -27152 41059 -27088
rect 40932 -27168 41059 -27152
rect 40932 -27232 40979 -27168
rect 41043 -27232 41059 -27168
rect 40932 -27248 41059 -27232
rect 40932 -27312 40979 -27248
rect 41043 -27312 41059 -27248
rect 40932 -27328 41059 -27312
rect 40932 -27392 40979 -27328
rect 41043 -27392 41059 -27328
rect 40932 -27408 41059 -27392
rect 40932 -27472 40979 -27408
rect 41043 -27472 41059 -27408
rect 40932 -27488 41059 -27472
rect 40932 -27552 40979 -27488
rect 41043 -27552 41059 -27488
rect 40932 -27568 41059 -27552
rect 40932 -27632 40979 -27568
rect 41043 -27632 41059 -27568
rect 40932 -27648 41059 -27632
rect 40932 -27712 40979 -27648
rect 41043 -27712 41059 -27648
rect 40932 -27728 41059 -27712
rect 40932 -27792 40979 -27728
rect 41043 -27792 41059 -27728
rect 40932 -27808 41059 -27792
rect 40932 -27872 40979 -27808
rect 41043 -27872 41059 -27808
rect 40932 -27888 41059 -27872
rect 40932 -27952 40979 -27888
rect 41043 -27952 41059 -27888
rect 40932 -27968 41059 -27952
rect 40932 -28032 40979 -27968
rect 41043 -28032 41059 -27968
rect 40932 -28048 41059 -28032
rect 40932 -28112 40979 -28048
rect 41043 -28112 41059 -28048
rect 40932 -28128 41059 -28112
rect 34613 -28208 34740 -28192
rect 34613 -28272 34660 -28208
rect 34724 -28272 34740 -28208
rect 34613 -28288 34740 -28272
rect 34613 -28412 34717 -28288
rect 34613 -28428 34740 -28412
rect 34613 -28492 34660 -28428
rect 34724 -28492 34740 -28428
rect 34613 -28508 34740 -28492
rect 28294 -28588 28421 -28572
rect 28294 -28652 28341 -28588
rect 28405 -28652 28421 -28588
rect 28294 -28668 28421 -28652
rect 28294 -28732 28341 -28668
rect 28405 -28732 28421 -28668
rect 28294 -28748 28421 -28732
rect 28294 -28812 28341 -28748
rect 28405 -28812 28421 -28748
rect 28294 -28828 28421 -28812
rect 28294 -28892 28341 -28828
rect 28405 -28892 28421 -28828
rect 28294 -28908 28421 -28892
rect 28294 -28972 28341 -28908
rect 28405 -28972 28421 -28908
rect 28294 -28988 28421 -28972
rect 28294 -29052 28341 -28988
rect 28405 -29052 28421 -28988
rect 28294 -29068 28421 -29052
rect 28294 -29132 28341 -29068
rect 28405 -29132 28421 -29068
rect 28294 -29148 28421 -29132
rect 28294 -29212 28341 -29148
rect 28405 -29212 28421 -29148
rect 28294 -29228 28421 -29212
rect 28294 -29292 28341 -29228
rect 28405 -29292 28421 -29228
rect 28294 -29308 28421 -29292
rect 28294 -29372 28341 -29308
rect 28405 -29372 28421 -29308
rect 28294 -29388 28421 -29372
rect 28294 -29452 28341 -29388
rect 28405 -29452 28421 -29388
rect 28294 -29468 28421 -29452
rect 28294 -29532 28341 -29468
rect 28405 -29532 28421 -29468
rect 28294 -29548 28421 -29532
rect 28294 -29612 28341 -29548
rect 28405 -29612 28421 -29548
rect 28294 -29628 28421 -29612
rect 28294 -29692 28341 -29628
rect 28405 -29692 28421 -29628
rect 28294 -29708 28421 -29692
rect 28294 -29772 28341 -29708
rect 28405 -29772 28421 -29708
rect 28294 -29788 28421 -29772
rect 28294 -29852 28341 -29788
rect 28405 -29852 28421 -29788
rect 28294 -29868 28421 -29852
rect 28294 -29932 28341 -29868
rect 28405 -29932 28421 -29868
rect 28294 -29948 28421 -29932
rect 28294 -30012 28341 -29948
rect 28405 -30012 28421 -29948
rect 28294 -30028 28421 -30012
rect 28294 -30092 28341 -30028
rect 28405 -30092 28421 -30028
rect 28294 -30108 28421 -30092
rect 28294 -30172 28341 -30108
rect 28405 -30172 28421 -30108
rect 28294 -30188 28421 -30172
rect 28294 -30252 28341 -30188
rect 28405 -30252 28421 -30188
rect 28294 -30268 28421 -30252
rect 28294 -30332 28341 -30268
rect 28405 -30332 28421 -30268
rect 28294 -30348 28421 -30332
rect 28294 -30412 28341 -30348
rect 28405 -30412 28421 -30348
rect 28294 -30428 28421 -30412
rect 28294 -30492 28341 -30428
rect 28405 -30492 28421 -30428
rect 28294 -30508 28421 -30492
rect 28294 -30572 28341 -30508
rect 28405 -30572 28421 -30508
rect 28294 -30588 28421 -30572
rect 28294 -30652 28341 -30588
rect 28405 -30652 28421 -30588
rect 28294 -30668 28421 -30652
rect 28294 -30732 28341 -30668
rect 28405 -30732 28421 -30668
rect 28294 -30748 28421 -30732
rect 28294 -30812 28341 -30748
rect 28405 -30812 28421 -30748
rect 28294 -30828 28421 -30812
rect 28294 -30892 28341 -30828
rect 28405 -30892 28421 -30828
rect 28294 -30908 28421 -30892
rect 28294 -30972 28341 -30908
rect 28405 -30972 28421 -30908
rect 28294 -30988 28421 -30972
rect 28294 -31052 28341 -30988
rect 28405 -31052 28421 -30988
rect 28294 -31068 28421 -31052
rect 28294 -31132 28341 -31068
rect 28405 -31132 28421 -31068
rect 28294 -31148 28421 -31132
rect 28294 -31212 28341 -31148
rect 28405 -31212 28421 -31148
rect 28294 -31228 28421 -31212
rect 28294 -31292 28341 -31228
rect 28405 -31292 28421 -31228
rect 28294 -31308 28421 -31292
rect 28294 -31372 28341 -31308
rect 28405 -31372 28421 -31308
rect 28294 -31388 28421 -31372
rect 28294 -31452 28341 -31388
rect 28405 -31452 28421 -31388
rect 28294 -31468 28421 -31452
rect 28294 -31532 28341 -31468
rect 28405 -31532 28421 -31468
rect 28294 -31548 28421 -31532
rect 28294 -31612 28341 -31548
rect 28405 -31612 28421 -31548
rect 28294 -31628 28421 -31612
rect 28294 -31692 28341 -31628
rect 28405 -31692 28421 -31628
rect 28294 -31708 28421 -31692
rect 28294 -31772 28341 -31708
rect 28405 -31772 28421 -31708
rect 28294 -31788 28421 -31772
rect 28294 -31852 28341 -31788
rect 28405 -31852 28421 -31788
rect 28294 -31868 28421 -31852
rect 28294 -31932 28341 -31868
rect 28405 -31932 28421 -31868
rect 28294 -31948 28421 -31932
rect 28294 -32012 28341 -31948
rect 28405 -32012 28421 -31948
rect 28294 -32028 28421 -32012
rect 28294 -32092 28341 -32028
rect 28405 -32092 28421 -32028
rect 28294 -32108 28421 -32092
rect 28294 -32172 28341 -32108
rect 28405 -32172 28421 -32108
rect 28294 -32188 28421 -32172
rect 28294 -32252 28341 -32188
rect 28405 -32252 28421 -32188
rect 28294 -32268 28421 -32252
rect 28294 -32332 28341 -32268
rect 28405 -32332 28421 -32268
rect 28294 -32348 28421 -32332
rect 28294 -32412 28341 -32348
rect 28405 -32412 28421 -32348
rect 28294 -32428 28421 -32412
rect 28294 -32492 28341 -32428
rect 28405 -32492 28421 -32428
rect 28294 -32508 28421 -32492
rect 28294 -32572 28341 -32508
rect 28405 -32572 28421 -32508
rect 28294 -32588 28421 -32572
rect 28294 -32652 28341 -32588
rect 28405 -32652 28421 -32588
rect 28294 -32668 28421 -32652
rect 28294 -32732 28341 -32668
rect 28405 -32732 28421 -32668
rect 28294 -32748 28421 -32732
rect 28294 -32812 28341 -32748
rect 28405 -32812 28421 -32748
rect 28294 -32828 28421 -32812
rect 28294 -32892 28341 -32828
rect 28405 -32892 28421 -32828
rect 28294 -32908 28421 -32892
rect 28294 -32972 28341 -32908
rect 28405 -32972 28421 -32908
rect 28294 -32988 28421 -32972
rect 28294 -33052 28341 -32988
rect 28405 -33052 28421 -32988
rect 28294 -33068 28421 -33052
rect 28294 -33132 28341 -33068
rect 28405 -33132 28421 -33068
rect 28294 -33148 28421 -33132
rect 28294 -33212 28341 -33148
rect 28405 -33212 28421 -33148
rect 28294 -33228 28421 -33212
rect 28294 -33292 28341 -33228
rect 28405 -33292 28421 -33228
rect 28294 -33308 28421 -33292
rect 28294 -33372 28341 -33308
rect 28405 -33372 28421 -33308
rect 28294 -33388 28421 -33372
rect 28294 -33452 28341 -33388
rect 28405 -33452 28421 -33388
rect 28294 -33468 28421 -33452
rect 28294 -33532 28341 -33468
rect 28405 -33532 28421 -33468
rect 28294 -33548 28421 -33532
rect 28294 -33612 28341 -33548
rect 28405 -33612 28421 -33548
rect 28294 -33628 28421 -33612
rect 28294 -33692 28341 -33628
rect 28405 -33692 28421 -33628
rect 28294 -33708 28421 -33692
rect 28294 -33772 28341 -33708
rect 28405 -33772 28421 -33708
rect 28294 -33788 28421 -33772
rect 28294 -33852 28341 -33788
rect 28405 -33852 28421 -33788
rect 28294 -33868 28421 -33852
rect 28294 -33932 28341 -33868
rect 28405 -33932 28421 -33868
rect 28294 -33948 28421 -33932
rect 28294 -34012 28341 -33948
rect 28405 -34012 28421 -33948
rect 28294 -34028 28421 -34012
rect 28294 -34092 28341 -34028
rect 28405 -34092 28421 -34028
rect 28294 -34108 28421 -34092
rect 28294 -34172 28341 -34108
rect 28405 -34172 28421 -34108
rect 28294 -34188 28421 -34172
rect 28294 -34252 28341 -34188
rect 28405 -34252 28421 -34188
rect 28294 -34268 28421 -34252
rect 28294 -34332 28341 -34268
rect 28405 -34332 28421 -34268
rect 28294 -34348 28421 -34332
rect 28294 -34412 28341 -34348
rect 28405 -34412 28421 -34348
rect 28294 -34428 28421 -34412
rect 21975 -34508 22102 -34492
rect 21975 -34572 22022 -34508
rect 22086 -34572 22102 -34508
rect 21975 -34588 22102 -34572
rect 21975 -34712 22079 -34588
rect 21975 -34728 22102 -34712
rect 21975 -34792 22022 -34728
rect 22086 -34792 22102 -34728
rect 21975 -34808 22102 -34792
rect 15656 -34888 15783 -34872
rect 15656 -34952 15703 -34888
rect 15767 -34952 15783 -34888
rect 15656 -34968 15783 -34952
rect 15656 -35032 15703 -34968
rect 15767 -35032 15783 -34968
rect 15656 -35048 15783 -35032
rect 15656 -35112 15703 -35048
rect 15767 -35112 15783 -35048
rect 15656 -35128 15783 -35112
rect 15656 -35192 15703 -35128
rect 15767 -35192 15783 -35128
rect 15656 -35208 15783 -35192
rect 15656 -35272 15703 -35208
rect 15767 -35272 15783 -35208
rect 15656 -35288 15783 -35272
rect 15656 -35352 15703 -35288
rect 15767 -35352 15783 -35288
rect 15656 -35368 15783 -35352
rect 15656 -35432 15703 -35368
rect 15767 -35432 15783 -35368
rect 15656 -35448 15783 -35432
rect 15656 -35512 15703 -35448
rect 15767 -35512 15783 -35448
rect 15656 -35528 15783 -35512
rect 15656 -35592 15703 -35528
rect 15767 -35592 15783 -35528
rect 15656 -35608 15783 -35592
rect 15656 -35672 15703 -35608
rect 15767 -35672 15783 -35608
rect 15656 -35688 15783 -35672
rect 15656 -35752 15703 -35688
rect 15767 -35752 15783 -35688
rect 15656 -35768 15783 -35752
rect 15656 -35832 15703 -35768
rect 15767 -35832 15783 -35768
rect 15656 -35848 15783 -35832
rect 15656 -35912 15703 -35848
rect 15767 -35912 15783 -35848
rect 15656 -35928 15783 -35912
rect 15656 -35992 15703 -35928
rect 15767 -35992 15783 -35928
rect 15656 -36008 15783 -35992
rect 15656 -36072 15703 -36008
rect 15767 -36072 15783 -36008
rect 15656 -36088 15783 -36072
rect 15656 -36152 15703 -36088
rect 15767 -36152 15783 -36088
rect 15656 -36168 15783 -36152
rect 15656 -36232 15703 -36168
rect 15767 -36232 15783 -36168
rect 15656 -36248 15783 -36232
rect 15656 -36312 15703 -36248
rect 15767 -36312 15783 -36248
rect 15656 -36328 15783 -36312
rect 15656 -36392 15703 -36328
rect 15767 -36392 15783 -36328
rect 15656 -36408 15783 -36392
rect 15656 -36472 15703 -36408
rect 15767 -36472 15783 -36408
rect 15656 -36488 15783 -36472
rect 15656 -36552 15703 -36488
rect 15767 -36552 15783 -36488
rect 15656 -36568 15783 -36552
rect 15656 -36632 15703 -36568
rect 15767 -36632 15783 -36568
rect 15656 -36648 15783 -36632
rect 15656 -36712 15703 -36648
rect 15767 -36712 15783 -36648
rect 15656 -36728 15783 -36712
rect 15656 -36792 15703 -36728
rect 15767 -36792 15783 -36728
rect 15656 -36808 15783 -36792
rect 15656 -36872 15703 -36808
rect 15767 -36872 15783 -36808
rect 15656 -36888 15783 -36872
rect 15656 -36952 15703 -36888
rect 15767 -36952 15783 -36888
rect 15656 -36968 15783 -36952
rect 15656 -37032 15703 -36968
rect 15767 -37032 15783 -36968
rect 15656 -37048 15783 -37032
rect 15656 -37112 15703 -37048
rect 15767 -37112 15783 -37048
rect 15656 -37128 15783 -37112
rect 15656 -37192 15703 -37128
rect 15767 -37192 15783 -37128
rect 15656 -37208 15783 -37192
rect 15656 -37272 15703 -37208
rect 15767 -37272 15783 -37208
rect 15656 -37288 15783 -37272
rect 15656 -37352 15703 -37288
rect 15767 -37352 15783 -37288
rect 15656 -37368 15783 -37352
rect 15656 -37432 15703 -37368
rect 15767 -37432 15783 -37368
rect 15656 -37448 15783 -37432
rect 15656 -37512 15703 -37448
rect 15767 -37512 15783 -37448
rect 15656 -37528 15783 -37512
rect 15656 -37592 15703 -37528
rect 15767 -37592 15783 -37528
rect 15656 -37608 15783 -37592
rect 15656 -37672 15703 -37608
rect 15767 -37672 15783 -37608
rect 15656 -37688 15783 -37672
rect 15656 -37752 15703 -37688
rect 15767 -37752 15783 -37688
rect 15656 -37768 15783 -37752
rect 15656 -37832 15703 -37768
rect 15767 -37832 15783 -37768
rect 15656 -37848 15783 -37832
rect 15656 -37912 15703 -37848
rect 15767 -37912 15783 -37848
rect 15656 -37928 15783 -37912
rect 15656 -37992 15703 -37928
rect 15767 -37992 15783 -37928
rect 15656 -38008 15783 -37992
rect 15656 -38072 15703 -38008
rect 15767 -38072 15783 -38008
rect 15656 -38088 15783 -38072
rect 15656 -38152 15703 -38088
rect 15767 -38152 15783 -38088
rect 15656 -38168 15783 -38152
rect 15656 -38232 15703 -38168
rect 15767 -38232 15783 -38168
rect 15656 -38248 15783 -38232
rect 15656 -38312 15703 -38248
rect 15767 -38312 15783 -38248
rect 15656 -38328 15783 -38312
rect 15656 -38392 15703 -38328
rect 15767 -38392 15783 -38328
rect 15656 -38408 15783 -38392
rect 15656 -38472 15703 -38408
rect 15767 -38472 15783 -38408
rect 15656 -38488 15783 -38472
rect 15656 -38552 15703 -38488
rect 15767 -38552 15783 -38488
rect 15656 -38568 15783 -38552
rect 15656 -38632 15703 -38568
rect 15767 -38632 15783 -38568
rect 15656 -38648 15783 -38632
rect 15656 -38712 15703 -38648
rect 15767 -38712 15783 -38648
rect 15656 -38728 15783 -38712
rect 15656 -38792 15703 -38728
rect 15767 -38792 15783 -38728
rect 15656 -38808 15783 -38792
rect 15656 -38872 15703 -38808
rect 15767 -38872 15783 -38808
rect 15656 -38888 15783 -38872
rect 15656 -38952 15703 -38888
rect 15767 -38952 15783 -38888
rect 15656 -38968 15783 -38952
rect 15656 -39032 15703 -38968
rect 15767 -39032 15783 -38968
rect 15656 -39048 15783 -39032
rect 15656 -39112 15703 -39048
rect 15767 -39112 15783 -39048
rect 15656 -39128 15783 -39112
rect 15656 -39192 15703 -39128
rect 15767 -39192 15783 -39128
rect 15656 -39208 15783 -39192
rect 15656 -39272 15703 -39208
rect 15767 -39272 15783 -39208
rect 15656 -39288 15783 -39272
rect 15656 -39352 15703 -39288
rect 15767 -39352 15783 -39288
rect 15656 -39368 15783 -39352
rect 15656 -39432 15703 -39368
rect 15767 -39432 15783 -39368
rect 15656 -39448 15783 -39432
rect 15656 -39512 15703 -39448
rect 15767 -39512 15783 -39448
rect 15656 -39528 15783 -39512
rect 15656 -39592 15703 -39528
rect 15767 -39592 15783 -39528
rect 15656 -39608 15783 -39592
rect 15656 -39672 15703 -39608
rect 15767 -39672 15783 -39608
rect 15656 -39688 15783 -39672
rect 15656 -39752 15703 -39688
rect 15767 -39752 15783 -39688
rect 15656 -39768 15783 -39752
rect 15656 -39832 15703 -39768
rect 15767 -39832 15783 -39768
rect 15656 -39848 15783 -39832
rect 15656 -39912 15703 -39848
rect 15767 -39912 15783 -39848
rect 15656 -39928 15783 -39912
rect 15656 -39992 15703 -39928
rect 15767 -39992 15783 -39928
rect 15656 -40008 15783 -39992
rect 15656 -40072 15703 -40008
rect 15767 -40072 15783 -40008
rect 15656 -40088 15783 -40072
rect 15656 -40152 15703 -40088
rect 15767 -40152 15783 -40088
rect 15656 -40168 15783 -40152
rect 15656 -40232 15703 -40168
rect 15767 -40232 15783 -40168
rect 15656 -40248 15783 -40232
rect 15656 -40312 15703 -40248
rect 15767 -40312 15783 -40248
rect 15656 -40328 15783 -40312
rect 15656 -40392 15703 -40328
rect 15767 -40392 15783 -40328
rect 15656 -40408 15783 -40392
rect 15656 -40472 15703 -40408
rect 15767 -40472 15783 -40408
rect 15656 -40488 15783 -40472
rect 15656 -40552 15703 -40488
rect 15767 -40552 15783 -40488
rect 15656 -40568 15783 -40552
rect 15656 -40632 15703 -40568
rect 15767 -40632 15783 -40568
rect 15656 -40648 15783 -40632
rect 15656 -40712 15703 -40648
rect 15767 -40712 15783 -40648
rect 15656 -40728 15783 -40712
rect 9337 -40808 9464 -40792
rect 9337 -40872 9384 -40808
rect 9448 -40872 9464 -40808
rect 9337 -40888 9464 -40872
rect 9337 -41012 9441 -40888
rect 9337 -41028 9464 -41012
rect 9337 -41092 9384 -41028
rect 9448 -41092 9464 -41028
rect 9337 -41108 9464 -41092
rect 3018 -41188 3145 -41172
rect 3018 -41252 3065 -41188
rect 3129 -41252 3145 -41188
rect 3018 -41268 3145 -41252
rect 3018 -41332 3065 -41268
rect 3129 -41332 3145 -41268
rect 3018 -41348 3145 -41332
rect 3018 -41412 3065 -41348
rect 3129 -41412 3145 -41348
rect 3018 -41428 3145 -41412
rect 3018 -41492 3065 -41428
rect 3129 -41492 3145 -41428
rect 3018 -41508 3145 -41492
rect 3018 -41572 3065 -41508
rect 3129 -41572 3145 -41508
rect 3018 -41588 3145 -41572
rect 3018 -41652 3065 -41588
rect 3129 -41652 3145 -41588
rect 3018 -41668 3145 -41652
rect 3018 -41732 3065 -41668
rect 3129 -41732 3145 -41668
rect 3018 -41748 3145 -41732
rect 3018 -41812 3065 -41748
rect 3129 -41812 3145 -41748
rect 3018 -41828 3145 -41812
rect 3018 -41892 3065 -41828
rect 3129 -41892 3145 -41828
rect 3018 -41908 3145 -41892
rect 3018 -41972 3065 -41908
rect 3129 -41972 3145 -41908
rect 3018 -41988 3145 -41972
rect 3018 -42052 3065 -41988
rect 3129 -42052 3145 -41988
rect 3018 -42068 3145 -42052
rect 3018 -42132 3065 -42068
rect 3129 -42132 3145 -42068
rect 3018 -42148 3145 -42132
rect 3018 -42212 3065 -42148
rect 3129 -42212 3145 -42148
rect 3018 -42228 3145 -42212
rect 3018 -42292 3065 -42228
rect 3129 -42292 3145 -42228
rect 3018 -42308 3145 -42292
rect 3018 -42372 3065 -42308
rect 3129 -42372 3145 -42308
rect 3018 -42388 3145 -42372
rect 3018 -42452 3065 -42388
rect 3129 -42452 3145 -42388
rect 3018 -42468 3145 -42452
rect 3018 -42532 3065 -42468
rect 3129 -42532 3145 -42468
rect 3018 -42548 3145 -42532
rect 3018 -42612 3065 -42548
rect 3129 -42612 3145 -42548
rect 3018 -42628 3145 -42612
rect 3018 -42692 3065 -42628
rect 3129 -42692 3145 -42628
rect 3018 -42708 3145 -42692
rect 3018 -42772 3065 -42708
rect 3129 -42772 3145 -42708
rect 3018 -42788 3145 -42772
rect 3018 -42852 3065 -42788
rect 3129 -42852 3145 -42788
rect 3018 -42868 3145 -42852
rect 3018 -42932 3065 -42868
rect 3129 -42932 3145 -42868
rect 3018 -42948 3145 -42932
rect 3018 -43012 3065 -42948
rect 3129 -43012 3145 -42948
rect 3018 -43028 3145 -43012
rect 3018 -43092 3065 -43028
rect 3129 -43092 3145 -43028
rect 3018 -43108 3145 -43092
rect 3018 -43172 3065 -43108
rect 3129 -43172 3145 -43108
rect 3018 -43188 3145 -43172
rect 3018 -43252 3065 -43188
rect 3129 -43252 3145 -43188
rect 3018 -43268 3145 -43252
rect 3018 -43332 3065 -43268
rect 3129 -43332 3145 -43268
rect 3018 -43348 3145 -43332
rect 3018 -43412 3065 -43348
rect 3129 -43412 3145 -43348
rect 3018 -43428 3145 -43412
rect 3018 -43492 3065 -43428
rect 3129 -43492 3145 -43428
rect 3018 -43508 3145 -43492
rect 3018 -43572 3065 -43508
rect 3129 -43572 3145 -43508
rect 3018 -43588 3145 -43572
rect 3018 -43652 3065 -43588
rect 3129 -43652 3145 -43588
rect 3018 -43668 3145 -43652
rect 3018 -43732 3065 -43668
rect 3129 -43732 3145 -43668
rect 3018 -43748 3145 -43732
rect 3018 -43812 3065 -43748
rect 3129 -43812 3145 -43748
rect 3018 -43828 3145 -43812
rect 3018 -43892 3065 -43828
rect 3129 -43892 3145 -43828
rect 3018 -43908 3145 -43892
rect 3018 -43972 3065 -43908
rect 3129 -43972 3145 -43908
rect 3018 -43988 3145 -43972
rect 3018 -44052 3065 -43988
rect 3129 -44052 3145 -43988
rect 3018 -44068 3145 -44052
rect 3018 -44132 3065 -44068
rect 3129 -44132 3145 -44068
rect 3018 -44148 3145 -44132
rect 3018 -44212 3065 -44148
rect 3129 -44212 3145 -44148
rect 3018 -44228 3145 -44212
rect 3018 -44292 3065 -44228
rect 3129 -44292 3145 -44228
rect 3018 -44308 3145 -44292
rect 3018 -44372 3065 -44308
rect 3129 -44372 3145 -44308
rect 3018 -44388 3145 -44372
rect 3018 -44452 3065 -44388
rect 3129 -44452 3145 -44388
rect 3018 -44468 3145 -44452
rect 3018 -44532 3065 -44468
rect 3129 -44532 3145 -44468
rect 3018 -44548 3145 -44532
rect 3018 -44612 3065 -44548
rect 3129 -44612 3145 -44548
rect 3018 -44628 3145 -44612
rect 3018 -44692 3065 -44628
rect 3129 -44692 3145 -44628
rect 3018 -44708 3145 -44692
rect 3018 -44772 3065 -44708
rect 3129 -44772 3145 -44708
rect 3018 -44788 3145 -44772
rect 3018 -44852 3065 -44788
rect 3129 -44852 3145 -44788
rect 3018 -44868 3145 -44852
rect 3018 -44932 3065 -44868
rect 3129 -44932 3145 -44868
rect 3018 -44948 3145 -44932
rect 3018 -45012 3065 -44948
rect 3129 -45012 3145 -44948
rect 3018 -45028 3145 -45012
rect 3018 -45092 3065 -45028
rect 3129 -45092 3145 -45028
rect 3018 -45108 3145 -45092
rect 3018 -45172 3065 -45108
rect 3129 -45172 3145 -45108
rect 3018 -45188 3145 -45172
rect 3018 -45252 3065 -45188
rect 3129 -45252 3145 -45188
rect 3018 -45268 3145 -45252
rect 3018 -45332 3065 -45268
rect 3129 -45332 3145 -45268
rect 3018 -45348 3145 -45332
rect 3018 -45412 3065 -45348
rect 3129 -45412 3145 -45348
rect 3018 -45428 3145 -45412
rect 3018 -45492 3065 -45428
rect 3129 -45492 3145 -45428
rect 3018 -45508 3145 -45492
rect 3018 -45572 3065 -45508
rect 3129 -45572 3145 -45508
rect 3018 -45588 3145 -45572
rect 3018 -45652 3065 -45588
rect 3129 -45652 3145 -45588
rect 3018 -45668 3145 -45652
rect 3018 -45732 3065 -45668
rect 3129 -45732 3145 -45668
rect 3018 -45748 3145 -45732
rect 3018 -45812 3065 -45748
rect 3129 -45812 3145 -45748
rect 3018 -45828 3145 -45812
rect 3018 -45892 3065 -45828
rect 3129 -45892 3145 -45828
rect 3018 -45908 3145 -45892
rect 3018 -45972 3065 -45908
rect 3129 -45972 3145 -45908
rect 3018 -45988 3145 -45972
rect 3018 -46052 3065 -45988
rect 3129 -46052 3145 -45988
rect 3018 -46068 3145 -46052
rect 3018 -46132 3065 -46068
rect 3129 -46132 3145 -46068
rect 3018 -46148 3145 -46132
rect 3018 -46212 3065 -46148
rect 3129 -46212 3145 -46148
rect 3018 -46228 3145 -46212
rect 3018 -46292 3065 -46228
rect 3129 -46292 3145 -46228
rect 3018 -46308 3145 -46292
rect 3018 -46372 3065 -46308
rect 3129 -46372 3145 -46308
rect 3018 -46388 3145 -46372
rect 3018 -46452 3065 -46388
rect 3129 -46452 3145 -46388
rect 3018 -46468 3145 -46452
rect 3018 -46532 3065 -46468
rect 3129 -46532 3145 -46468
rect 3018 -46548 3145 -46532
rect 3018 -46612 3065 -46548
rect 3129 -46612 3145 -46548
rect 3018 -46628 3145 -46612
rect 3018 -46692 3065 -46628
rect 3129 -46692 3145 -46628
rect 3018 -46708 3145 -46692
rect 3018 -46772 3065 -46708
rect 3129 -46772 3145 -46708
rect 3018 -46788 3145 -46772
rect 3018 -46852 3065 -46788
rect 3129 -46852 3145 -46788
rect 3018 -46868 3145 -46852
rect 3018 -46932 3065 -46868
rect 3129 -46932 3145 -46868
rect 3018 -46948 3145 -46932
rect 3018 -47012 3065 -46948
rect 3129 -47012 3145 -46948
rect 3018 -47028 3145 -47012
rect -3301 -47108 -3174 -47092
rect -3301 -47172 -3254 -47108
rect -3190 -47172 -3174 -47108
rect -3301 -47188 -3174 -47172
rect -3301 -47250 -3197 -47188
rect -102 -47250 2 -47061
rect 3018 -47092 3065 -47028
rect 3129 -47092 3145 -47028
rect 3308 -41148 9230 -41139
rect 3308 -47052 3317 -41148
rect 9221 -47052 9230 -41148
rect 3308 -47061 9230 -47052
rect 9337 -41172 9384 -41108
rect 9448 -41172 9464 -41108
rect 12536 -41139 12640 -40761
rect 15656 -40792 15703 -40728
rect 15767 -40792 15783 -40728
rect 15946 -34848 21868 -34839
rect 15946 -40752 15955 -34848
rect 21859 -40752 21868 -34848
rect 15946 -40761 21868 -40752
rect 21975 -34872 22022 -34808
rect 22086 -34872 22102 -34808
rect 25174 -34839 25278 -34461
rect 28294 -34492 28341 -34428
rect 28405 -34492 28421 -34428
rect 28584 -28548 34506 -28539
rect 28584 -34452 28593 -28548
rect 34497 -34452 34506 -28548
rect 28584 -34461 34506 -34452
rect 34613 -28572 34660 -28508
rect 34724 -28572 34740 -28508
rect 37812 -28539 37916 -28161
rect 40932 -28192 40979 -28128
rect 41043 -28192 41059 -28128
rect 41222 -22248 47144 -22239
rect 41222 -28152 41231 -22248
rect 47135 -28152 47144 -22248
rect 41222 -28161 47144 -28152
rect 47251 -22272 47298 -22208
rect 47362 -22272 47378 -22208
rect 47251 -22288 47378 -22272
rect 47251 -22352 47298 -22288
rect 47362 -22352 47378 -22288
rect 47251 -22368 47378 -22352
rect 47251 -22432 47298 -22368
rect 47362 -22432 47378 -22368
rect 47251 -22448 47378 -22432
rect 47251 -22512 47298 -22448
rect 47362 -22512 47378 -22448
rect 47251 -22528 47378 -22512
rect 47251 -22592 47298 -22528
rect 47362 -22592 47378 -22528
rect 47251 -22608 47378 -22592
rect 47251 -22672 47298 -22608
rect 47362 -22672 47378 -22608
rect 47251 -22688 47378 -22672
rect 47251 -22752 47298 -22688
rect 47362 -22752 47378 -22688
rect 47251 -22768 47378 -22752
rect 47251 -22832 47298 -22768
rect 47362 -22832 47378 -22768
rect 47251 -22848 47378 -22832
rect 47251 -22912 47298 -22848
rect 47362 -22912 47378 -22848
rect 47251 -22928 47378 -22912
rect 47251 -22992 47298 -22928
rect 47362 -22992 47378 -22928
rect 47251 -23008 47378 -22992
rect 47251 -23072 47298 -23008
rect 47362 -23072 47378 -23008
rect 47251 -23088 47378 -23072
rect 47251 -23152 47298 -23088
rect 47362 -23152 47378 -23088
rect 47251 -23168 47378 -23152
rect 47251 -23232 47298 -23168
rect 47362 -23232 47378 -23168
rect 47251 -23248 47378 -23232
rect 47251 -23312 47298 -23248
rect 47362 -23312 47378 -23248
rect 47251 -23328 47378 -23312
rect 47251 -23392 47298 -23328
rect 47362 -23392 47378 -23328
rect 47251 -23408 47378 -23392
rect 47251 -23472 47298 -23408
rect 47362 -23472 47378 -23408
rect 47251 -23488 47378 -23472
rect 47251 -23552 47298 -23488
rect 47362 -23552 47378 -23488
rect 47251 -23568 47378 -23552
rect 47251 -23632 47298 -23568
rect 47362 -23632 47378 -23568
rect 47251 -23648 47378 -23632
rect 47251 -23712 47298 -23648
rect 47362 -23712 47378 -23648
rect 47251 -23728 47378 -23712
rect 47251 -23792 47298 -23728
rect 47362 -23792 47378 -23728
rect 47251 -23808 47378 -23792
rect 47251 -23872 47298 -23808
rect 47362 -23872 47378 -23808
rect 47251 -23888 47378 -23872
rect 47251 -23952 47298 -23888
rect 47362 -23952 47378 -23888
rect 47251 -23968 47378 -23952
rect 47251 -24032 47298 -23968
rect 47362 -24032 47378 -23968
rect 47251 -24048 47378 -24032
rect 47251 -24112 47298 -24048
rect 47362 -24112 47378 -24048
rect 47251 -24128 47378 -24112
rect 47251 -24192 47298 -24128
rect 47362 -24192 47378 -24128
rect 47251 -24208 47378 -24192
rect 47251 -24272 47298 -24208
rect 47362 -24272 47378 -24208
rect 47251 -24288 47378 -24272
rect 47251 -24352 47298 -24288
rect 47362 -24352 47378 -24288
rect 47251 -24368 47378 -24352
rect 47251 -24432 47298 -24368
rect 47362 -24432 47378 -24368
rect 47251 -24448 47378 -24432
rect 47251 -24512 47298 -24448
rect 47362 -24512 47378 -24448
rect 47251 -24528 47378 -24512
rect 47251 -24592 47298 -24528
rect 47362 -24592 47378 -24528
rect 47251 -24608 47378 -24592
rect 47251 -24672 47298 -24608
rect 47362 -24672 47378 -24608
rect 47251 -24688 47378 -24672
rect 47251 -24752 47298 -24688
rect 47362 -24752 47378 -24688
rect 47251 -24768 47378 -24752
rect 47251 -24832 47298 -24768
rect 47362 -24832 47378 -24768
rect 47251 -24848 47378 -24832
rect 47251 -24912 47298 -24848
rect 47362 -24912 47378 -24848
rect 47251 -24928 47378 -24912
rect 47251 -24992 47298 -24928
rect 47362 -24992 47378 -24928
rect 47251 -25008 47378 -24992
rect 47251 -25072 47298 -25008
rect 47362 -25072 47378 -25008
rect 47251 -25088 47378 -25072
rect 47251 -25152 47298 -25088
rect 47362 -25152 47378 -25088
rect 47251 -25168 47378 -25152
rect 47251 -25232 47298 -25168
rect 47362 -25232 47378 -25168
rect 47251 -25248 47378 -25232
rect 47251 -25312 47298 -25248
rect 47362 -25312 47378 -25248
rect 47251 -25328 47378 -25312
rect 47251 -25392 47298 -25328
rect 47362 -25392 47378 -25328
rect 47251 -25408 47378 -25392
rect 47251 -25472 47298 -25408
rect 47362 -25472 47378 -25408
rect 47251 -25488 47378 -25472
rect 47251 -25552 47298 -25488
rect 47362 -25552 47378 -25488
rect 47251 -25568 47378 -25552
rect 47251 -25632 47298 -25568
rect 47362 -25632 47378 -25568
rect 47251 -25648 47378 -25632
rect 47251 -25712 47298 -25648
rect 47362 -25712 47378 -25648
rect 47251 -25728 47378 -25712
rect 47251 -25792 47298 -25728
rect 47362 -25792 47378 -25728
rect 47251 -25808 47378 -25792
rect 47251 -25872 47298 -25808
rect 47362 -25872 47378 -25808
rect 47251 -25888 47378 -25872
rect 47251 -25952 47298 -25888
rect 47362 -25952 47378 -25888
rect 47251 -25968 47378 -25952
rect 47251 -26032 47298 -25968
rect 47362 -26032 47378 -25968
rect 47251 -26048 47378 -26032
rect 47251 -26112 47298 -26048
rect 47362 -26112 47378 -26048
rect 47251 -26128 47378 -26112
rect 47251 -26192 47298 -26128
rect 47362 -26192 47378 -26128
rect 47251 -26208 47378 -26192
rect 47251 -26272 47298 -26208
rect 47362 -26272 47378 -26208
rect 47251 -26288 47378 -26272
rect 47251 -26352 47298 -26288
rect 47362 -26352 47378 -26288
rect 47251 -26368 47378 -26352
rect 47251 -26432 47298 -26368
rect 47362 -26432 47378 -26368
rect 47251 -26448 47378 -26432
rect 47251 -26512 47298 -26448
rect 47362 -26512 47378 -26448
rect 47251 -26528 47378 -26512
rect 47251 -26592 47298 -26528
rect 47362 -26592 47378 -26528
rect 47251 -26608 47378 -26592
rect 47251 -26672 47298 -26608
rect 47362 -26672 47378 -26608
rect 47251 -26688 47378 -26672
rect 47251 -26752 47298 -26688
rect 47362 -26752 47378 -26688
rect 47251 -26768 47378 -26752
rect 47251 -26832 47298 -26768
rect 47362 -26832 47378 -26768
rect 47251 -26848 47378 -26832
rect 47251 -26912 47298 -26848
rect 47362 -26912 47378 -26848
rect 47251 -26928 47378 -26912
rect 47251 -26992 47298 -26928
rect 47362 -26992 47378 -26928
rect 47251 -27008 47378 -26992
rect 47251 -27072 47298 -27008
rect 47362 -27072 47378 -27008
rect 47251 -27088 47378 -27072
rect 47251 -27152 47298 -27088
rect 47362 -27152 47378 -27088
rect 47251 -27168 47378 -27152
rect 47251 -27232 47298 -27168
rect 47362 -27232 47378 -27168
rect 47251 -27248 47378 -27232
rect 47251 -27312 47298 -27248
rect 47362 -27312 47378 -27248
rect 47251 -27328 47378 -27312
rect 47251 -27392 47298 -27328
rect 47362 -27392 47378 -27328
rect 47251 -27408 47378 -27392
rect 47251 -27472 47298 -27408
rect 47362 -27472 47378 -27408
rect 47251 -27488 47378 -27472
rect 47251 -27552 47298 -27488
rect 47362 -27552 47378 -27488
rect 47251 -27568 47378 -27552
rect 47251 -27632 47298 -27568
rect 47362 -27632 47378 -27568
rect 47251 -27648 47378 -27632
rect 47251 -27712 47298 -27648
rect 47362 -27712 47378 -27648
rect 47251 -27728 47378 -27712
rect 47251 -27792 47298 -27728
rect 47362 -27792 47378 -27728
rect 47251 -27808 47378 -27792
rect 47251 -27872 47298 -27808
rect 47362 -27872 47378 -27808
rect 47251 -27888 47378 -27872
rect 47251 -27952 47298 -27888
rect 47362 -27952 47378 -27888
rect 47251 -27968 47378 -27952
rect 47251 -28032 47298 -27968
rect 47362 -28032 47378 -27968
rect 47251 -28048 47378 -28032
rect 47251 -28112 47298 -28048
rect 47362 -28112 47378 -28048
rect 47251 -28128 47378 -28112
rect 40932 -28208 41059 -28192
rect 40932 -28272 40979 -28208
rect 41043 -28272 41059 -28208
rect 40932 -28288 41059 -28272
rect 40932 -28412 41036 -28288
rect 40932 -28428 41059 -28412
rect 40932 -28492 40979 -28428
rect 41043 -28492 41059 -28428
rect 40932 -28508 41059 -28492
rect 34613 -28588 34740 -28572
rect 34613 -28652 34660 -28588
rect 34724 -28652 34740 -28588
rect 34613 -28668 34740 -28652
rect 34613 -28732 34660 -28668
rect 34724 -28732 34740 -28668
rect 34613 -28748 34740 -28732
rect 34613 -28812 34660 -28748
rect 34724 -28812 34740 -28748
rect 34613 -28828 34740 -28812
rect 34613 -28892 34660 -28828
rect 34724 -28892 34740 -28828
rect 34613 -28908 34740 -28892
rect 34613 -28972 34660 -28908
rect 34724 -28972 34740 -28908
rect 34613 -28988 34740 -28972
rect 34613 -29052 34660 -28988
rect 34724 -29052 34740 -28988
rect 34613 -29068 34740 -29052
rect 34613 -29132 34660 -29068
rect 34724 -29132 34740 -29068
rect 34613 -29148 34740 -29132
rect 34613 -29212 34660 -29148
rect 34724 -29212 34740 -29148
rect 34613 -29228 34740 -29212
rect 34613 -29292 34660 -29228
rect 34724 -29292 34740 -29228
rect 34613 -29308 34740 -29292
rect 34613 -29372 34660 -29308
rect 34724 -29372 34740 -29308
rect 34613 -29388 34740 -29372
rect 34613 -29452 34660 -29388
rect 34724 -29452 34740 -29388
rect 34613 -29468 34740 -29452
rect 34613 -29532 34660 -29468
rect 34724 -29532 34740 -29468
rect 34613 -29548 34740 -29532
rect 34613 -29612 34660 -29548
rect 34724 -29612 34740 -29548
rect 34613 -29628 34740 -29612
rect 34613 -29692 34660 -29628
rect 34724 -29692 34740 -29628
rect 34613 -29708 34740 -29692
rect 34613 -29772 34660 -29708
rect 34724 -29772 34740 -29708
rect 34613 -29788 34740 -29772
rect 34613 -29852 34660 -29788
rect 34724 -29852 34740 -29788
rect 34613 -29868 34740 -29852
rect 34613 -29932 34660 -29868
rect 34724 -29932 34740 -29868
rect 34613 -29948 34740 -29932
rect 34613 -30012 34660 -29948
rect 34724 -30012 34740 -29948
rect 34613 -30028 34740 -30012
rect 34613 -30092 34660 -30028
rect 34724 -30092 34740 -30028
rect 34613 -30108 34740 -30092
rect 34613 -30172 34660 -30108
rect 34724 -30172 34740 -30108
rect 34613 -30188 34740 -30172
rect 34613 -30252 34660 -30188
rect 34724 -30252 34740 -30188
rect 34613 -30268 34740 -30252
rect 34613 -30332 34660 -30268
rect 34724 -30332 34740 -30268
rect 34613 -30348 34740 -30332
rect 34613 -30412 34660 -30348
rect 34724 -30412 34740 -30348
rect 34613 -30428 34740 -30412
rect 34613 -30492 34660 -30428
rect 34724 -30492 34740 -30428
rect 34613 -30508 34740 -30492
rect 34613 -30572 34660 -30508
rect 34724 -30572 34740 -30508
rect 34613 -30588 34740 -30572
rect 34613 -30652 34660 -30588
rect 34724 -30652 34740 -30588
rect 34613 -30668 34740 -30652
rect 34613 -30732 34660 -30668
rect 34724 -30732 34740 -30668
rect 34613 -30748 34740 -30732
rect 34613 -30812 34660 -30748
rect 34724 -30812 34740 -30748
rect 34613 -30828 34740 -30812
rect 34613 -30892 34660 -30828
rect 34724 -30892 34740 -30828
rect 34613 -30908 34740 -30892
rect 34613 -30972 34660 -30908
rect 34724 -30972 34740 -30908
rect 34613 -30988 34740 -30972
rect 34613 -31052 34660 -30988
rect 34724 -31052 34740 -30988
rect 34613 -31068 34740 -31052
rect 34613 -31132 34660 -31068
rect 34724 -31132 34740 -31068
rect 34613 -31148 34740 -31132
rect 34613 -31212 34660 -31148
rect 34724 -31212 34740 -31148
rect 34613 -31228 34740 -31212
rect 34613 -31292 34660 -31228
rect 34724 -31292 34740 -31228
rect 34613 -31308 34740 -31292
rect 34613 -31372 34660 -31308
rect 34724 -31372 34740 -31308
rect 34613 -31388 34740 -31372
rect 34613 -31452 34660 -31388
rect 34724 -31452 34740 -31388
rect 34613 -31468 34740 -31452
rect 34613 -31532 34660 -31468
rect 34724 -31532 34740 -31468
rect 34613 -31548 34740 -31532
rect 34613 -31612 34660 -31548
rect 34724 -31612 34740 -31548
rect 34613 -31628 34740 -31612
rect 34613 -31692 34660 -31628
rect 34724 -31692 34740 -31628
rect 34613 -31708 34740 -31692
rect 34613 -31772 34660 -31708
rect 34724 -31772 34740 -31708
rect 34613 -31788 34740 -31772
rect 34613 -31852 34660 -31788
rect 34724 -31852 34740 -31788
rect 34613 -31868 34740 -31852
rect 34613 -31932 34660 -31868
rect 34724 -31932 34740 -31868
rect 34613 -31948 34740 -31932
rect 34613 -32012 34660 -31948
rect 34724 -32012 34740 -31948
rect 34613 -32028 34740 -32012
rect 34613 -32092 34660 -32028
rect 34724 -32092 34740 -32028
rect 34613 -32108 34740 -32092
rect 34613 -32172 34660 -32108
rect 34724 -32172 34740 -32108
rect 34613 -32188 34740 -32172
rect 34613 -32252 34660 -32188
rect 34724 -32252 34740 -32188
rect 34613 -32268 34740 -32252
rect 34613 -32332 34660 -32268
rect 34724 -32332 34740 -32268
rect 34613 -32348 34740 -32332
rect 34613 -32412 34660 -32348
rect 34724 -32412 34740 -32348
rect 34613 -32428 34740 -32412
rect 34613 -32492 34660 -32428
rect 34724 -32492 34740 -32428
rect 34613 -32508 34740 -32492
rect 34613 -32572 34660 -32508
rect 34724 -32572 34740 -32508
rect 34613 -32588 34740 -32572
rect 34613 -32652 34660 -32588
rect 34724 -32652 34740 -32588
rect 34613 -32668 34740 -32652
rect 34613 -32732 34660 -32668
rect 34724 -32732 34740 -32668
rect 34613 -32748 34740 -32732
rect 34613 -32812 34660 -32748
rect 34724 -32812 34740 -32748
rect 34613 -32828 34740 -32812
rect 34613 -32892 34660 -32828
rect 34724 -32892 34740 -32828
rect 34613 -32908 34740 -32892
rect 34613 -32972 34660 -32908
rect 34724 -32972 34740 -32908
rect 34613 -32988 34740 -32972
rect 34613 -33052 34660 -32988
rect 34724 -33052 34740 -32988
rect 34613 -33068 34740 -33052
rect 34613 -33132 34660 -33068
rect 34724 -33132 34740 -33068
rect 34613 -33148 34740 -33132
rect 34613 -33212 34660 -33148
rect 34724 -33212 34740 -33148
rect 34613 -33228 34740 -33212
rect 34613 -33292 34660 -33228
rect 34724 -33292 34740 -33228
rect 34613 -33308 34740 -33292
rect 34613 -33372 34660 -33308
rect 34724 -33372 34740 -33308
rect 34613 -33388 34740 -33372
rect 34613 -33452 34660 -33388
rect 34724 -33452 34740 -33388
rect 34613 -33468 34740 -33452
rect 34613 -33532 34660 -33468
rect 34724 -33532 34740 -33468
rect 34613 -33548 34740 -33532
rect 34613 -33612 34660 -33548
rect 34724 -33612 34740 -33548
rect 34613 -33628 34740 -33612
rect 34613 -33692 34660 -33628
rect 34724 -33692 34740 -33628
rect 34613 -33708 34740 -33692
rect 34613 -33772 34660 -33708
rect 34724 -33772 34740 -33708
rect 34613 -33788 34740 -33772
rect 34613 -33852 34660 -33788
rect 34724 -33852 34740 -33788
rect 34613 -33868 34740 -33852
rect 34613 -33932 34660 -33868
rect 34724 -33932 34740 -33868
rect 34613 -33948 34740 -33932
rect 34613 -34012 34660 -33948
rect 34724 -34012 34740 -33948
rect 34613 -34028 34740 -34012
rect 34613 -34092 34660 -34028
rect 34724 -34092 34740 -34028
rect 34613 -34108 34740 -34092
rect 34613 -34172 34660 -34108
rect 34724 -34172 34740 -34108
rect 34613 -34188 34740 -34172
rect 34613 -34252 34660 -34188
rect 34724 -34252 34740 -34188
rect 34613 -34268 34740 -34252
rect 34613 -34332 34660 -34268
rect 34724 -34332 34740 -34268
rect 34613 -34348 34740 -34332
rect 34613 -34412 34660 -34348
rect 34724 -34412 34740 -34348
rect 34613 -34428 34740 -34412
rect 28294 -34508 28421 -34492
rect 28294 -34572 28341 -34508
rect 28405 -34572 28421 -34508
rect 28294 -34588 28421 -34572
rect 28294 -34712 28398 -34588
rect 28294 -34728 28421 -34712
rect 28294 -34792 28341 -34728
rect 28405 -34792 28421 -34728
rect 28294 -34808 28421 -34792
rect 21975 -34888 22102 -34872
rect 21975 -34952 22022 -34888
rect 22086 -34952 22102 -34888
rect 21975 -34968 22102 -34952
rect 21975 -35032 22022 -34968
rect 22086 -35032 22102 -34968
rect 21975 -35048 22102 -35032
rect 21975 -35112 22022 -35048
rect 22086 -35112 22102 -35048
rect 21975 -35128 22102 -35112
rect 21975 -35192 22022 -35128
rect 22086 -35192 22102 -35128
rect 21975 -35208 22102 -35192
rect 21975 -35272 22022 -35208
rect 22086 -35272 22102 -35208
rect 21975 -35288 22102 -35272
rect 21975 -35352 22022 -35288
rect 22086 -35352 22102 -35288
rect 21975 -35368 22102 -35352
rect 21975 -35432 22022 -35368
rect 22086 -35432 22102 -35368
rect 21975 -35448 22102 -35432
rect 21975 -35512 22022 -35448
rect 22086 -35512 22102 -35448
rect 21975 -35528 22102 -35512
rect 21975 -35592 22022 -35528
rect 22086 -35592 22102 -35528
rect 21975 -35608 22102 -35592
rect 21975 -35672 22022 -35608
rect 22086 -35672 22102 -35608
rect 21975 -35688 22102 -35672
rect 21975 -35752 22022 -35688
rect 22086 -35752 22102 -35688
rect 21975 -35768 22102 -35752
rect 21975 -35832 22022 -35768
rect 22086 -35832 22102 -35768
rect 21975 -35848 22102 -35832
rect 21975 -35912 22022 -35848
rect 22086 -35912 22102 -35848
rect 21975 -35928 22102 -35912
rect 21975 -35992 22022 -35928
rect 22086 -35992 22102 -35928
rect 21975 -36008 22102 -35992
rect 21975 -36072 22022 -36008
rect 22086 -36072 22102 -36008
rect 21975 -36088 22102 -36072
rect 21975 -36152 22022 -36088
rect 22086 -36152 22102 -36088
rect 21975 -36168 22102 -36152
rect 21975 -36232 22022 -36168
rect 22086 -36232 22102 -36168
rect 21975 -36248 22102 -36232
rect 21975 -36312 22022 -36248
rect 22086 -36312 22102 -36248
rect 21975 -36328 22102 -36312
rect 21975 -36392 22022 -36328
rect 22086 -36392 22102 -36328
rect 21975 -36408 22102 -36392
rect 21975 -36472 22022 -36408
rect 22086 -36472 22102 -36408
rect 21975 -36488 22102 -36472
rect 21975 -36552 22022 -36488
rect 22086 -36552 22102 -36488
rect 21975 -36568 22102 -36552
rect 21975 -36632 22022 -36568
rect 22086 -36632 22102 -36568
rect 21975 -36648 22102 -36632
rect 21975 -36712 22022 -36648
rect 22086 -36712 22102 -36648
rect 21975 -36728 22102 -36712
rect 21975 -36792 22022 -36728
rect 22086 -36792 22102 -36728
rect 21975 -36808 22102 -36792
rect 21975 -36872 22022 -36808
rect 22086 -36872 22102 -36808
rect 21975 -36888 22102 -36872
rect 21975 -36952 22022 -36888
rect 22086 -36952 22102 -36888
rect 21975 -36968 22102 -36952
rect 21975 -37032 22022 -36968
rect 22086 -37032 22102 -36968
rect 21975 -37048 22102 -37032
rect 21975 -37112 22022 -37048
rect 22086 -37112 22102 -37048
rect 21975 -37128 22102 -37112
rect 21975 -37192 22022 -37128
rect 22086 -37192 22102 -37128
rect 21975 -37208 22102 -37192
rect 21975 -37272 22022 -37208
rect 22086 -37272 22102 -37208
rect 21975 -37288 22102 -37272
rect 21975 -37352 22022 -37288
rect 22086 -37352 22102 -37288
rect 21975 -37368 22102 -37352
rect 21975 -37432 22022 -37368
rect 22086 -37432 22102 -37368
rect 21975 -37448 22102 -37432
rect 21975 -37512 22022 -37448
rect 22086 -37512 22102 -37448
rect 21975 -37528 22102 -37512
rect 21975 -37592 22022 -37528
rect 22086 -37592 22102 -37528
rect 21975 -37608 22102 -37592
rect 21975 -37672 22022 -37608
rect 22086 -37672 22102 -37608
rect 21975 -37688 22102 -37672
rect 21975 -37752 22022 -37688
rect 22086 -37752 22102 -37688
rect 21975 -37768 22102 -37752
rect 21975 -37832 22022 -37768
rect 22086 -37832 22102 -37768
rect 21975 -37848 22102 -37832
rect 21975 -37912 22022 -37848
rect 22086 -37912 22102 -37848
rect 21975 -37928 22102 -37912
rect 21975 -37992 22022 -37928
rect 22086 -37992 22102 -37928
rect 21975 -38008 22102 -37992
rect 21975 -38072 22022 -38008
rect 22086 -38072 22102 -38008
rect 21975 -38088 22102 -38072
rect 21975 -38152 22022 -38088
rect 22086 -38152 22102 -38088
rect 21975 -38168 22102 -38152
rect 21975 -38232 22022 -38168
rect 22086 -38232 22102 -38168
rect 21975 -38248 22102 -38232
rect 21975 -38312 22022 -38248
rect 22086 -38312 22102 -38248
rect 21975 -38328 22102 -38312
rect 21975 -38392 22022 -38328
rect 22086 -38392 22102 -38328
rect 21975 -38408 22102 -38392
rect 21975 -38472 22022 -38408
rect 22086 -38472 22102 -38408
rect 21975 -38488 22102 -38472
rect 21975 -38552 22022 -38488
rect 22086 -38552 22102 -38488
rect 21975 -38568 22102 -38552
rect 21975 -38632 22022 -38568
rect 22086 -38632 22102 -38568
rect 21975 -38648 22102 -38632
rect 21975 -38712 22022 -38648
rect 22086 -38712 22102 -38648
rect 21975 -38728 22102 -38712
rect 21975 -38792 22022 -38728
rect 22086 -38792 22102 -38728
rect 21975 -38808 22102 -38792
rect 21975 -38872 22022 -38808
rect 22086 -38872 22102 -38808
rect 21975 -38888 22102 -38872
rect 21975 -38952 22022 -38888
rect 22086 -38952 22102 -38888
rect 21975 -38968 22102 -38952
rect 21975 -39032 22022 -38968
rect 22086 -39032 22102 -38968
rect 21975 -39048 22102 -39032
rect 21975 -39112 22022 -39048
rect 22086 -39112 22102 -39048
rect 21975 -39128 22102 -39112
rect 21975 -39192 22022 -39128
rect 22086 -39192 22102 -39128
rect 21975 -39208 22102 -39192
rect 21975 -39272 22022 -39208
rect 22086 -39272 22102 -39208
rect 21975 -39288 22102 -39272
rect 21975 -39352 22022 -39288
rect 22086 -39352 22102 -39288
rect 21975 -39368 22102 -39352
rect 21975 -39432 22022 -39368
rect 22086 -39432 22102 -39368
rect 21975 -39448 22102 -39432
rect 21975 -39512 22022 -39448
rect 22086 -39512 22102 -39448
rect 21975 -39528 22102 -39512
rect 21975 -39592 22022 -39528
rect 22086 -39592 22102 -39528
rect 21975 -39608 22102 -39592
rect 21975 -39672 22022 -39608
rect 22086 -39672 22102 -39608
rect 21975 -39688 22102 -39672
rect 21975 -39752 22022 -39688
rect 22086 -39752 22102 -39688
rect 21975 -39768 22102 -39752
rect 21975 -39832 22022 -39768
rect 22086 -39832 22102 -39768
rect 21975 -39848 22102 -39832
rect 21975 -39912 22022 -39848
rect 22086 -39912 22102 -39848
rect 21975 -39928 22102 -39912
rect 21975 -39992 22022 -39928
rect 22086 -39992 22102 -39928
rect 21975 -40008 22102 -39992
rect 21975 -40072 22022 -40008
rect 22086 -40072 22102 -40008
rect 21975 -40088 22102 -40072
rect 21975 -40152 22022 -40088
rect 22086 -40152 22102 -40088
rect 21975 -40168 22102 -40152
rect 21975 -40232 22022 -40168
rect 22086 -40232 22102 -40168
rect 21975 -40248 22102 -40232
rect 21975 -40312 22022 -40248
rect 22086 -40312 22102 -40248
rect 21975 -40328 22102 -40312
rect 21975 -40392 22022 -40328
rect 22086 -40392 22102 -40328
rect 21975 -40408 22102 -40392
rect 21975 -40472 22022 -40408
rect 22086 -40472 22102 -40408
rect 21975 -40488 22102 -40472
rect 21975 -40552 22022 -40488
rect 22086 -40552 22102 -40488
rect 21975 -40568 22102 -40552
rect 21975 -40632 22022 -40568
rect 22086 -40632 22102 -40568
rect 21975 -40648 22102 -40632
rect 21975 -40712 22022 -40648
rect 22086 -40712 22102 -40648
rect 21975 -40728 22102 -40712
rect 15656 -40808 15783 -40792
rect 15656 -40872 15703 -40808
rect 15767 -40872 15783 -40808
rect 15656 -40888 15783 -40872
rect 15656 -41012 15760 -40888
rect 15656 -41028 15783 -41012
rect 15656 -41092 15703 -41028
rect 15767 -41092 15783 -41028
rect 15656 -41108 15783 -41092
rect 9337 -41188 9464 -41172
rect 9337 -41252 9384 -41188
rect 9448 -41252 9464 -41188
rect 9337 -41268 9464 -41252
rect 9337 -41332 9384 -41268
rect 9448 -41332 9464 -41268
rect 9337 -41348 9464 -41332
rect 9337 -41412 9384 -41348
rect 9448 -41412 9464 -41348
rect 9337 -41428 9464 -41412
rect 9337 -41492 9384 -41428
rect 9448 -41492 9464 -41428
rect 9337 -41508 9464 -41492
rect 9337 -41572 9384 -41508
rect 9448 -41572 9464 -41508
rect 9337 -41588 9464 -41572
rect 9337 -41652 9384 -41588
rect 9448 -41652 9464 -41588
rect 9337 -41668 9464 -41652
rect 9337 -41732 9384 -41668
rect 9448 -41732 9464 -41668
rect 9337 -41748 9464 -41732
rect 9337 -41812 9384 -41748
rect 9448 -41812 9464 -41748
rect 9337 -41828 9464 -41812
rect 9337 -41892 9384 -41828
rect 9448 -41892 9464 -41828
rect 9337 -41908 9464 -41892
rect 9337 -41972 9384 -41908
rect 9448 -41972 9464 -41908
rect 9337 -41988 9464 -41972
rect 9337 -42052 9384 -41988
rect 9448 -42052 9464 -41988
rect 9337 -42068 9464 -42052
rect 9337 -42132 9384 -42068
rect 9448 -42132 9464 -42068
rect 9337 -42148 9464 -42132
rect 9337 -42212 9384 -42148
rect 9448 -42212 9464 -42148
rect 9337 -42228 9464 -42212
rect 9337 -42292 9384 -42228
rect 9448 -42292 9464 -42228
rect 9337 -42308 9464 -42292
rect 9337 -42372 9384 -42308
rect 9448 -42372 9464 -42308
rect 9337 -42388 9464 -42372
rect 9337 -42452 9384 -42388
rect 9448 -42452 9464 -42388
rect 9337 -42468 9464 -42452
rect 9337 -42532 9384 -42468
rect 9448 -42532 9464 -42468
rect 9337 -42548 9464 -42532
rect 9337 -42612 9384 -42548
rect 9448 -42612 9464 -42548
rect 9337 -42628 9464 -42612
rect 9337 -42692 9384 -42628
rect 9448 -42692 9464 -42628
rect 9337 -42708 9464 -42692
rect 9337 -42772 9384 -42708
rect 9448 -42772 9464 -42708
rect 9337 -42788 9464 -42772
rect 9337 -42852 9384 -42788
rect 9448 -42852 9464 -42788
rect 9337 -42868 9464 -42852
rect 9337 -42932 9384 -42868
rect 9448 -42932 9464 -42868
rect 9337 -42948 9464 -42932
rect 9337 -43012 9384 -42948
rect 9448 -43012 9464 -42948
rect 9337 -43028 9464 -43012
rect 9337 -43092 9384 -43028
rect 9448 -43092 9464 -43028
rect 9337 -43108 9464 -43092
rect 9337 -43172 9384 -43108
rect 9448 -43172 9464 -43108
rect 9337 -43188 9464 -43172
rect 9337 -43252 9384 -43188
rect 9448 -43252 9464 -43188
rect 9337 -43268 9464 -43252
rect 9337 -43332 9384 -43268
rect 9448 -43332 9464 -43268
rect 9337 -43348 9464 -43332
rect 9337 -43412 9384 -43348
rect 9448 -43412 9464 -43348
rect 9337 -43428 9464 -43412
rect 9337 -43492 9384 -43428
rect 9448 -43492 9464 -43428
rect 9337 -43508 9464 -43492
rect 9337 -43572 9384 -43508
rect 9448 -43572 9464 -43508
rect 9337 -43588 9464 -43572
rect 9337 -43652 9384 -43588
rect 9448 -43652 9464 -43588
rect 9337 -43668 9464 -43652
rect 9337 -43732 9384 -43668
rect 9448 -43732 9464 -43668
rect 9337 -43748 9464 -43732
rect 9337 -43812 9384 -43748
rect 9448 -43812 9464 -43748
rect 9337 -43828 9464 -43812
rect 9337 -43892 9384 -43828
rect 9448 -43892 9464 -43828
rect 9337 -43908 9464 -43892
rect 9337 -43972 9384 -43908
rect 9448 -43972 9464 -43908
rect 9337 -43988 9464 -43972
rect 9337 -44052 9384 -43988
rect 9448 -44052 9464 -43988
rect 9337 -44068 9464 -44052
rect 9337 -44132 9384 -44068
rect 9448 -44132 9464 -44068
rect 9337 -44148 9464 -44132
rect 9337 -44212 9384 -44148
rect 9448 -44212 9464 -44148
rect 9337 -44228 9464 -44212
rect 9337 -44292 9384 -44228
rect 9448 -44292 9464 -44228
rect 9337 -44308 9464 -44292
rect 9337 -44372 9384 -44308
rect 9448 -44372 9464 -44308
rect 9337 -44388 9464 -44372
rect 9337 -44452 9384 -44388
rect 9448 -44452 9464 -44388
rect 9337 -44468 9464 -44452
rect 9337 -44532 9384 -44468
rect 9448 -44532 9464 -44468
rect 9337 -44548 9464 -44532
rect 9337 -44612 9384 -44548
rect 9448 -44612 9464 -44548
rect 9337 -44628 9464 -44612
rect 9337 -44692 9384 -44628
rect 9448 -44692 9464 -44628
rect 9337 -44708 9464 -44692
rect 9337 -44772 9384 -44708
rect 9448 -44772 9464 -44708
rect 9337 -44788 9464 -44772
rect 9337 -44852 9384 -44788
rect 9448 -44852 9464 -44788
rect 9337 -44868 9464 -44852
rect 9337 -44932 9384 -44868
rect 9448 -44932 9464 -44868
rect 9337 -44948 9464 -44932
rect 9337 -45012 9384 -44948
rect 9448 -45012 9464 -44948
rect 9337 -45028 9464 -45012
rect 9337 -45092 9384 -45028
rect 9448 -45092 9464 -45028
rect 9337 -45108 9464 -45092
rect 9337 -45172 9384 -45108
rect 9448 -45172 9464 -45108
rect 9337 -45188 9464 -45172
rect 9337 -45252 9384 -45188
rect 9448 -45252 9464 -45188
rect 9337 -45268 9464 -45252
rect 9337 -45332 9384 -45268
rect 9448 -45332 9464 -45268
rect 9337 -45348 9464 -45332
rect 9337 -45412 9384 -45348
rect 9448 -45412 9464 -45348
rect 9337 -45428 9464 -45412
rect 9337 -45492 9384 -45428
rect 9448 -45492 9464 -45428
rect 9337 -45508 9464 -45492
rect 9337 -45572 9384 -45508
rect 9448 -45572 9464 -45508
rect 9337 -45588 9464 -45572
rect 9337 -45652 9384 -45588
rect 9448 -45652 9464 -45588
rect 9337 -45668 9464 -45652
rect 9337 -45732 9384 -45668
rect 9448 -45732 9464 -45668
rect 9337 -45748 9464 -45732
rect 9337 -45812 9384 -45748
rect 9448 -45812 9464 -45748
rect 9337 -45828 9464 -45812
rect 9337 -45892 9384 -45828
rect 9448 -45892 9464 -45828
rect 9337 -45908 9464 -45892
rect 9337 -45972 9384 -45908
rect 9448 -45972 9464 -45908
rect 9337 -45988 9464 -45972
rect 9337 -46052 9384 -45988
rect 9448 -46052 9464 -45988
rect 9337 -46068 9464 -46052
rect 9337 -46132 9384 -46068
rect 9448 -46132 9464 -46068
rect 9337 -46148 9464 -46132
rect 9337 -46212 9384 -46148
rect 9448 -46212 9464 -46148
rect 9337 -46228 9464 -46212
rect 9337 -46292 9384 -46228
rect 9448 -46292 9464 -46228
rect 9337 -46308 9464 -46292
rect 9337 -46372 9384 -46308
rect 9448 -46372 9464 -46308
rect 9337 -46388 9464 -46372
rect 9337 -46452 9384 -46388
rect 9448 -46452 9464 -46388
rect 9337 -46468 9464 -46452
rect 9337 -46532 9384 -46468
rect 9448 -46532 9464 -46468
rect 9337 -46548 9464 -46532
rect 9337 -46612 9384 -46548
rect 9448 -46612 9464 -46548
rect 9337 -46628 9464 -46612
rect 9337 -46692 9384 -46628
rect 9448 -46692 9464 -46628
rect 9337 -46708 9464 -46692
rect 9337 -46772 9384 -46708
rect 9448 -46772 9464 -46708
rect 9337 -46788 9464 -46772
rect 9337 -46852 9384 -46788
rect 9448 -46852 9464 -46788
rect 9337 -46868 9464 -46852
rect 9337 -46932 9384 -46868
rect 9448 -46932 9464 -46868
rect 9337 -46948 9464 -46932
rect 9337 -47012 9384 -46948
rect 9448 -47012 9464 -46948
rect 9337 -47028 9464 -47012
rect 3018 -47108 3145 -47092
rect 3018 -47172 3065 -47108
rect 3129 -47172 3145 -47108
rect 3018 -47188 3145 -47172
rect 3018 -47250 3122 -47188
rect 6217 -47250 6321 -47061
rect 9337 -47092 9384 -47028
rect 9448 -47092 9464 -47028
rect 9627 -41148 15549 -41139
rect 9627 -47052 9636 -41148
rect 15540 -47052 15549 -41148
rect 9627 -47061 15549 -47052
rect 15656 -41172 15703 -41108
rect 15767 -41172 15783 -41108
rect 18855 -41139 18959 -40761
rect 21975 -40792 22022 -40728
rect 22086 -40792 22102 -40728
rect 22265 -34848 28187 -34839
rect 22265 -40752 22274 -34848
rect 28178 -40752 28187 -34848
rect 22265 -40761 28187 -40752
rect 28294 -34872 28341 -34808
rect 28405 -34872 28421 -34808
rect 31493 -34839 31597 -34461
rect 34613 -34492 34660 -34428
rect 34724 -34492 34740 -34428
rect 34903 -28548 40825 -28539
rect 34903 -34452 34912 -28548
rect 40816 -34452 40825 -28548
rect 34903 -34461 40825 -34452
rect 40932 -28572 40979 -28508
rect 41043 -28572 41059 -28508
rect 44131 -28539 44235 -28161
rect 47251 -28192 47298 -28128
rect 47362 -28192 47378 -28128
rect 47251 -28208 47378 -28192
rect 47251 -28272 47298 -28208
rect 47362 -28272 47378 -28208
rect 47251 -28288 47378 -28272
rect 47251 -28412 47355 -28288
rect 47251 -28428 47378 -28412
rect 47251 -28492 47298 -28428
rect 47362 -28492 47378 -28428
rect 47251 -28508 47378 -28492
rect 40932 -28588 41059 -28572
rect 40932 -28652 40979 -28588
rect 41043 -28652 41059 -28588
rect 40932 -28668 41059 -28652
rect 40932 -28732 40979 -28668
rect 41043 -28732 41059 -28668
rect 40932 -28748 41059 -28732
rect 40932 -28812 40979 -28748
rect 41043 -28812 41059 -28748
rect 40932 -28828 41059 -28812
rect 40932 -28892 40979 -28828
rect 41043 -28892 41059 -28828
rect 40932 -28908 41059 -28892
rect 40932 -28972 40979 -28908
rect 41043 -28972 41059 -28908
rect 40932 -28988 41059 -28972
rect 40932 -29052 40979 -28988
rect 41043 -29052 41059 -28988
rect 40932 -29068 41059 -29052
rect 40932 -29132 40979 -29068
rect 41043 -29132 41059 -29068
rect 40932 -29148 41059 -29132
rect 40932 -29212 40979 -29148
rect 41043 -29212 41059 -29148
rect 40932 -29228 41059 -29212
rect 40932 -29292 40979 -29228
rect 41043 -29292 41059 -29228
rect 40932 -29308 41059 -29292
rect 40932 -29372 40979 -29308
rect 41043 -29372 41059 -29308
rect 40932 -29388 41059 -29372
rect 40932 -29452 40979 -29388
rect 41043 -29452 41059 -29388
rect 40932 -29468 41059 -29452
rect 40932 -29532 40979 -29468
rect 41043 -29532 41059 -29468
rect 40932 -29548 41059 -29532
rect 40932 -29612 40979 -29548
rect 41043 -29612 41059 -29548
rect 40932 -29628 41059 -29612
rect 40932 -29692 40979 -29628
rect 41043 -29692 41059 -29628
rect 40932 -29708 41059 -29692
rect 40932 -29772 40979 -29708
rect 41043 -29772 41059 -29708
rect 40932 -29788 41059 -29772
rect 40932 -29852 40979 -29788
rect 41043 -29852 41059 -29788
rect 40932 -29868 41059 -29852
rect 40932 -29932 40979 -29868
rect 41043 -29932 41059 -29868
rect 40932 -29948 41059 -29932
rect 40932 -30012 40979 -29948
rect 41043 -30012 41059 -29948
rect 40932 -30028 41059 -30012
rect 40932 -30092 40979 -30028
rect 41043 -30092 41059 -30028
rect 40932 -30108 41059 -30092
rect 40932 -30172 40979 -30108
rect 41043 -30172 41059 -30108
rect 40932 -30188 41059 -30172
rect 40932 -30252 40979 -30188
rect 41043 -30252 41059 -30188
rect 40932 -30268 41059 -30252
rect 40932 -30332 40979 -30268
rect 41043 -30332 41059 -30268
rect 40932 -30348 41059 -30332
rect 40932 -30412 40979 -30348
rect 41043 -30412 41059 -30348
rect 40932 -30428 41059 -30412
rect 40932 -30492 40979 -30428
rect 41043 -30492 41059 -30428
rect 40932 -30508 41059 -30492
rect 40932 -30572 40979 -30508
rect 41043 -30572 41059 -30508
rect 40932 -30588 41059 -30572
rect 40932 -30652 40979 -30588
rect 41043 -30652 41059 -30588
rect 40932 -30668 41059 -30652
rect 40932 -30732 40979 -30668
rect 41043 -30732 41059 -30668
rect 40932 -30748 41059 -30732
rect 40932 -30812 40979 -30748
rect 41043 -30812 41059 -30748
rect 40932 -30828 41059 -30812
rect 40932 -30892 40979 -30828
rect 41043 -30892 41059 -30828
rect 40932 -30908 41059 -30892
rect 40932 -30972 40979 -30908
rect 41043 -30972 41059 -30908
rect 40932 -30988 41059 -30972
rect 40932 -31052 40979 -30988
rect 41043 -31052 41059 -30988
rect 40932 -31068 41059 -31052
rect 40932 -31132 40979 -31068
rect 41043 -31132 41059 -31068
rect 40932 -31148 41059 -31132
rect 40932 -31212 40979 -31148
rect 41043 -31212 41059 -31148
rect 40932 -31228 41059 -31212
rect 40932 -31292 40979 -31228
rect 41043 -31292 41059 -31228
rect 40932 -31308 41059 -31292
rect 40932 -31372 40979 -31308
rect 41043 -31372 41059 -31308
rect 40932 -31388 41059 -31372
rect 40932 -31452 40979 -31388
rect 41043 -31452 41059 -31388
rect 40932 -31468 41059 -31452
rect 40932 -31532 40979 -31468
rect 41043 -31532 41059 -31468
rect 40932 -31548 41059 -31532
rect 40932 -31612 40979 -31548
rect 41043 -31612 41059 -31548
rect 40932 -31628 41059 -31612
rect 40932 -31692 40979 -31628
rect 41043 -31692 41059 -31628
rect 40932 -31708 41059 -31692
rect 40932 -31772 40979 -31708
rect 41043 -31772 41059 -31708
rect 40932 -31788 41059 -31772
rect 40932 -31852 40979 -31788
rect 41043 -31852 41059 -31788
rect 40932 -31868 41059 -31852
rect 40932 -31932 40979 -31868
rect 41043 -31932 41059 -31868
rect 40932 -31948 41059 -31932
rect 40932 -32012 40979 -31948
rect 41043 -32012 41059 -31948
rect 40932 -32028 41059 -32012
rect 40932 -32092 40979 -32028
rect 41043 -32092 41059 -32028
rect 40932 -32108 41059 -32092
rect 40932 -32172 40979 -32108
rect 41043 -32172 41059 -32108
rect 40932 -32188 41059 -32172
rect 40932 -32252 40979 -32188
rect 41043 -32252 41059 -32188
rect 40932 -32268 41059 -32252
rect 40932 -32332 40979 -32268
rect 41043 -32332 41059 -32268
rect 40932 -32348 41059 -32332
rect 40932 -32412 40979 -32348
rect 41043 -32412 41059 -32348
rect 40932 -32428 41059 -32412
rect 40932 -32492 40979 -32428
rect 41043 -32492 41059 -32428
rect 40932 -32508 41059 -32492
rect 40932 -32572 40979 -32508
rect 41043 -32572 41059 -32508
rect 40932 -32588 41059 -32572
rect 40932 -32652 40979 -32588
rect 41043 -32652 41059 -32588
rect 40932 -32668 41059 -32652
rect 40932 -32732 40979 -32668
rect 41043 -32732 41059 -32668
rect 40932 -32748 41059 -32732
rect 40932 -32812 40979 -32748
rect 41043 -32812 41059 -32748
rect 40932 -32828 41059 -32812
rect 40932 -32892 40979 -32828
rect 41043 -32892 41059 -32828
rect 40932 -32908 41059 -32892
rect 40932 -32972 40979 -32908
rect 41043 -32972 41059 -32908
rect 40932 -32988 41059 -32972
rect 40932 -33052 40979 -32988
rect 41043 -33052 41059 -32988
rect 40932 -33068 41059 -33052
rect 40932 -33132 40979 -33068
rect 41043 -33132 41059 -33068
rect 40932 -33148 41059 -33132
rect 40932 -33212 40979 -33148
rect 41043 -33212 41059 -33148
rect 40932 -33228 41059 -33212
rect 40932 -33292 40979 -33228
rect 41043 -33292 41059 -33228
rect 40932 -33308 41059 -33292
rect 40932 -33372 40979 -33308
rect 41043 -33372 41059 -33308
rect 40932 -33388 41059 -33372
rect 40932 -33452 40979 -33388
rect 41043 -33452 41059 -33388
rect 40932 -33468 41059 -33452
rect 40932 -33532 40979 -33468
rect 41043 -33532 41059 -33468
rect 40932 -33548 41059 -33532
rect 40932 -33612 40979 -33548
rect 41043 -33612 41059 -33548
rect 40932 -33628 41059 -33612
rect 40932 -33692 40979 -33628
rect 41043 -33692 41059 -33628
rect 40932 -33708 41059 -33692
rect 40932 -33772 40979 -33708
rect 41043 -33772 41059 -33708
rect 40932 -33788 41059 -33772
rect 40932 -33852 40979 -33788
rect 41043 -33852 41059 -33788
rect 40932 -33868 41059 -33852
rect 40932 -33932 40979 -33868
rect 41043 -33932 41059 -33868
rect 40932 -33948 41059 -33932
rect 40932 -34012 40979 -33948
rect 41043 -34012 41059 -33948
rect 40932 -34028 41059 -34012
rect 40932 -34092 40979 -34028
rect 41043 -34092 41059 -34028
rect 40932 -34108 41059 -34092
rect 40932 -34172 40979 -34108
rect 41043 -34172 41059 -34108
rect 40932 -34188 41059 -34172
rect 40932 -34252 40979 -34188
rect 41043 -34252 41059 -34188
rect 40932 -34268 41059 -34252
rect 40932 -34332 40979 -34268
rect 41043 -34332 41059 -34268
rect 40932 -34348 41059 -34332
rect 40932 -34412 40979 -34348
rect 41043 -34412 41059 -34348
rect 40932 -34428 41059 -34412
rect 34613 -34508 34740 -34492
rect 34613 -34572 34660 -34508
rect 34724 -34572 34740 -34508
rect 34613 -34588 34740 -34572
rect 34613 -34712 34717 -34588
rect 34613 -34728 34740 -34712
rect 34613 -34792 34660 -34728
rect 34724 -34792 34740 -34728
rect 34613 -34808 34740 -34792
rect 28294 -34888 28421 -34872
rect 28294 -34952 28341 -34888
rect 28405 -34952 28421 -34888
rect 28294 -34968 28421 -34952
rect 28294 -35032 28341 -34968
rect 28405 -35032 28421 -34968
rect 28294 -35048 28421 -35032
rect 28294 -35112 28341 -35048
rect 28405 -35112 28421 -35048
rect 28294 -35128 28421 -35112
rect 28294 -35192 28341 -35128
rect 28405 -35192 28421 -35128
rect 28294 -35208 28421 -35192
rect 28294 -35272 28341 -35208
rect 28405 -35272 28421 -35208
rect 28294 -35288 28421 -35272
rect 28294 -35352 28341 -35288
rect 28405 -35352 28421 -35288
rect 28294 -35368 28421 -35352
rect 28294 -35432 28341 -35368
rect 28405 -35432 28421 -35368
rect 28294 -35448 28421 -35432
rect 28294 -35512 28341 -35448
rect 28405 -35512 28421 -35448
rect 28294 -35528 28421 -35512
rect 28294 -35592 28341 -35528
rect 28405 -35592 28421 -35528
rect 28294 -35608 28421 -35592
rect 28294 -35672 28341 -35608
rect 28405 -35672 28421 -35608
rect 28294 -35688 28421 -35672
rect 28294 -35752 28341 -35688
rect 28405 -35752 28421 -35688
rect 28294 -35768 28421 -35752
rect 28294 -35832 28341 -35768
rect 28405 -35832 28421 -35768
rect 28294 -35848 28421 -35832
rect 28294 -35912 28341 -35848
rect 28405 -35912 28421 -35848
rect 28294 -35928 28421 -35912
rect 28294 -35992 28341 -35928
rect 28405 -35992 28421 -35928
rect 28294 -36008 28421 -35992
rect 28294 -36072 28341 -36008
rect 28405 -36072 28421 -36008
rect 28294 -36088 28421 -36072
rect 28294 -36152 28341 -36088
rect 28405 -36152 28421 -36088
rect 28294 -36168 28421 -36152
rect 28294 -36232 28341 -36168
rect 28405 -36232 28421 -36168
rect 28294 -36248 28421 -36232
rect 28294 -36312 28341 -36248
rect 28405 -36312 28421 -36248
rect 28294 -36328 28421 -36312
rect 28294 -36392 28341 -36328
rect 28405 -36392 28421 -36328
rect 28294 -36408 28421 -36392
rect 28294 -36472 28341 -36408
rect 28405 -36472 28421 -36408
rect 28294 -36488 28421 -36472
rect 28294 -36552 28341 -36488
rect 28405 -36552 28421 -36488
rect 28294 -36568 28421 -36552
rect 28294 -36632 28341 -36568
rect 28405 -36632 28421 -36568
rect 28294 -36648 28421 -36632
rect 28294 -36712 28341 -36648
rect 28405 -36712 28421 -36648
rect 28294 -36728 28421 -36712
rect 28294 -36792 28341 -36728
rect 28405 -36792 28421 -36728
rect 28294 -36808 28421 -36792
rect 28294 -36872 28341 -36808
rect 28405 -36872 28421 -36808
rect 28294 -36888 28421 -36872
rect 28294 -36952 28341 -36888
rect 28405 -36952 28421 -36888
rect 28294 -36968 28421 -36952
rect 28294 -37032 28341 -36968
rect 28405 -37032 28421 -36968
rect 28294 -37048 28421 -37032
rect 28294 -37112 28341 -37048
rect 28405 -37112 28421 -37048
rect 28294 -37128 28421 -37112
rect 28294 -37192 28341 -37128
rect 28405 -37192 28421 -37128
rect 28294 -37208 28421 -37192
rect 28294 -37272 28341 -37208
rect 28405 -37272 28421 -37208
rect 28294 -37288 28421 -37272
rect 28294 -37352 28341 -37288
rect 28405 -37352 28421 -37288
rect 28294 -37368 28421 -37352
rect 28294 -37432 28341 -37368
rect 28405 -37432 28421 -37368
rect 28294 -37448 28421 -37432
rect 28294 -37512 28341 -37448
rect 28405 -37512 28421 -37448
rect 28294 -37528 28421 -37512
rect 28294 -37592 28341 -37528
rect 28405 -37592 28421 -37528
rect 28294 -37608 28421 -37592
rect 28294 -37672 28341 -37608
rect 28405 -37672 28421 -37608
rect 28294 -37688 28421 -37672
rect 28294 -37752 28341 -37688
rect 28405 -37752 28421 -37688
rect 28294 -37768 28421 -37752
rect 28294 -37832 28341 -37768
rect 28405 -37832 28421 -37768
rect 28294 -37848 28421 -37832
rect 28294 -37912 28341 -37848
rect 28405 -37912 28421 -37848
rect 28294 -37928 28421 -37912
rect 28294 -37992 28341 -37928
rect 28405 -37992 28421 -37928
rect 28294 -38008 28421 -37992
rect 28294 -38072 28341 -38008
rect 28405 -38072 28421 -38008
rect 28294 -38088 28421 -38072
rect 28294 -38152 28341 -38088
rect 28405 -38152 28421 -38088
rect 28294 -38168 28421 -38152
rect 28294 -38232 28341 -38168
rect 28405 -38232 28421 -38168
rect 28294 -38248 28421 -38232
rect 28294 -38312 28341 -38248
rect 28405 -38312 28421 -38248
rect 28294 -38328 28421 -38312
rect 28294 -38392 28341 -38328
rect 28405 -38392 28421 -38328
rect 28294 -38408 28421 -38392
rect 28294 -38472 28341 -38408
rect 28405 -38472 28421 -38408
rect 28294 -38488 28421 -38472
rect 28294 -38552 28341 -38488
rect 28405 -38552 28421 -38488
rect 28294 -38568 28421 -38552
rect 28294 -38632 28341 -38568
rect 28405 -38632 28421 -38568
rect 28294 -38648 28421 -38632
rect 28294 -38712 28341 -38648
rect 28405 -38712 28421 -38648
rect 28294 -38728 28421 -38712
rect 28294 -38792 28341 -38728
rect 28405 -38792 28421 -38728
rect 28294 -38808 28421 -38792
rect 28294 -38872 28341 -38808
rect 28405 -38872 28421 -38808
rect 28294 -38888 28421 -38872
rect 28294 -38952 28341 -38888
rect 28405 -38952 28421 -38888
rect 28294 -38968 28421 -38952
rect 28294 -39032 28341 -38968
rect 28405 -39032 28421 -38968
rect 28294 -39048 28421 -39032
rect 28294 -39112 28341 -39048
rect 28405 -39112 28421 -39048
rect 28294 -39128 28421 -39112
rect 28294 -39192 28341 -39128
rect 28405 -39192 28421 -39128
rect 28294 -39208 28421 -39192
rect 28294 -39272 28341 -39208
rect 28405 -39272 28421 -39208
rect 28294 -39288 28421 -39272
rect 28294 -39352 28341 -39288
rect 28405 -39352 28421 -39288
rect 28294 -39368 28421 -39352
rect 28294 -39432 28341 -39368
rect 28405 -39432 28421 -39368
rect 28294 -39448 28421 -39432
rect 28294 -39512 28341 -39448
rect 28405 -39512 28421 -39448
rect 28294 -39528 28421 -39512
rect 28294 -39592 28341 -39528
rect 28405 -39592 28421 -39528
rect 28294 -39608 28421 -39592
rect 28294 -39672 28341 -39608
rect 28405 -39672 28421 -39608
rect 28294 -39688 28421 -39672
rect 28294 -39752 28341 -39688
rect 28405 -39752 28421 -39688
rect 28294 -39768 28421 -39752
rect 28294 -39832 28341 -39768
rect 28405 -39832 28421 -39768
rect 28294 -39848 28421 -39832
rect 28294 -39912 28341 -39848
rect 28405 -39912 28421 -39848
rect 28294 -39928 28421 -39912
rect 28294 -39992 28341 -39928
rect 28405 -39992 28421 -39928
rect 28294 -40008 28421 -39992
rect 28294 -40072 28341 -40008
rect 28405 -40072 28421 -40008
rect 28294 -40088 28421 -40072
rect 28294 -40152 28341 -40088
rect 28405 -40152 28421 -40088
rect 28294 -40168 28421 -40152
rect 28294 -40232 28341 -40168
rect 28405 -40232 28421 -40168
rect 28294 -40248 28421 -40232
rect 28294 -40312 28341 -40248
rect 28405 -40312 28421 -40248
rect 28294 -40328 28421 -40312
rect 28294 -40392 28341 -40328
rect 28405 -40392 28421 -40328
rect 28294 -40408 28421 -40392
rect 28294 -40472 28341 -40408
rect 28405 -40472 28421 -40408
rect 28294 -40488 28421 -40472
rect 28294 -40552 28341 -40488
rect 28405 -40552 28421 -40488
rect 28294 -40568 28421 -40552
rect 28294 -40632 28341 -40568
rect 28405 -40632 28421 -40568
rect 28294 -40648 28421 -40632
rect 28294 -40712 28341 -40648
rect 28405 -40712 28421 -40648
rect 28294 -40728 28421 -40712
rect 21975 -40808 22102 -40792
rect 21975 -40872 22022 -40808
rect 22086 -40872 22102 -40808
rect 21975 -40888 22102 -40872
rect 21975 -41012 22079 -40888
rect 21975 -41028 22102 -41012
rect 21975 -41092 22022 -41028
rect 22086 -41092 22102 -41028
rect 21975 -41108 22102 -41092
rect 15656 -41188 15783 -41172
rect 15656 -41252 15703 -41188
rect 15767 -41252 15783 -41188
rect 15656 -41268 15783 -41252
rect 15656 -41332 15703 -41268
rect 15767 -41332 15783 -41268
rect 15656 -41348 15783 -41332
rect 15656 -41412 15703 -41348
rect 15767 -41412 15783 -41348
rect 15656 -41428 15783 -41412
rect 15656 -41492 15703 -41428
rect 15767 -41492 15783 -41428
rect 15656 -41508 15783 -41492
rect 15656 -41572 15703 -41508
rect 15767 -41572 15783 -41508
rect 15656 -41588 15783 -41572
rect 15656 -41652 15703 -41588
rect 15767 -41652 15783 -41588
rect 15656 -41668 15783 -41652
rect 15656 -41732 15703 -41668
rect 15767 -41732 15783 -41668
rect 15656 -41748 15783 -41732
rect 15656 -41812 15703 -41748
rect 15767 -41812 15783 -41748
rect 15656 -41828 15783 -41812
rect 15656 -41892 15703 -41828
rect 15767 -41892 15783 -41828
rect 15656 -41908 15783 -41892
rect 15656 -41972 15703 -41908
rect 15767 -41972 15783 -41908
rect 15656 -41988 15783 -41972
rect 15656 -42052 15703 -41988
rect 15767 -42052 15783 -41988
rect 15656 -42068 15783 -42052
rect 15656 -42132 15703 -42068
rect 15767 -42132 15783 -42068
rect 15656 -42148 15783 -42132
rect 15656 -42212 15703 -42148
rect 15767 -42212 15783 -42148
rect 15656 -42228 15783 -42212
rect 15656 -42292 15703 -42228
rect 15767 -42292 15783 -42228
rect 15656 -42308 15783 -42292
rect 15656 -42372 15703 -42308
rect 15767 -42372 15783 -42308
rect 15656 -42388 15783 -42372
rect 15656 -42452 15703 -42388
rect 15767 -42452 15783 -42388
rect 15656 -42468 15783 -42452
rect 15656 -42532 15703 -42468
rect 15767 -42532 15783 -42468
rect 15656 -42548 15783 -42532
rect 15656 -42612 15703 -42548
rect 15767 -42612 15783 -42548
rect 15656 -42628 15783 -42612
rect 15656 -42692 15703 -42628
rect 15767 -42692 15783 -42628
rect 15656 -42708 15783 -42692
rect 15656 -42772 15703 -42708
rect 15767 -42772 15783 -42708
rect 15656 -42788 15783 -42772
rect 15656 -42852 15703 -42788
rect 15767 -42852 15783 -42788
rect 15656 -42868 15783 -42852
rect 15656 -42932 15703 -42868
rect 15767 -42932 15783 -42868
rect 15656 -42948 15783 -42932
rect 15656 -43012 15703 -42948
rect 15767 -43012 15783 -42948
rect 15656 -43028 15783 -43012
rect 15656 -43092 15703 -43028
rect 15767 -43092 15783 -43028
rect 15656 -43108 15783 -43092
rect 15656 -43172 15703 -43108
rect 15767 -43172 15783 -43108
rect 15656 -43188 15783 -43172
rect 15656 -43252 15703 -43188
rect 15767 -43252 15783 -43188
rect 15656 -43268 15783 -43252
rect 15656 -43332 15703 -43268
rect 15767 -43332 15783 -43268
rect 15656 -43348 15783 -43332
rect 15656 -43412 15703 -43348
rect 15767 -43412 15783 -43348
rect 15656 -43428 15783 -43412
rect 15656 -43492 15703 -43428
rect 15767 -43492 15783 -43428
rect 15656 -43508 15783 -43492
rect 15656 -43572 15703 -43508
rect 15767 -43572 15783 -43508
rect 15656 -43588 15783 -43572
rect 15656 -43652 15703 -43588
rect 15767 -43652 15783 -43588
rect 15656 -43668 15783 -43652
rect 15656 -43732 15703 -43668
rect 15767 -43732 15783 -43668
rect 15656 -43748 15783 -43732
rect 15656 -43812 15703 -43748
rect 15767 -43812 15783 -43748
rect 15656 -43828 15783 -43812
rect 15656 -43892 15703 -43828
rect 15767 -43892 15783 -43828
rect 15656 -43908 15783 -43892
rect 15656 -43972 15703 -43908
rect 15767 -43972 15783 -43908
rect 15656 -43988 15783 -43972
rect 15656 -44052 15703 -43988
rect 15767 -44052 15783 -43988
rect 15656 -44068 15783 -44052
rect 15656 -44132 15703 -44068
rect 15767 -44132 15783 -44068
rect 15656 -44148 15783 -44132
rect 15656 -44212 15703 -44148
rect 15767 -44212 15783 -44148
rect 15656 -44228 15783 -44212
rect 15656 -44292 15703 -44228
rect 15767 -44292 15783 -44228
rect 15656 -44308 15783 -44292
rect 15656 -44372 15703 -44308
rect 15767 -44372 15783 -44308
rect 15656 -44388 15783 -44372
rect 15656 -44452 15703 -44388
rect 15767 -44452 15783 -44388
rect 15656 -44468 15783 -44452
rect 15656 -44532 15703 -44468
rect 15767 -44532 15783 -44468
rect 15656 -44548 15783 -44532
rect 15656 -44612 15703 -44548
rect 15767 -44612 15783 -44548
rect 15656 -44628 15783 -44612
rect 15656 -44692 15703 -44628
rect 15767 -44692 15783 -44628
rect 15656 -44708 15783 -44692
rect 15656 -44772 15703 -44708
rect 15767 -44772 15783 -44708
rect 15656 -44788 15783 -44772
rect 15656 -44852 15703 -44788
rect 15767 -44852 15783 -44788
rect 15656 -44868 15783 -44852
rect 15656 -44932 15703 -44868
rect 15767 -44932 15783 -44868
rect 15656 -44948 15783 -44932
rect 15656 -45012 15703 -44948
rect 15767 -45012 15783 -44948
rect 15656 -45028 15783 -45012
rect 15656 -45092 15703 -45028
rect 15767 -45092 15783 -45028
rect 15656 -45108 15783 -45092
rect 15656 -45172 15703 -45108
rect 15767 -45172 15783 -45108
rect 15656 -45188 15783 -45172
rect 15656 -45252 15703 -45188
rect 15767 -45252 15783 -45188
rect 15656 -45268 15783 -45252
rect 15656 -45332 15703 -45268
rect 15767 -45332 15783 -45268
rect 15656 -45348 15783 -45332
rect 15656 -45412 15703 -45348
rect 15767 -45412 15783 -45348
rect 15656 -45428 15783 -45412
rect 15656 -45492 15703 -45428
rect 15767 -45492 15783 -45428
rect 15656 -45508 15783 -45492
rect 15656 -45572 15703 -45508
rect 15767 -45572 15783 -45508
rect 15656 -45588 15783 -45572
rect 15656 -45652 15703 -45588
rect 15767 -45652 15783 -45588
rect 15656 -45668 15783 -45652
rect 15656 -45732 15703 -45668
rect 15767 -45732 15783 -45668
rect 15656 -45748 15783 -45732
rect 15656 -45812 15703 -45748
rect 15767 -45812 15783 -45748
rect 15656 -45828 15783 -45812
rect 15656 -45892 15703 -45828
rect 15767 -45892 15783 -45828
rect 15656 -45908 15783 -45892
rect 15656 -45972 15703 -45908
rect 15767 -45972 15783 -45908
rect 15656 -45988 15783 -45972
rect 15656 -46052 15703 -45988
rect 15767 -46052 15783 -45988
rect 15656 -46068 15783 -46052
rect 15656 -46132 15703 -46068
rect 15767 -46132 15783 -46068
rect 15656 -46148 15783 -46132
rect 15656 -46212 15703 -46148
rect 15767 -46212 15783 -46148
rect 15656 -46228 15783 -46212
rect 15656 -46292 15703 -46228
rect 15767 -46292 15783 -46228
rect 15656 -46308 15783 -46292
rect 15656 -46372 15703 -46308
rect 15767 -46372 15783 -46308
rect 15656 -46388 15783 -46372
rect 15656 -46452 15703 -46388
rect 15767 -46452 15783 -46388
rect 15656 -46468 15783 -46452
rect 15656 -46532 15703 -46468
rect 15767 -46532 15783 -46468
rect 15656 -46548 15783 -46532
rect 15656 -46612 15703 -46548
rect 15767 -46612 15783 -46548
rect 15656 -46628 15783 -46612
rect 15656 -46692 15703 -46628
rect 15767 -46692 15783 -46628
rect 15656 -46708 15783 -46692
rect 15656 -46772 15703 -46708
rect 15767 -46772 15783 -46708
rect 15656 -46788 15783 -46772
rect 15656 -46852 15703 -46788
rect 15767 -46852 15783 -46788
rect 15656 -46868 15783 -46852
rect 15656 -46932 15703 -46868
rect 15767 -46932 15783 -46868
rect 15656 -46948 15783 -46932
rect 15656 -47012 15703 -46948
rect 15767 -47012 15783 -46948
rect 15656 -47028 15783 -47012
rect 9337 -47108 9464 -47092
rect 9337 -47172 9384 -47108
rect 9448 -47172 9464 -47108
rect 9337 -47188 9464 -47172
rect 9337 -47250 9441 -47188
rect 12536 -47250 12640 -47061
rect 15656 -47092 15703 -47028
rect 15767 -47092 15783 -47028
rect 15946 -41148 21868 -41139
rect 15946 -47052 15955 -41148
rect 21859 -47052 21868 -41148
rect 15946 -47061 21868 -47052
rect 21975 -41172 22022 -41108
rect 22086 -41172 22102 -41108
rect 25174 -41139 25278 -40761
rect 28294 -40792 28341 -40728
rect 28405 -40792 28421 -40728
rect 28584 -34848 34506 -34839
rect 28584 -40752 28593 -34848
rect 34497 -40752 34506 -34848
rect 28584 -40761 34506 -40752
rect 34613 -34872 34660 -34808
rect 34724 -34872 34740 -34808
rect 37812 -34839 37916 -34461
rect 40932 -34492 40979 -34428
rect 41043 -34492 41059 -34428
rect 41222 -28548 47144 -28539
rect 41222 -34452 41231 -28548
rect 47135 -34452 47144 -28548
rect 41222 -34461 47144 -34452
rect 47251 -28572 47298 -28508
rect 47362 -28572 47378 -28508
rect 47251 -28588 47378 -28572
rect 47251 -28652 47298 -28588
rect 47362 -28652 47378 -28588
rect 47251 -28668 47378 -28652
rect 47251 -28732 47298 -28668
rect 47362 -28732 47378 -28668
rect 47251 -28748 47378 -28732
rect 47251 -28812 47298 -28748
rect 47362 -28812 47378 -28748
rect 47251 -28828 47378 -28812
rect 47251 -28892 47298 -28828
rect 47362 -28892 47378 -28828
rect 47251 -28908 47378 -28892
rect 47251 -28972 47298 -28908
rect 47362 -28972 47378 -28908
rect 47251 -28988 47378 -28972
rect 47251 -29052 47298 -28988
rect 47362 -29052 47378 -28988
rect 47251 -29068 47378 -29052
rect 47251 -29132 47298 -29068
rect 47362 -29132 47378 -29068
rect 47251 -29148 47378 -29132
rect 47251 -29212 47298 -29148
rect 47362 -29212 47378 -29148
rect 47251 -29228 47378 -29212
rect 47251 -29292 47298 -29228
rect 47362 -29292 47378 -29228
rect 47251 -29308 47378 -29292
rect 47251 -29372 47298 -29308
rect 47362 -29372 47378 -29308
rect 47251 -29388 47378 -29372
rect 47251 -29452 47298 -29388
rect 47362 -29452 47378 -29388
rect 47251 -29468 47378 -29452
rect 47251 -29532 47298 -29468
rect 47362 -29532 47378 -29468
rect 47251 -29548 47378 -29532
rect 47251 -29612 47298 -29548
rect 47362 -29612 47378 -29548
rect 47251 -29628 47378 -29612
rect 47251 -29692 47298 -29628
rect 47362 -29692 47378 -29628
rect 47251 -29708 47378 -29692
rect 47251 -29772 47298 -29708
rect 47362 -29772 47378 -29708
rect 47251 -29788 47378 -29772
rect 47251 -29852 47298 -29788
rect 47362 -29852 47378 -29788
rect 47251 -29868 47378 -29852
rect 47251 -29932 47298 -29868
rect 47362 -29932 47378 -29868
rect 47251 -29948 47378 -29932
rect 47251 -30012 47298 -29948
rect 47362 -30012 47378 -29948
rect 47251 -30028 47378 -30012
rect 47251 -30092 47298 -30028
rect 47362 -30092 47378 -30028
rect 47251 -30108 47378 -30092
rect 47251 -30172 47298 -30108
rect 47362 -30172 47378 -30108
rect 47251 -30188 47378 -30172
rect 47251 -30252 47298 -30188
rect 47362 -30252 47378 -30188
rect 47251 -30268 47378 -30252
rect 47251 -30332 47298 -30268
rect 47362 -30332 47378 -30268
rect 47251 -30348 47378 -30332
rect 47251 -30412 47298 -30348
rect 47362 -30412 47378 -30348
rect 47251 -30428 47378 -30412
rect 47251 -30492 47298 -30428
rect 47362 -30492 47378 -30428
rect 47251 -30508 47378 -30492
rect 47251 -30572 47298 -30508
rect 47362 -30572 47378 -30508
rect 47251 -30588 47378 -30572
rect 47251 -30652 47298 -30588
rect 47362 -30652 47378 -30588
rect 47251 -30668 47378 -30652
rect 47251 -30732 47298 -30668
rect 47362 -30732 47378 -30668
rect 47251 -30748 47378 -30732
rect 47251 -30812 47298 -30748
rect 47362 -30812 47378 -30748
rect 47251 -30828 47378 -30812
rect 47251 -30892 47298 -30828
rect 47362 -30892 47378 -30828
rect 47251 -30908 47378 -30892
rect 47251 -30972 47298 -30908
rect 47362 -30972 47378 -30908
rect 47251 -30988 47378 -30972
rect 47251 -31052 47298 -30988
rect 47362 -31052 47378 -30988
rect 47251 -31068 47378 -31052
rect 47251 -31132 47298 -31068
rect 47362 -31132 47378 -31068
rect 47251 -31148 47378 -31132
rect 47251 -31212 47298 -31148
rect 47362 -31212 47378 -31148
rect 47251 -31228 47378 -31212
rect 47251 -31292 47298 -31228
rect 47362 -31292 47378 -31228
rect 47251 -31308 47378 -31292
rect 47251 -31372 47298 -31308
rect 47362 -31372 47378 -31308
rect 47251 -31388 47378 -31372
rect 47251 -31452 47298 -31388
rect 47362 -31452 47378 -31388
rect 47251 -31468 47378 -31452
rect 47251 -31532 47298 -31468
rect 47362 -31532 47378 -31468
rect 47251 -31548 47378 -31532
rect 47251 -31612 47298 -31548
rect 47362 -31612 47378 -31548
rect 47251 -31628 47378 -31612
rect 47251 -31692 47298 -31628
rect 47362 -31692 47378 -31628
rect 47251 -31708 47378 -31692
rect 47251 -31772 47298 -31708
rect 47362 -31772 47378 -31708
rect 47251 -31788 47378 -31772
rect 47251 -31852 47298 -31788
rect 47362 -31852 47378 -31788
rect 47251 -31868 47378 -31852
rect 47251 -31932 47298 -31868
rect 47362 -31932 47378 -31868
rect 47251 -31948 47378 -31932
rect 47251 -32012 47298 -31948
rect 47362 -32012 47378 -31948
rect 47251 -32028 47378 -32012
rect 47251 -32092 47298 -32028
rect 47362 -32092 47378 -32028
rect 47251 -32108 47378 -32092
rect 47251 -32172 47298 -32108
rect 47362 -32172 47378 -32108
rect 47251 -32188 47378 -32172
rect 47251 -32252 47298 -32188
rect 47362 -32252 47378 -32188
rect 47251 -32268 47378 -32252
rect 47251 -32332 47298 -32268
rect 47362 -32332 47378 -32268
rect 47251 -32348 47378 -32332
rect 47251 -32412 47298 -32348
rect 47362 -32412 47378 -32348
rect 47251 -32428 47378 -32412
rect 47251 -32492 47298 -32428
rect 47362 -32492 47378 -32428
rect 47251 -32508 47378 -32492
rect 47251 -32572 47298 -32508
rect 47362 -32572 47378 -32508
rect 47251 -32588 47378 -32572
rect 47251 -32652 47298 -32588
rect 47362 -32652 47378 -32588
rect 47251 -32668 47378 -32652
rect 47251 -32732 47298 -32668
rect 47362 -32732 47378 -32668
rect 47251 -32748 47378 -32732
rect 47251 -32812 47298 -32748
rect 47362 -32812 47378 -32748
rect 47251 -32828 47378 -32812
rect 47251 -32892 47298 -32828
rect 47362 -32892 47378 -32828
rect 47251 -32908 47378 -32892
rect 47251 -32972 47298 -32908
rect 47362 -32972 47378 -32908
rect 47251 -32988 47378 -32972
rect 47251 -33052 47298 -32988
rect 47362 -33052 47378 -32988
rect 47251 -33068 47378 -33052
rect 47251 -33132 47298 -33068
rect 47362 -33132 47378 -33068
rect 47251 -33148 47378 -33132
rect 47251 -33212 47298 -33148
rect 47362 -33212 47378 -33148
rect 47251 -33228 47378 -33212
rect 47251 -33292 47298 -33228
rect 47362 -33292 47378 -33228
rect 47251 -33308 47378 -33292
rect 47251 -33372 47298 -33308
rect 47362 -33372 47378 -33308
rect 47251 -33388 47378 -33372
rect 47251 -33452 47298 -33388
rect 47362 -33452 47378 -33388
rect 47251 -33468 47378 -33452
rect 47251 -33532 47298 -33468
rect 47362 -33532 47378 -33468
rect 47251 -33548 47378 -33532
rect 47251 -33612 47298 -33548
rect 47362 -33612 47378 -33548
rect 47251 -33628 47378 -33612
rect 47251 -33692 47298 -33628
rect 47362 -33692 47378 -33628
rect 47251 -33708 47378 -33692
rect 47251 -33772 47298 -33708
rect 47362 -33772 47378 -33708
rect 47251 -33788 47378 -33772
rect 47251 -33852 47298 -33788
rect 47362 -33852 47378 -33788
rect 47251 -33868 47378 -33852
rect 47251 -33932 47298 -33868
rect 47362 -33932 47378 -33868
rect 47251 -33948 47378 -33932
rect 47251 -34012 47298 -33948
rect 47362 -34012 47378 -33948
rect 47251 -34028 47378 -34012
rect 47251 -34092 47298 -34028
rect 47362 -34092 47378 -34028
rect 47251 -34108 47378 -34092
rect 47251 -34172 47298 -34108
rect 47362 -34172 47378 -34108
rect 47251 -34188 47378 -34172
rect 47251 -34252 47298 -34188
rect 47362 -34252 47378 -34188
rect 47251 -34268 47378 -34252
rect 47251 -34332 47298 -34268
rect 47362 -34332 47378 -34268
rect 47251 -34348 47378 -34332
rect 47251 -34412 47298 -34348
rect 47362 -34412 47378 -34348
rect 47251 -34428 47378 -34412
rect 40932 -34508 41059 -34492
rect 40932 -34572 40979 -34508
rect 41043 -34572 41059 -34508
rect 40932 -34588 41059 -34572
rect 40932 -34712 41036 -34588
rect 40932 -34728 41059 -34712
rect 40932 -34792 40979 -34728
rect 41043 -34792 41059 -34728
rect 40932 -34808 41059 -34792
rect 34613 -34888 34740 -34872
rect 34613 -34952 34660 -34888
rect 34724 -34952 34740 -34888
rect 34613 -34968 34740 -34952
rect 34613 -35032 34660 -34968
rect 34724 -35032 34740 -34968
rect 34613 -35048 34740 -35032
rect 34613 -35112 34660 -35048
rect 34724 -35112 34740 -35048
rect 34613 -35128 34740 -35112
rect 34613 -35192 34660 -35128
rect 34724 -35192 34740 -35128
rect 34613 -35208 34740 -35192
rect 34613 -35272 34660 -35208
rect 34724 -35272 34740 -35208
rect 34613 -35288 34740 -35272
rect 34613 -35352 34660 -35288
rect 34724 -35352 34740 -35288
rect 34613 -35368 34740 -35352
rect 34613 -35432 34660 -35368
rect 34724 -35432 34740 -35368
rect 34613 -35448 34740 -35432
rect 34613 -35512 34660 -35448
rect 34724 -35512 34740 -35448
rect 34613 -35528 34740 -35512
rect 34613 -35592 34660 -35528
rect 34724 -35592 34740 -35528
rect 34613 -35608 34740 -35592
rect 34613 -35672 34660 -35608
rect 34724 -35672 34740 -35608
rect 34613 -35688 34740 -35672
rect 34613 -35752 34660 -35688
rect 34724 -35752 34740 -35688
rect 34613 -35768 34740 -35752
rect 34613 -35832 34660 -35768
rect 34724 -35832 34740 -35768
rect 34613 -35848 34740 -35832
rect 34613 -35912 34660 -35848
rect 34724 -35912 34740 -35848
rect 34613 -35928 34740 -35912
rect 34613 -35992 34660 -35928
rect 34724 -35992 34740 -35928
rect 34613 -36008 34740 -35992
rect 34613 -36072 34660 -36008
rect 34724 -36072 34740 -36008
rect 34613 -36088 34740 -36072
rect 34613 -36152 34660 -36088
rect 34724 -36152 34740 -36088
rect 34613 -36168 34740 -36152
rect 34613 -36232 34660 -36168
rect 34724 -36232 34740 -36168
rect 34613 -36248 34740 -36232
rect 34613 -36312 34660 -36248
rect 34724 -36312 34740 -36248
rect 34613 -36328 34740 -36312
rect 34613 -36392 34660 -36328
rect 34724 -36392 34740 -36328
rect 34613 -36408 34740 -36392
rect 34613 -36472 34660 -36408
rect 34724 -36472 34740 -36408
rect 34613 -36488 34740 -36472
rect 34613 -36552 34660 -36488
rect 34724 -36552 34740 -36488
rect 34613 -36568 34740 -36552
rect 34613 -36632 34660 -36568
rect 34724 -36632 34740 -36568
rect 34613 -36648 34740 -36632
rect 34613 -36712 34660 -36648
rect 34724 -36712 34740 -36648
rect 34613 -36728 34740 -36712
rect 34613 -36792 34660 -36728
rect 34724 -36792 34740 -36728
rect 34613 -36808 34740 -36792
rect 34613 -36872 34660 -36808
rect 34724 -36872 34740 -36808
rect 34613 -36888 34740 -36872
rect 34613 -36952 34660 -36888
rect 34724 -36952 34740 -36888
rect 34613 -36968 34740 -36952
rect 34613 -37032 34660 -36968
rect 34724 -37032 34740 -36968
rect 34613 -37048 34740 -37032
rect 34613 -37112 34660 -37048
rect 34724 -37112 34740 -37048
rect 34613 -37128 34740 -37112
rect 34613 -37192 34660 -37128
rect 34724 -37192 34740 -37128
rect 34613 -37208 34740 -37192
rect 34613 -37272 34660 -37208
rect 34724 -37272 34740 -37208
rect 34613 -37288 34740 -37272
rect 34613 -37352 34660 -37288
rect 34724 -37352 34740 -37288
rect 34613 -37368 34740 -37352
rect 34613 -37432 34660 -37368
rect 34724 -37432 34740 -37368
rect 34613 -37448 34740 -37432
rect 34613 -37512 34660 -37448
rect 34724 -37512 34740 -37448
rect 34613 -37528 34740 -37512
rect 34613 -37592 34660 -37528
rect 34724 -37592 34740 -37528
rect 34613 -37608 34740 -37592
rect 34613 -37672 34660 -37608
rect 34724 -37672 34740 -37608
rect 34613 -37688 34740 -37672
rect 34613 -37752 34660 -37688
rect 34724 -37752 34740 -37688
rect 34613 -37768 34740 -37752
rect 34613 -37832 34660 -37768
rect 34724 -37832 34740 -37768
rect 34613 -37848 34740 -37832
rect 34613 -37912 34660 -37848
rect 34724 -37912 34740 -37848
rect 34613 -37928 34740 -37912
rect 34613 -37992 34660 -37928
rect 34724 -37992 34740 -37928
rect 34613 -38008 34740 -37992
rect 34613 -38072 34660 -38008
rect 34724 -38072 34740 -38008
rect 34613 -38088 34740 -38072
rect 34613 -38152 34660 -38088
rect 34724 -38152 34740 -38088
rect 34613 -38168 34740 -38152
rect 34613 -38232 34660 -38168
rect 34724 -38232 34740 -38168
rect 34613 -38248 34740 -38232
rect 34613 -38312 34660 -38248
rect 34724 -38312 34740 -38248
rect 34613 -38328 34740 -38312
rect 34613 -38392 34660 -38328
rect 34724 -38392 34740 -38328
rect 34613 -38408 34740 -38392
rect 34613 -38472 34660 -38408
rect 34724 -38472 34740 -38408
rect 34613 -38488 34740 -38472
rect 34613 -38552 34660 -38488
rect 34724 -38552 34740 -38488
rect 34613 -38568 34740 -38552
rect 34613 -38632 34660 -38568
rect 34724 -38632 34740 -38568
rect 34613 -38648 34740 -38632
rect 34613 -38712 34660 -38648
rect 34724 -38712 34740 -38648
rect 34613 -38728 34740 -38712
rect 34613 -38792 34660 -38728
rect 34724 -38792 34740 -38728
rect 34613 -38808 34740 -38792
rect 34613 -38872 34660 -38808
rect 34724 -38872 34740 -38808
rect 34613 -38888 34740 -38872
rect 34613 -38952 34660 -38888
rect 34724 -38952 34740 -38888
rect 34613 -38968 34740 -38952
rect 34613 -39032 34660 -38968
rect 34724 -39032 34740 -38968
rect 34613 -39048 34740 -39032
rect 34613 -39112 34660 -39048
rect 34724 -39112 34740 -39048
rect 34613 -39128 34740 -39112
rect 34613 -39192 34660 -39128
rect 34724 -39192 34740 -39128
rect 34613 -39208 34740 -39192
rect 34613 -39272 34660 -39208
rect 34724 -39272 34740 -39208
rect 34613 -39288 34740 -39272
rect 34613 -39352 34660 -39288
rect 34724 -39352 34740 -39288
rect 34613 -39368 34740 -39352
rect 34613 -39432 34660 -39368
rect 34724 -39432 34740 -39368
rect 34613 -39448 34740 -39432
rect 34613 -39512 34660 -39448
rect 34724 -39512 34740 -39448
rect 34613 -39528 34740 -39512
rect 34613 -39592 34660 -39528
rect 34724 -39592 34740 -39528
rect 34613 -39608 34740 -39592
rect 34613 -39672 34660 -39608
rect 34724 -39672 34740 -39608
rect 34613 -39688 34740 -39672
rect 34613 -39752 34660 -39688
rect 34724 -39752 34740 -39688
rect 34613 -39768 34740 -39752
rect 34613 -39832 34660 -39768
rect 34724 -39832 34740 -39768
rect 34613 -39848 34740 -39832
rect 34613 -39912 34660 -39848
rect 34724 -39912 34740 -39848
rect 34613 -39928 34740 -39912
rect 34613 -39992 34660 -39928
rect 34724 -39992 34740 -39928
rect 34613 -40008 34740 -39992
rect 34613 -40072 34660 -40008
rect 34724 -40072 34740 -40008
rect 34613 -40088 34740 -40072
rect 34613 -40152 34660 -40088
rect 34724 -40152 34740 -40088
rect 34613 -40168 34740 -40152
rect 34613 -40232 34660 -40168
rect 34724 -40232 34740 -40168
rect 34613 -40248 34740 -40232
rect 34613 -40312 34660 -40248
rect 34724 -40312 34740 -40248
rect 34613 -40328 34740 -40312
rect 34613 -40392 34660 -40328
rect 34724 -40392 34740 -40328
rect 34613 -40408 34740 -40392
rect 34613 -40472 34660 -40408
rect 34724 -40472 34740 -40408
rect 34613 -40488 34740 -40472
rect 34613 -40552 34660 -40488
rect 34724 -40552 34740 -40488
rect 34613 -40568 34740 -40552
rect 34613 -40632 34660 -40568
rect 34724 -40632 34740 -40568
rect 34613 -40648 34740 -40632
rect 34613 -40712 34660 -40648
rect 34724 -40712 34740 -40648
rect 34613 -40728 34740 -40712
rect 28294 -40808 28421 -40792
rect 28294 -40872 28341 -40808
rect 28405 -40872 28421 -40808
rect 28294 -40888 28421 -40872
rect 28294 -41012 28398 -40888
rect 28294 -41028 28421 -41012
rect 28294 -41092 28341 -41028
rect 28405 -41092 28421 -41028
rect 28294 -41108 28421 -41092
rect 21975 -41188 22102 -41172
rect 21975 -41252 22022 -41188
rect 22086 -41252 22102 -41188
rect 21975 -41268 22102 -41252
rect 21975 -41332 22022 -41268
rect 22086 -41332 22102 -41268
rect 21975 -41348 22102 -41332
rect 21975 -41412 22022 -41348
rect 22086 -41412 22102 -41348
rect 21975 -41428 22102 -41412
rect 21975 -41492 22022 -41428
rect 22086 -41492 22102 -41428
rect 21975 -41508 22102 -41492
rect 21975 -41572 22022 -41508
rect 22086 -41572 22102 -41508
rect 21975 -41588 22102 -41572
rect 21975 -41652 22022 -41588
rect 22086 -41652 22102 -41588
rect 21975 -41668 22102 -41652
rect 21975 -41732 22022 -41668
rect 22086 -41732 22102 -41668
rect 21975 -41748 22102 -41732
rect 21975 -41812 22022 -41748
rect 22086 -41812 22102 -41748
rect 21975 -41828 22102 -41812
rect 21975 -41892 22022 -41828
rect 22086 -41892 22102 -41828
rect 21975 -41908 22102 -41892
rect 21975 -41972 22022 -41908
rect 22086 -41972 22102 -41908
rect 21975 -41988 22102 -41972
rect 21975 -42052 22022 -41988
rect 22086 -42052 22102 -41988
rect 21975 -42068 22102 -42052
rect 21975 -42132 22022 -42068
rect 22086 -42132 22102 -42068
rect 21975 -42148 22102 -42132
rect 21975 -42212 22022 -42148
rect 22086 -42212 22102 -42148
rect 21975 -42228 22102 -42212
rect 21975 -42292 22022 -42228
rect 22086 -42292 22102 -42228
rect 21975 -42308 22102 -42292
rect 21975 -42372 22022 -42308
rect 22086 -42372 22102 -42308
rect 21975 -42388 22102 -42372
rect 21975 -42452 22022 -42388
rect 22086 -42452 22102 -42388
rect 21975 -42468 22102 -42452
rect 21975 -42532 22022 -42468
rect 22086 -42532 22102 -42468
rect 21975 -42548 22102 -42532
rect 21975 -42612 22022 -42548
rect 22086 -42612 22102 -42548
rect 21975 -42628 22102 -42612
rect 21975 -42692 22022 -42628
rect 22086 -42692 22102 -42628
rect 21975 -42708 22102 -42692
rect 21975 -42772 22022 -42708
rect 22086 -42772 22102 -42708
rect 21975 -42788 22102 -42772
rect 21975 -42852 22022 -42788
rect 22086 -42852 22102 -42788
rect 21975 -42868 22102 -42852
rect 21975 -42932 22022 -42868
rect 22086 -42932 22102 -42868
rect 21975 -42948 22102 -42932
rect 21975 -43012 22022 -42948
rect 22086 -43012 22102 -42948
rect 21975 -43028 22102 -43012
rect 21975 -43092 22022 -43028
rect 22086 -43092 22102 -43028
rect 21975 -43108 22102 -43092
rect 21975 -43172 22022 -43108
rect 22086 -43172 22102 -43108
rect 21975 -43188 22102 -43172
rect 21975 -43252 22022 -43188
rect 22086 -43252 22102 -43188
rect 21975 -43268 22102 -43252
rect 21975 -43332 22022 -43268
rect 22086 -43332 22102 -43268
rect 21975 -43348 22102 -43332
rect 21975 -43412 22022 -43348
rect 22086 -43412 22102 -43348
rect 21975 -43428 22102 -43412
rect 21975 -43492 22022 -43428
rect 22086 -43492 22102 -43428
rect 21975 -43508 22102 -43492
rect 21975 -43572 22022 -43508
rect 22086 -43572 22102 -43508
rect 21975 -43588 22102 -43572
rect 21975 -43652 22022 -43588
rect 22086 -43652 22102 -43588
rect 21975 -43668 22102 -43652
rect 21975 -43732 22022 -43668
rect 22086 -43732 22102 -43668
rect 21975 -43748 22102 -43732
rect 21975 -43812 22022 -43748
rect 22086 -43812 22102 -43748
rect 21975 -43828 22102 -43812
rect 21975 -43892 22022 -43828
rect 22086 -43892 22102 -43828
rect 21975 -43908 22102 -43892
rect 21975 -43972 22022 -43908
rect 22086 -43972 22102 -43908
rect 21975 -43988 22102 -43972
rect 21975 -44052 22022 -43988
rect 22086 -44052 22102 -43988
rect 21975 -44068 22102 -44052
rect 21975 -44132 22022 -44068
rect 22086 -44132 22102 -44068
rect 21975 -44148 22102 -44132
rect 21975 -44212 22022 -44148
rect 22086 -44212 22102 -44148
rect 21975 -44228 22102 -44212
rect 21975 -44292 22022 -44228
rect 22086 -44292 22102 -44228
rect 21975 -44308 22102 -44292
rect 21975 -44372 22022 -44308
rect 22086 -44372 22102 -44308
rect 21975 -44388 22102 -44372
rect 21975 -44452 22022 -44388
rect 22086 -44452 22102 -44388
rect 21975 -44468 22102 -44452
rect 21975 -44532 22022 -44468
rect 22086 -44532 22102 -44468
rect 21975 -44548 22102 -44532
rect 21975 -44612 22022 -44548
rect 22086 -44612 22102 -44548
rect 21975 -44628 22102 -44612
rect 21975 -44692 22022 -44628
rect 22086 -44692 22102 -44628
rect 21975 -44708 22102 -44692
rect 21975 -44772 22022 -44708
rect 22086 -44772 22102 -44708
rect 21975 -44788 22102 -44772
rect 21975 -44852 22022 -44788
rect 22086 -44852 22102 -44788
rect 21975 -44868 22102 -44852
rect 21975 -44932 22022 -44868
rect 22086 -44932 22102 -44868
rect 21975 -44948 22102 -44932
rect 21975 -45012 22022 -44948
rect 22086 -45012 22102 -44948
rect 21975 -45028 22102 -45012
rect 21975 -45092 22022 -45028
rect 22086 -45092 22102 -45028
rect 21975 -45108 22102 -45092
rect 21975 -45172 22022 -45108
rect 22086 -45172 22102 -45108
rect 21975 -45188 22102 -45172
rect 21975 -45252 22022 -45188
rect 22086 -45252 22102 -45188
rect 21975 -45268 22102 -45252
rect 21975 -45332 22022 -45268
rect 22086 -45332 22102 -45268
rect 21975 -45348 22102 -45332
rect 21975 -45412 22022 -45348
rect 22086 -45412 22102 -45348
rect 21975 -45428 22102 -45412
rect 21975 -45492 22022 -45428
rect 22086 -45492 22102 -45428
rect 21975 -45508 22102 -45492
rect 21975 -45572 22022 -45508
rect 22086 -45572 22102 -45508
rect 21975 -45588 22102 -45572
rect 21975 -45652 22022 -45588
rect 22086 -45652 22102 -45588
rect 21975 -45668 22102 -45652
rect 21975 -45732 22022 -45668
rect 22086 -45732 22102 -45668
rect 21975 -45748 22102 -45732
rect 21975 -45812 22022 -45748
rect 22086 -45812 22102 -45748
rect 21975 -45828 22102 -45812
rect 21975 -45892 22022 -45828
rect 22086 -45892 22102 -45828
rect 21975 -45908 22102 -45892
rect 21975 -45972 22022 -45908
rect 22086 -45972 22102 -45908
rect 21975 -45988 22102 -45972
rect 21975 -46052 22022 -45988
rect 22086 -46052 22102 -45988
rect 21975 -46068 22102 -46052
rect 21975 -46132 22022 -46068
rect 22086 -46132 22102 -46068
rect 21975 -46148 22102 -46132
rect 21975 -46212 22022 -46148
rect 22086 -46212 22102 -46148
rect 21975 -46228 22102 -46212
rect 21975 -46292 22022 -46228
rect 22086 -46292 22102 -46228
rect 21975 -46308 22102 -46292
rect 21975 -46372 22022 -46308
rect 22086 -46372 22102 -46308
rect 21975 -46388 22102 -46372
rect 21975 -46452 22022 -46388
rect 22086 -46452 22102 -46388
rect 21975 -46468 22102 -46452
rect 21975 -46532 22022 -46468
rect 22086 -46532 22102 -46468
rect 21975 -46548 22102 -46532
rect 21975 -46612 22022 -46548
rect 22086 -46612 22102 -46548
rect 21975 -46628 22102 -46612
rect 21975 -46692 22022 -46628
rect 22086 -46692 22102 -46628
rect 21975 -46708 22102 -46692
rect 21975 -46772 22022 -46708
rect 22086 -46772 22102 -46708
rect 21975 -46788 22102 -46772
rect 21975 -46852 22022 -46788
rect 22086 -46852 22102 -46788
rect 21975 -46868 22102 -46852
rect 21975 -46932 22022 -46868
rect 22086 -46932 22102 -46868
rect 21975 -46948 22102 -46932
rect 21975 -47012 22022 -46948
rect 22086 -47012 22102 -46948
rect 21975 -47028 22102 -47012
rect 15656 -47108 15783 -47092
rect 15656 -47172 15703 -47108
rect 15767 -47172 15783 -47108
rect 15656 -47188 15783 -47172
rect 15656 -47250 15760 -47188
rect 18855 -47250 18959 -47061
rect 21975 -47092 22022 -47028
rect 22086 -47092 22102 -47028
rect 22265 -41148 28187 -41139
rect 22265 -47052 22274 -41148
rect 28178 -47052 28187 -41148
rect 22265 -47061 28187 -47052
rect 28294 -41172 28341 -41108
rect 28405 -41172 28421 -41108
rect 31493 -41139 31597 -40761
rect 34613 -40792 34660 -40728
rect 34724 -40792 34740 -40728
rect 34903 -34848 40825 -34839
rect 34903 -40752 34912 -34848
rect 40816 -40752 40825 -34848
rect 34903 -40761 40825 -40752
rect 40932 -34872 40979 -34808
rect 41043 -34872 41059 -34808
rect 44131 -34839 44235 -34461
rect 47251 -34492 47298 -34428
rect 47362 -34492 47378 -34428
rect 47251 -34508 47378 -34492
rect 47251 -34572 47298 -34508
rect 47362 -34572 47378 -34508
rect 47251 -34588 47378 -34572
rect 47251 -34712 47355 -34588
rect 47251 -34728 47378 -34712
rect 47251 -34792 47298 -34728
rect 47362 -34792 47378 -34728
rect 47251 -34808 47378 -34792
rect 40932 -34888 41059 -34872
rect 40932 -34952 40979 -34888
rect 41043 -34952 41059 -34888
rect 40932 -34968 41059 -34952
rect 40932 -35032 40979 -34968
rect 41043 -35032 41059 -34968
rect 40932 -35048 41059 -35032
rect 40932 -35112 40979 -35048
rect 41043 -35112 41059 -35048
rect 40932 -35128 41059 -35112
rect 40932 -35192 40979 -35128
rect 41043 -35192 41059 -35128
rect 40932 -35208 41059 -35192
rect 40932 -35272 40979 -35208
rect 41043 -35272 41059 -35208
rect 40932 -35288 41059 -35272
rect 40932 -35352 40979 -35288
rect 41043 -35352 41059 -35288
rect 40932 -35368 41059 -35352
rect 40932 -35432 40979 -35368
rect 41043 -35432 41059 -35368
rect 40932 -35448 41059 -35432
rect 40932 -35512 40979 -35448
rect 41043 -35512 41059 -35448
rect 40932 -35528 41059 -35512
rect 40932 -35592 40979 -35528
rect 41043 -35592 41059 -35528
rect 40932 -35608 41059 -35592
rect 40932 -35672 40979 -35608
rect 41043 -35672 41059 -35608
rect 40932 -35688 41059 -35672
rect 40932 -35752 40979 -35688
rect 41043 -35752 41059 -35688
rect 40932 -35768 41059 -35752
rect 40932 -35832 40979 -35768
rect 41043 -35832 41059 -35768
rect 40932 -35848 41059 -35832
rect 40932 -35912 40979 -35848
rect 41043 -35912 41059 -35848
rect 40932 -35928 41059 -35912
rect 40932 -35992 40979 -35928
rect 41043 -35992 41059 -35928
rect 40932 -36008 41059 -35992
rect 40932 -36072 40979 -36008
rect 41043 -36072 41059 -36008
rect 40932 -36088 41059 -36072
rect 40932 -36152 40979 -36088
rect 41043 -36152 41059 -36088
rect 40932 -36168 41059 -36152
rect 40932 -36232 40979 -36168
rect 41043 -36232 41059 -36168
rect 40932 -36248 41059 -36232
rect 40932 -36312 40979 -36248
rect 41043 -36312 41059 -36248
rect 40932 -36328 41059 -36312
rect 40932 -36392 40979 -36328
rect 41043 -36392 41059 -36328
rect 40932 -36408 41059 -36392
rect 40932 -36472 40979 -36408
rect 41043 -36472 41059 -36408
rect 40932 -36488 41059 -36472
rect 40932 -36552 40979 -36488
rect 41043 -36552 41059 -36488
rect 40932 -36568 41059 -36552
rect 40932 -36632 40979 -36568
rect 41043 -36632 41059 -36568
rect 40932 -36648 41059 -36632
rect 40932 -36712 40979 -36648
rect 41043 -36712 41059 -36648
rect 40932 -36728 41059 -36712
rect 40932 -36792 40979 -36728
rect 41043 -36792 41059 -36728
rect 40932 -36808 41059 -36792
rect 40932 -36872 40979 -36808
rect 41043 -36872 41059 -36808
rect 40932 -36888 41059 -36872
rect 40932 -36952 40979 -36888
rect 41043 -36952 41059 -36888
rect 40932 -36968 41059 -36952
rect 40932 -37032 40979 -36968
rect 41043 -37032 41059 -36968
rect 40932 -37048 41059 -37032
rect 40932 -37112 40979 -37048
rect 41043 -37112 41059 -37048
rect 40932 -37128 41059 -37112
rect 40932 -37192 40979 -37128
rect 41043 -37192 41059 -37128
rect 40932 -37208 41059 -37192
rect 40932 -37272 40979 -37208
rect 41043 -37272 41059 -37208
rect 40932 -37288 41059 -37272
rect 40932 -37352 40979 -37288
rect 41043 -37352 41059 -37288
rect 40932 -37368 41059 -37352
rect 40932 -37432 40979 -37368
rect 41043 -37432 41059 -37368
rect 40932 -37448 41059 -37432
rect 40932 -37512 40979 -37448
rect 41043 -37512 41059 -37448
rect 40932 -37528 41059 -37512
rect 40932 -37592 40979 -37528
rect 41043 -37592 41059 -37528
rect 40932 -37608 41059 -37592
rect 40932 -37672 40979 -37608
rect 41043 -37672 41059 -37608
rect 40932 -37688 41059 -37672
rect 40932 -37752 40979 -37688
rect 41043 -37752 41059 -37688
rect 40932 -37768 41059 -37752
rect 40932 -37832 40979 -37768
rect 41043 -37832 41059 -37768
rect 40932 -37848 41059 -37832
rect 40932 -37912 40979 -37848
rect 41043 -37912 41059 -37848
rect 40932 -37928 41059 -37912
rect 40932 -37992 40979 -37928
rect 41043 -37992 41059 -37928
rect 40932 -38008 41059 -37992
rect 40932 -38072 40979 -38008
rect 41043 -38072 41059 -38008
rect 40932 -38088 41059 -38072
rect 40932 -38152 40979 -38088
rect 41043 -38152 41059 -38088
rect 40932 -38168 41059 -38152
rect 40932 -38232 40979 -38168
rect 41043 -38232 41059 -38168
rect 40932 -38248 41059 -38232
rect 40932 -38312 40979 -38248
rect 41043 -38312 41059 -38248
rect 40932 -38328 41059 -38312
rect 40932 -38392 40979 -38328
rect 41043 -38392 41059 -38328
rect 40932 -38408 41059 -38392
rect 40932 -38472 40979 -38408
rect 41043 -38472 41059 -38408
rect 40932 -38488 41059 -38472
rect 40932 -38552 40979 -38488
rect 41043 -38552 41059 -38488
rect 40932 -38568 41059 -38552
rect 40932 -38632 40979 -38568
rect 41043 -38632 41059 -38568
rect 40932 -38648 41059 -38632
rect 40932 -38712 40979 -38648
rect 41043 -38712 41059 -38648
rect 40932 -38728 41059 -38712
rect 40932 -38792 40979 -38728
rect 41043 -38792 41059 -38728
rect 40932 -38808 41059 -38792
rect 40932 -38872 40979 -38808
rect 41043 -38872 41059 -38808
rect 40932 -38888 41059 -38872
rect 40932 -38952 40979 -38888
rect 41043 -38952 41059 -38888
rect 40932 -38968 41059 -38952
rect 40932 -39032 40979 -38968
rect 41043 -39032 41059 -38968
rect 40932 -39048 41059 -39032
rect 40932 -39112 40979 -39048
rect 41043 -39112 41059 -39048
rect 40932 -39128 41059 -39112
rect 40932 -39192 40979 -39128
rect 41043 -39192 41059 -39128
rect 40932 -39208 41059 -39192
rect 40932 -39272 40979 -39208
rect 41043 -39272 41059 -39208
rect 40932 -39288 41059 -39272
rect 40932 -39352 40979 -39288
rect 41043 -39352 41059 -39288
rect 40932 -39368 41059 -39352
rect 40932 -39432 40979 -39368
rect 41043 -39432 41059 -39368
rect 40932 -39448 41059 -39432
rect 40932 -39512 40979 -39448
rect 41043 -39512 41059 -39448
rect 40932 -39528 41059 -39512
rect 40932 -39592 40979 -39528
rect 41043 -39592 41059 -39528
rect 40932 -39608 41059 -39592
rect 40932 -39672 40979 -39608
rect 41043 -39672 41059 -39608
rect 40932 -39688 41059 -39672
rect 40932 -39752 40979 -39688
rect 41043 -39752 41059 -39688
rect 40932 -39768 41059 -39752
rect 40932 -39832 40979 -39768
rect 41043 -39832 41059 -39768
rect 40932 -39848 41059 -39832
rect 40932 -39912 40979 -39848
rect 41043 -39912 41059 -39848
rect 40932 -39928 41059 -39912
rect 40932 -39992 40979 -39928
rect 41043 -39992 41059 -39928
rect 40932 -40008 41059 -39992
rect 40932 -40072 40979 -40008
rect 41043 -40072 41059 -40008
rect 40932 -40088 41059 -40072
rect 40932 -40152 40979 -40088
rect 41043 -40152 41059 -40088
rect 40932 -40168 41059 -40152
rect 40932 -40232 40979 -40168
rect 41043 -40232 41059 -40168
rect 40932 -40248 41059 -40232
rect 40932 -40312 40979 -40248
rect 41043 -40312 41059 -40248
rect 40932 -40328 41059 -40312
rect 40932 -40392 40979 -40328
rect 41043 -40392 41059 -40328
rect 40932 -40408 41059 -40392
rect 40932 -40472 40979 -40408
rect 41043 -40472 41059 -40408
rect 40932 -40488 41059 -40472
rect 40932 -40552 40979 -40488
rect 41043 -40552 41059 -40488
rect 40932 -40568 41059 -40552
rect 40932 -40632 40979 -40568
rect 41043 -40632 41059 -40568
rect 40932 -40648 41059 -40632
rect 40932 -40712 40979 -40648
rect 41043 -40712 41059 -40648
rect 40932 -40728 41059 -40712
rect 34613 -40808 34740 -40792
rect 34613 -40872 34660 -40808
rect 34724 -40872 34740 -40808
rect 34613 -40888 34740 -40872
rect 34613 -41012 34717 -40888
rect 34613 -41028 34740 -41012
rect 34613 -41092 34660 -41028
rect 34724 -41092 34740 -41028
rect 34613 -41108 34740 -41092
rect 28294 -41188 28421 -41172
rect 28294 -41252 28341 -41188
rect 28405 -41252 28421 -41188
rect 28294 -41268 28421 -41252
rect 28294 -41332 28341 -41268
rect 28405 -41332 28421 -41268
rect 28294 -41348 28421 -41332
rect 28294 -41412 28341 -41348
rect 28405 -41412 28421 -41348
rect 28294 -41428 28421 -41412
rect 28294 -41492 28341 -41428
rect 28405 -41492 28421 -41428
rect 28294 -41508 28421 -41492
rect 28294 -41572 28341 -41508
rect 28405 -41572 28421 -41508
rect 28294 -41588 28421 -41572
rect 28294 -41652 28341 -41588
rect 28405 -41652 28421 -41588
rect 28294 -41668 28421 -41652
rect 28294 -41732 28341 -41668
rect 28405 -41732 28421 -41668
rect 28294 -41748 28421 -41732
rect 28294 -41812 28341 -41748
rect 28405 -41812 28421 -41748
rect 28294 -41828 28421 -41812
rect 28294 -41892 28341 -41828
rect 28405 -41892 28421 -41828
rect 28294 -41908 28421 -41892
rect 28294 -41972 28341 -41908
rect 28405 -41972 28421 -41908
rect 28294 -41988 28421 -41972
rect 28294 -42052 28341 -41988
rect 28405 -42052 28421 -41988
rect 28294 -42068 28421 -42052
rect 28294 -42132 28341 -42068
rect 28405 -42132 28421 -42068
rect 28294 -42148 28421 -42132
rect 28294 -42212 28341 -42148
rect 28405 -42212 28421 -42148
rect 28294 -42228 28421 -42212
rect 28294 -42292 28341 -42228
rect 28405 -42292 28421 -42228
rect 28294 -42308 28421 -42292
rect 28294 -42372 28341 -42308
rect 28405 -42372 28421 -42308
rect 28294 -42388 28421 -42372
rect 28294 -42452 28341 -42388
rect 28405 -42452 28421 -42388
rect 28294 -42468 28421 -42452
rect 28294 -42532 28341 -42468
rect 28405 -42532 28421 -42468
rect 28294 -42548 28421 -42532
rect 28294 -42612 28341 -42548
rect 28405 -42612 28421 -42548
rect 28294 -42628 28421 -42612
rect 28294 -42692 28341 -42628
rect 28405 -42692 28421 -42628
rect 28294 -42708 28421 -42692
rect 28294 -42772 28341 -42708
rect 28405 -42772 28421 -42708
rect 28294 -42788 28421 -42772
rect 28294 -42852 28341 -42788
rect 28405 -42852 28421 -42788
rect 28294 -42868 28421 -42852
rect 28294 -42932 28341 -42868
rect 28405 -42932 28421 -42868
rect 28294 -42948 28421 -42932
rect 28294 -43012 28341 -42948
rect 28405 -43012 28421 -42948
rect 28294 -43028 28421 -43012
rect 28294 -43092 28341 -43028
rect 28405 -43092 28421 -43028
rect 28294 -43108 28421 -43092
rect 28294 -43172 28341 -43108
rect 28405 -43172 28421 -43108
rect 28294 -43188 28421 -43172
rect 28294 -43252 28341 -43188
rect 28405 -43252 28421 -43188
rect 28294 -43268 28421 -43252
rect 28294 -43332 28341 -43268
rect 28405 -43332 28421 -43268
rect 28294 -43348 28421 -43332
rect 28294 -43412 28341 -43348
rect 28405 -43412 28421 -43348
rect 28294 -43428 28421 -43412
rect 28294 -43492 28341 -43428
rect 28405 -43492 28421 -43428
rect 28294 -43508 28421 -43492
rect 28294 -43572 28341 -43508
rect 28405 -43572 28421 -43508
rect 28294 -43588 28421 -43572
rect 28294 -43652 28341 -43588
rect 28405 -43652 28421 -43588
rect 28294 -43668 28421 -43652
rect 28294 -43732 28341 -43668
rect 28405 -43732 28421 -43668
rect 28294 -43748 28421 -43732
rect 28294 -43812 28341 -43748
rect 28405 -43812 28421 -43748
rect 28294 -43828 28421 -43812
rect 28294 -43892 28341 -43828
rect 28405 -43892 28421 -43828
rect 28294 -43908 28421 -43892
rect 28294 -43972 28341 -43908
rect 28405 -43972 28421 -43908
rect 28294 -43988 28421 -43972
rect 28294 -44052 28341 -43988
rect 28405 -44052 28421 -43988
rect 28294 -44068 28421 -44052
rect 28294 -44132 28341 -44068
rect 28405 -44132 28421 -44068
rect 28294 -44148 28421 -44132
rect 28294 -44212 28341 -44148
rect 28405 -44212 28421 -44148
rect 28294 -44228 28421 -44212
rect 28294 -44292 28341 -44228
rect 28405 -44292 28421 -44228
rect 28294 -44308 28421 -44292
rect 28294 -44372 28341 -44308
rect 28405 -44372 28421 -44308
rect 28294 -44388 28421 -44372
rect 28294 -44452 28341 -44388
rect 28405 -44452 28421 -44388
rect 28294 -44468 28421 -44452
rect 28294 -44532 28341 -44468
rect 28405 -44532 28421 -44468
rect 28294 -44548 28421 -44532
rect 28294 -44612 28341 -44548
rect 28405 -44612 28421 -44548
rect 28294 -44628 28421 -44612
rect 28294 -44692 28341 -44628
rect 28405 -44692 28421 -44628
rect 28294 -44708 28421 -44692
rect 28294 -44772 28341 -44708
rect 28405 -44772 28421 -44708
rect 28294 -44788 28421 -44772
rect 28294 -44852 28341 -44788
rect 28405 -44852 28421 -44788
rect 28294 -44868 28421 -44852
rect 28294 -44932 28341 -44868
rect 28405 -44932 28421 -44868
rect 28294 -44948 28421 -44932
rect 28294 -45012 28341 -44948
rect 28405 -45012 28421 -44948
rect 28294 -45028 28421 -45012
rect 28294 -45092 28341 -45028
rect 28405 -45092 28421 -45028
rect 28294 -45108 28421 -45092
rect 28294 -45172 28341 -45108
rect 28405 -45172 28421 -45108
rect 28294 -45188 28421 -45172
rect 28294 -45252 28341 -45188
rect 28405 -45252 28421 -45188
rect 28294 -45268 28421 -45252
rect 28294 -45332 28341 -45268
rect 28405 -45332 28421 -45268
rect 28294 -45348 28421 -45332
rect 28294 -45412 28341 -45348
rect 28405 -45412 28421 -45348
rect 28294 -45428 28421 -45412
rect 28294 -45492 28341 -45428
rect 28405 -45492 28421 -45428
rect 28294 -45508 28421 -45492
rect 28294 -45572 28341 -45508
rect 28405 -45572 28421 -45508
rect 28294 -45588 28421 -45572
rect 28294 -45652 28341 -45588
rect 28405 -45652 28421 -45588
rect 28294 -45668 28421 -45652
rect 28294 -45732 28341 -45668
rect 28405 -45732 28421 -45668
rect 28294 -45748 28421 -45732
rect 28294 -45812 28341 -45748
rect 28405 -45812 28421 -45748
rect 28294 -45828 28421 -45812
rect 28294 -45892 28341 -45828
rect 28405 -45892 28421 -45828
rect 28294 -45908 28421 -45892
rect 28294 -45972 28341 -45908
rect 28405 -45972 28421 -45908
rect 28294 -45988 28421 -45972
rect 28294 -46052 28341 -45988
rect 28405 -46052 28421 -45988
rect 28294 -46068 28421 -46052
rect 28294 -46132 28341 -46068
rect 28405 -46132 28421 -46068
rect 28294 -46148 28421 -46132
rect 28294 -46212 28341 -46148
rect 28405 -46212 28421 -46148
rect 28294 -46228 28421 -46212
rect 28294 -46292 28341 -46228
rect 28405 -46292 28421 -46228
rect 28294 -46308 28421 -46292
rect 28294 -46372 28341 -46308
rect 28405 -46372 28421 -46308
rect 28294 -46388 28421 -46372
rect 28294 -46452 28341 -46388
rect 28405 -46452 28421 -46388
rect 28294 -46468 28421 -46452
rect 28294 -46532 28341 -46468
rect 28405 -46532 28421 -46468
rect 28294 -46548 28421 -46532
rect 28294 -46612 28341 -46548
rect 28405 -46612 28421 -46548
rect 28294 -46628 28421 -46612
rect 28294 -46692 28341 -46628
rect 28405 -46692 28421 -46628
rect 28294 -46708 28421 -46692
rect 28294 -46772 28341 -46708
rect 28405 -46772 28421 -46708
rect 28294 -46788 28421 -46772
rect 28294 -46852 28341 -46788
rect 28405 -46852 28421 -46788
rect 28294 -46868 28421 -46852
rect 28294 -46932 28341 -46868
rect 28405 -46932 28421 -46868
rect 28294 -46948 28421 -46932
rect 28294 -47012 28341 -46948
rect 28405 -47012 28421 -46948
rect 28294 -47028 28421 -47012
rect 21975 -47108 22102 -47092
rect 21975 -47172 22022 -47108
rect 22086 -47172 22102 -47108
rect 21975 -47188 22102 -47172
rect 21975 -47250 22079 -47188
rect 25174 -47250 25278 -47061
rect 28294 -47092 28341 -47028
rect 28405 -47092 28421 -47028
rect 28584 -41148 34506 -41139
rect 28584 -47052 28593 -41148
rect 34497 -47052 34506 -41148
rect 28584 -47061 34506 -47052
rect 34613 -41172 34660 -41108
rect 34724 -41172 34740 -41108
rect 37812 -41139 37916 -40761
rect 40932 -40792 40979 -40728
rect 41043 -40792 41059 -40728
rect 41222 -34848 47144 -34839
rect 41222 -40752 41231 -34848
rect 47135 -40752 47144 -34848
rect 41222 -40761 47144 -40752
rect 47251 -34872 47298 -34808
rect 47362 -34872 47378 -34808
rect 47251 -34888 47378 -34872
rect 47251 -34952 47298 -34888
rect 47362 -34952 47378 -34888
rect 47251 -34968 47378 -34952
rect 47251 -35032 47298 -34968
rect 47362 -35032 47378 -34968
rect 47251 -35048 47378 -35032
rect 47251 -35112 47298 -35048
rect 47362 -35112 47378 -35048
rect 47251 -35128 47378 -35112
rect 47251 -35192 47298 -35128
rect 47362 -35192 47378 -35128
rect 47251 -35208 47378 -35192
rect 47251 -35272 47298 -35208
rect 47362 -35272 47378 -35208
rect 47251 -35288 47378 -35272
rect 47251 -35352 47298 -35288
rect 47362 -35352 47378 -35288
rect 47251 -35368 47378 -35352
rect 47251 -35432 47298 -35368
rect 47362 -35432 47378 -35368
rect 47251 -35448 47378 -35432
rect 47251 -35512 47298 -35448
rect 47362 -35512 47378 -35448
rect 47251 -35528 47378 -35512
rect 47251 -35592 47298 -35528
rect 47362 -35592 47378 -35528
rect 47251 -35608 47378 -35592
rect 47251 -35672 47298 -35608
rect 47362 -35672 47378 -35608
rect 47251 -35688 47378 -35672
rect 47251 -35752 47298 -35688
rect 47362 -35752 47378 -35688
rect 47251 -35768 47378 -35752
rect 47251 -35832 47298 -35768
rect 47362 -35832 47378 -35768
rect 47251 -35848 47378 -35832
rect 47251 -35912 47298 -35848
rect 47362 -35912 47378 -35848
rect 47251 -35928 47378 -35912
rect 47251 -35992 47298 -35928
rect 47362 -35992 47378 -35928
rect 47251 -36008 47378 -35992
rect 47251 -36072 47298 -36008
rect 47362 -36072 47378 -36008
rect 47251 -36088 47378 -36072
rect 47251 -36152 47298 -36088
rect 47362 -36152 47378 -36088
rect 47251 -36168 47378 -36152
rect 47251 -36232 47298 -36168
rect 47362 -36232 47378 -36168
rect 47251 -36248 47378 -36232
rect 47251 -36312 47298 -36248
rect 47362 -36312 47378 -36248
rect 47251 -36328 47378 -36312
rect 47251 -36392 47298 -36328
rect 47362 -36392 47378 -36328
rect 47251 -36408 47378 -36392
rect 47251 -36472 47298 -36408
rect 47362 -36472 47378 -36408
rect 47251 -36488 47378 -36472
rect 47251 -36552 47298 -36488
rect 47362 -36552 47378 -36488
rect 47251 -36568 47378 -36552
rect 47251 -36632 47298 -36568
rect 47362 -36632 47378 -36568
rect 47251 -36648 47378 -36632
rect 47251 -36712 47298 -36648
rect 47362 -36712 47378 -36648
rect 47251 -36728 47378 -36712
rect 47251 -36792 47298 -36728
rect 47362 -36792 47378 -36728
rect 47251 -36808 47378 -36792
rect 47251 -36872 47298 -36808
rect 47362 -36872 47378 -36808
rect 47251 -36888 47378 -36872
rect 47251 -36952 47298 -36888
rect 47362 -36952 47378 -36888
rect 47251 -36968 47378 -36952
rect 47251 -37032 47298 -36968
rect 47362 -37032 47378 -36968
rect 47251 -37048 47378 -37032
rect 47251 -37112 47298 -37048
rect 47362 -37112 47378 -37048
rect 47251 -37128 47378 -37112
rect 47251 -37192 47298 -37128
rect 47362 -37192 47378 -37128
rect 47251 -37208 47378 -37192
rect 47251 -37272 47298 -37208
rect 47362 -37272 47378 -37208
rect 47251 -37288 47378 -37272
rect 47251 -37352 47298 -37288
rect 47362 -37352 47378 -37288
rect 47251 -37368 47378 -37352
rect 47251 -37432 47298 -37368
rect 47362 -37432 47378 -37368
rect 47251 -37448 47378 -37432
rect 47251 -37512 47298 -37448
rect 47362 -37512 47378 -37448
rect 47251 -37528 47378 -37512
rect 47251 -37592 47298 -37528
rect 47362 -37592 47378 -37528
rect 47251 -37608 47378 -37592
rect 47251 -37672 47298 -37608
rect 47362 -37672 47378 -37608
rect 47251 -37688 47378 -37672
rect 47251 -37752 47298 -37688
rect 47362 -37752 47378 -37688
rect 47251 -37768 47378 -37752
rect 47251 -37832 47298 -37768
rect 47362 -37832 47378 -37768
rect 47251 -37848 47378 -37832
rect 47251 -37912 47298 -37848
rect 47362 -37912 47378 -37848
rect 47251 -37928 47378 -37912
rect 47251 -37992 47298 -37928
rect 47362 -37992 47378 -37928
rect 47251 -38008 47378 -37992
rect 47251 -38072 47298 -38008
rect 47362 -38072 47378 -38008
rect 47251 -38088 47378 -38072
rect 47251 -38152 47298 -38088
rect 47362 -38152 47378 -38088
rect 47251 -38168 47378 -38152
rect 47251 -38232 47298 -38168
rect 47362 -38232 47378 -38168
rect 47251 -38248 47378 -38232
rect 47251 -38312 47298 -38248
rect 47362 -38312 47378 -38248
rect 47251 -38328 47378 -38312
rect 47251 -38392 47298 -38328
rect 47362 -38392 47378 -38328
rect 47251 -38408 47378 -38392
rect 47251 -38472 47298 -38408
rect 47362 -38472 47378 -38408
rect 47251 -38488 47378 -38472
rect 47251 -38552 47298 -38488
rect 47362 -38552 47378 -38488
rect 47251 -38568 47378 -38552
rect 47251 -38632 47298 -38568
rect 47362 -38632 47378 -38568
rect 47251 -38648 47378 -38632
rect 47251 -38712 47298 -38648
rect 47362 -38712 47378 -38648
rect 47251 -38728 47378 -38712
rect 47251 -38792 47298 -38728
rect 47362 -38792 47378 -38728
rect 47251 -38808 47378 -38792
rect 47251 -38872 47298 -38808
rect 47362 -38872 47378 -38808
rect 47251 -38888 47378 -38872
rect 47251 -38952 47298 -38888
rect 47362 -38952 47378 -38888
rect 47251 -38968 47378 -38952
rect 47251 -39032 47298 -38968
rect 47362 -39032 47378 -38968
rect 47251 -39048 47378 -39032
rect 47251 -39112 47298 -39048
rect 47362 -39112 47378 -39048
rect 47251 -39128 47378 -39112
rect 47251 -39192 47298 -39128
rect 47362 -39192 47378 -39128
rect 47251 -39208 47378 -39192
rect 47251 -39272 47298 -39208
rect 47362 -39272 47378 -39208
rect 47251 -39288 47378 -39272
rect 47251 -39352 47298 -39288
rect 47362 -39352 47378 -39288
rect 47251 -39368 47378 -39352
rect 47251 -39432 47298 -39368
rect 47362 -39432 47378 -39368
rect 47251 -39448 47378 -39432
rect 47251 -39512 47298 -39448
rect 47362 -39512 47378 -39448
rect 47251 -39528 47378 -39512
rect 47251 -39592 47298 -39528
rect 47362 -39592 47378 -39528
rect 47251 -39608 47378 -39592
rect 47251 -39672 47298 -39608
rect 47362 -39672 47378 -39608
rect 47251 -39688 47378 -39672
rect 47251 -39752 47298 -39688
rect 47362 -39752 47378 -39688
rect 47251 -39768 47378 -39752
rect 47251 -39832 47298 -39768
rect 47362 -39832 47378 -39768
rect 47251 -39848 47378 -39832
rect 47251 -39912 47298 -39848
rect 47362 -39912 47378 -39848
rect 47251 -39928 47378 -39912
rect 47251 -39992 47298 -39928
rect 47362 -39992 47378 -39928
rect 47251 -40008 47378 -39992
rect 47251 -40072 47298 -40008
rect 47362 -40072 47378 -40008
rect 47251 -40088 47378 -40072
rect 47251 -40152 47298 -40088
rect 47362 -40152 47378 -40088
rect 47251 -40168 47378 -40152
rect 47251 -40232 47298 -40168
rect 47362 -40232 47378 -40168
rect 47251 -40248 47378 -40232
rect 47251 -40312 47298 -40248
rect 47362 -40312 47378 -40248
rect 47251 -40328 47378 -40312
rect 47251 -40392 47298 -40328
rect 47362 -40392 47378 -40328
rect 47251 -40408 47378 -40392
rect 47251 -40472 47298 -40408
rect 47362 -40472 47378 -40408
rect 47251 -40488 47378 -40472
rect 47251 -40552 47298 -40488
rect 47362 -40552 47378 -40488
rect 47251 -40568 47378 -40552
rect 47251 -40632 47298 -40568
rect 47362 -40632 47378 -40568
rect 47251 -40648 47378 -40632
rect 47251 -40712 47298 -40648
rect 47362 -40712 47378 -40648
rect 47251 -40728 47378 -40712
rect 40932 -40808 41059 -40792
rect 40932 -40872 40979 -40808
rect 41043 -40872 41059 -40808
rect 40932 -40888 41059 -40872
rect 40932 -41012 41036 -40888
rect 40932 -41028 41059 -41012
rect 40932 -41092 40979 -41028
rect 41043 -41092 41059 -41028
rect 40932 -41108 41059 -41092
rect 34613 -41188 34740 -41172
rect 34613 -41252 34660 -41188
rect 34724 -41252 34740 -41188
rect 34613 -41268 34740 -41252
rect 34613 -41332 34660 -41268
rect 34724 -41332 34740 -41268
rect 34613 -41348 34740 -41332
rect 34613 -41412 34660 -41348
rect 34724 -41412 34740 -41348
rect 34613 -41428 34740 -41412
rect 34613 -41492 34660 -41428
rect 34724 -41492 34740 -41428
rect 34613 -41508 34740 -41492
rect 34613 -41572 34660 -41508
rect 34724 -41572 34740 -41508
rect 34613 -41588 34740 -41572
rect 34613 -41652 34660 -41588
rect 34724 -41652 34740 -41588
rect 34613 -41668 34740 -41652
rect 34613 -41732 34660 -41668
rect 34724 -41732 34740 -41668
rect 34613 -41748 34740 -41732
rect 34613 -41812 34660 -41748
rect 34724 -41812 34740 -41748
rect 34613 -41828 34740 -41812
rect 34613 -41892 34660 -41828
rect 34724 -41892 34740 -41828
rect 34613 -41908 34740 -41892
rect 34613 -41972 34660 -41908
rect 34724 -41972 34740 -41908
rect 34613 -41988 34740 -41972
rect 34613 -42052 34660 -41988
rect 34724 -42052 34740 -41988
rect 34613 -42068 34740 -42052
rect 34613 -42132 34660 -42068
rect 34724 -42132 34740 -42068
rect 34613 -42148 34740 -42132
rect 34613 -42212 34660 -42148
rect 34724 -42212 34740 -42148
rect 34613 -42228 34740 -42212
rect 34613 -42292 34660 -42228
rect 34724 -42292 34740 -42228
rect 34613 -42308 34740 -42292
rect 34613 -42372 34660 -42308
rect 34724 -42372 34740 -42308
rect 34613 -42388 34740 -42372
rect 34613 -42452 34660 -42388
rect 34724 -42452 34740 -42388
rect 34613 -42468 34740 -42452
rect 34613 -42532 34660 -42468
rect 34724 -42532 34740 -42468
rect 34613 -42548 34740 -42532
rect 34613 -42612 34660 -42548
rect 34724 -42612 34740 -42548
rect 34613 -42628 34740 -42612
rect 34613 -42692 34660 -42628
rect 34724 -42692 34740 -42628
rect 34613 -42708 34740 -42692
rect 34613 -42772 34660 -42708
rect 34724 -42772 34740 -42708
rect 34613 -42788 34740 -42772
rect 34613 -42852 34660 -42788
rect 34724 -42852 34740 -42788
rect 34613 -42868 34740 -42852
rect 34613 -42932 34660 -42868
rect 34724 -42932 34740 -42868
rect 34613 -42948 34740 -42932
rect 34613 -43012 34660 -42948
rect 34724 -43012 34740 -42948
rect 34613 -43028 34740 -43012
rect 34613 -43092 34660 -43028
rect 34724 -43092 34740 -43028
rect 34613 -43108 34740 -43092
rect 34613 -43172 34660 -43108
rect 34724 -43172 34740 -43108
rect 34613 -43188 34740 -43172
rect 34613 -43252 34660 -43188
rect 34724 -43252 34740 -43188
rect 34613 -43268 34740 -43252
rect 34613 -43332 34660 -43268
rect 34724 -43332 34740 -43268
rect 34613 -43348 34740 -43332
rect 34613 -43412 34660 -43348
rect 34724 -43412 34740 -43348
rect 34613 -43428 34740 -43412
rect 34613 -43492 34660 -43428
rect 34724 -43492 34740 -43428
rect 34613 -43508 34740 -43492
rect 34613 -43572 34660 -43508
rect 34724 -43572 34740 -43508
rect 34613 -43588 34740 -43572
rect 34613 -43652 34660 -43588
rect 34724 -43652 34740 -43588
rect 34613 -43668 34740 -43652
rect 34613 -43732 34660 -43668
rect 34724 -43732 34740 -43668
rect 34613 -43748 34740 -43732
rect 34613 -43812 34660 -43748
rect 34724 -43812 34740 -43748
rect 34613 -43828 34740 -43812
rect 34613 -43892 34660 -43828
rect 34724 -43892 34740 -43828
rect 34613 -43908 34740 -43892
rect 34613 -43972 34660 -43908
rect 34724 -43972 34740 -43908
rect 34613 -43988 34740 -43972
rect 34613 -44052 34660 -43988
rect 34724 -44052 34740 -43988
rect 34613 -44068 34740 -44052
rect 34613 -44132 34660 -44068
rect 34724 -44132 34740 -44068
rect 34613 -44148 34740 -44132
rect 34613 -44212 34660 -44148
rect 34724 -44212 34740 -44148
rect 34613 -44228 34740 -44212
rect 34613 -44292 34660 -44228
rect 34724 -44292 34740 -44228
rect 34613 -44308 34740 -44292
rect 34613 -44372 34660 -44308
rect 34724 -44372 34740 -44308
rect 34613 -44388 34740 -44372
rect 34613 -44452 34660 -44388
rect 34724 -44452 34740 -44388
rect 34613 -44468 34740 -44452
rect 34613 -44532 34660 -44468
rect 34724 -44532 34740 -44468
rect 34613 -44548 34740 -44532
rect 34613 -44612 34660 -44548
rect 34724 -44612 34740 -44548
rect 34613 -44628 34740 -44612
rect 34613 -44692 34660 -44628
rect 34724 -44692 34740 -44628
rect 34613 -44708 34740 -44692
rect 34613 -44772 34660 -44708
rect 34724 -44772 34740 -44708
rect 34613 -44788 34740 -44772
rect 34613 -44852 34660 -44788
rect 34724 -44852 34740 -44788
rect 34613 -44868 34740 -44852
rect 34613 -44932 34660 -44868
rect 34724 -44932 34740 -44868
rect 34613 -44948 34740 -44932
rect 34613 -45012 34660 -44948
rect 34724 -45012 34740 -44948
rect 34613 -45028 34740 -45012
rect 34613 -45092 34660 -45028
rect 34724 -45092 34740 -45028
rect 34613 -45108 34740 -45092
rect 34613 -45172 34660 -45108
rect 34724 -45172 34740 -45108
rect 34613 -45188 34740 -45172
rect 34613 -45252 34660 -45188
rect 34724 -45252 34740 -45188
rect 34613 -45268 34740 -45252
rect 34613 -45332 34660 -45268
rect 34724 -45332 34740 -45268
rect 34613 -45348 34740 -45332
rect 34613 -45412 34660 -45348
rect 34724 -45412 34740 -45348
rect 34613 -45428 34740 -45412
rect 34613 -45492 34660 -45428
rect 34724 -45492 34740 -45428
rect 34613 -45508 34740 -45492
rect 34613 -45572 34660 -45508
rect 34724 -45572 34740 -45508
rect 34613 -45588 34740 -45572
rect 34613 -45652 34660 -45588
rect 34724 -45652 34740 -45588
rect 34613 -45668 34740 -45652
rect 34613 -45732 34660 -45668
rect 34724 -45732 34740 -45668
rect 34613 -45748 34740 -45732
rect 34613 -45812 34660 -45748
rect 34724 -45812 34740 -45748
rect 34613 -45828 34740 -45812
rect 34613 -45892 34660 -45828
rect 34724 -45892 34740 -45828
rect 34613 -45908 34740 -45892
rect 34613 -45972 34660 -45908
rect 34724 -45972 34740 -45908
rect 34613 -45988 34740 -45972
rect 34613 -46052 34660 -45988
rect 34724 -46052 34740 -45988
rect 34613 -46068 34740 -46052
rect 34613 -46132 34660 -46068
rect 34724 -46132 34740 -46068
rect 34613 -46148 34740 -46132
rect 34613 -46212 34660 -46148
rect 34724 -46212 34740 -46148
rect 34613 -46228 34740 -46212
rect 34613 -46292 34660 -46228
rect 34724 -46292 34740 -46228
rect 34613 -46308 34740 -46292
rect 34613 -46372 34660 -46308
rect 34724 -46372 34740 -46308
rect 34613 -46388 34740 -46372
rect 34613 -46452 34660 -46388
rect 34724 -46452 34740 -46388
rect 34613 -46468 34740 -46452
rect 34613 -46532 34660 -46468
rect 34724 -46532 34740 -46468
rect 34613 -46548 34740 -46532
rect 34613 -46612 34660 -46548
rect 34724 -46612 34740 -46548
rect 34613 -46628 34740 -46612
rect 34613 -46692 34660 -46628
rect 34724 -46692 34740 -46628
rect 34613 -46708 34740 -46692
rect 34613 -46772 34660 -46708
rect 34724 -46772 34740 -46708
rect 34613 -46788 34740 -46772
rect 34613 -46852 34660 -46788
rect 34724 -46852 34740 -46788
rect 34613 -46868 34740 -46852
rect 34613 -46932 34660 -46868
rect 34724 -46932 34740 -46868
rect 34613 -46948 34740 -46932
rect 34613 -47012 34660 -46948
rect 34724 -47012 34740 -46948
rect 34613 -47028 34740 -47012
rect 28294 -47108 28421 -47092
rect 28294 -47172 28341 -47108
rect 28405 -47172 28421 -47108
rect 28294 -47188 28421 -47172
rect 28294 -47250 28398 -47188
rect 31493 -47250 31597 -47061
rect 34613 -47092 34660 -47028
rect 34724 -47092 34740 -47028
rect 34903 -41148 40825 -41139
rect 34903 -47052 34912 -41148
rect 40816 -47052 40825 -41148
rect 34903 -47061 40825 -47052
rect 40932 -41172 40979 -41108
rect 41043 -41172 41059 -41108
rect 44131 -41139 44235 -40761
rect 47251 -40792 47298 -40728
rect 47362 -40792 47378 -40728
rect 47251 -40808 47378 -40792
rect 47251 -40872 47298 -40808
rect 47362 -40872 47378 -40808
rect 47251 -40888 47378 -40872
rect 47251 -41012 47355 -40888
rect 47251 -41028 47378 -41012
rect 47251 -41092 47298 -41028
rect 47362 -41092 47378 -41028
rect 47251 -41108 47378 -41092
rect 40932 -41188 41059 -41172
rect 40932 -41252 40979 -41188
rect 41043 -41252 41059 -41188
rect 40932 -41268 41059 -41252
rect 40932 -41332 40979 -41268
rect 41043 -41332 41059 -41268
rect 40932 -41348 41059 -41332
rect 40932 -41412 40979 -41348
rect 41043 -41412 41059 -41348
rect 40932 -41428 41059 -41412
rect 40932 -41492 40979 -41428
rect 41043 -41492 41059 -41428
rect 40932 -41508 41059 -41492
rect 40932 -41572 40979 -41508
rect 41043 -41572 41059 -41508
rect 40932 -41588 41059 -41572
rect 40932 -41652 40979 -41588
rect 41043 -41652 41059 -41588
rect 40932 -41668 41059 -41652
rect 40932 -41732 40979 -41668
rect 41043 -41732 41059 -41668
rect 40932 -41748 41059 -41732
rect 40932 -41812 40979 -41748
rect 41043 -41812 41059 -41748
rect 40932 -41828 41059 -41812
rect 40932 -41892 40979 -41828
rect 41043 -41892 41059 -41828
rect 40932 -41908 41059 -41892
rect 40932 -41972 40979 -41908
rect 41043 -41972 41059 -41908
rect 40932 -41988 41059 -41972
rect 40932 -42052 40979 -41988
rect 41043 -42052 41059 -41988
rect 40932 -42068 41059 -42052
rect 40932 -42132 40979 -42068
rect 41043 -42132 41059 -42068
rect 40932 -42148 41059 -42132
rect 40932 -42212 40979 -42148
rect 41043 -42212 41059 -42148
rect 40932 -42228 41059 -42212
rect 40932 -42292 40979 -42228
rect 41043 -42292 41059 -42228
rect 40932 -42308 41059 -42292
rect 40932 -42372 40979 -42308
rect 41043 -42372 41059 -42308
rect 40932 -42388 41059 -42372
rect 40932 -42452 40979 -42388
rect 41043 -42452 41059 -42388
rect 40932 -42468 41059 -42452
rect 40932 -42532 40979 -42468
rect 41043 -42532 41059 -42468
rect 40932 -42548 41059 -42532
rect 40932 -42612 40979 -42548
rect 41043 -42612 41059 -42548
rect 40932 -42628 41059 -42612
rect 40932 -42692 40979 -42628
rect 41043 -42692 41059 -42628
rect 40932 -42708 41059 -42692
rect 40932 -42772 40979 -42708
rect 41043 -42772 41059 -42708
rect 40932 -42788 41059 -42772
rect 40932 -42852 40979 -42788
rect 41043 -42852 41059 -42788
rect 40932 -42868 41059 -42852
rect 40932 -42932 40979 -42868
rect 41043 -42932 41059 -42868
rect 40932 -42948 41059 -42932
rect 40932 -43012 40979 -42948
rect 41043 -43012 41059 -42948
rect 40932 -43028 41059 -43012
rect 40932 -43092 40979 -43028
rect 41043 -43092 41059 -43028
rect 40932 -43108 41059 -43092
rect 40932 -43172 40979 -43108
rect 41043 -43172 41059 -43108
rect 40932 -43188 41059 -43172
rect 40932 -43252 40979 -43188
rect 41043 -43252 41059 -43188
rect 40932 -43268 41059 -43252
rect 40932 -43332 40979 -43268
rect 41043 -43332 41059 -43268
rect 40932 -43348 41059 -43332
rect 40932 -43412 40979 -43348
rect 41043 -43412 41059 -43348
rect 40932 -43428 41059 -43412
rect 40932 -43492 40979 -43428
rect 41043 -43492 41059 -43428
rect 40932 -43508 41059 -43492
rect 40932 -43572 40979 -43508
rect 41043 -43572 41059 -43508
rect 40932 -43588 41059 -43572
rect 40932 -43652 40979 -43588
rect 41043 -43652 41059 -43588
rect 40932 -43668 41059 -43652
rect 40932 -43732 40979 -43668
rect 41043 -43732 41059 -43668
rect 40932 -43748 41059 -43732
rect 40932 -43812 40979 -43748
rect 41043 -43812 41059 -43748
rect 40932 -43828 41059 -43812
rect 40932 -43892 40979 -43828
rect 41043 -43892 41059 -43828
rect 40932 -43908 41059 -43892
rect 40932 -43972 40979 -43908
rect 41043 -43972 41059 -43908
rect 40932 -43988 41059 -43972
rect 40932 -44052 40979 -43988
rect 41043 -44052 41059 -43988
rect 40932 -44068 41059 -44052
rect 40932 -44132 40979 -44068
rect 41043 -44132 41059 -44068
rect 40932 -44148 41059 -44132
rect 40932 -44212 40979 -44148
rect 41043 -44212 41059 -44148
rect 40932 -44228 41059 -44212
rect 40932 -44292 40979 -44228
rect 41043 -44292 41059 -44228
rect 40932 -44308 41059 -44292
rect 40932 -44372 40979 -44308
rect 41043 -44372 41059 -44308
rect 40932 -44388 41059 -44372
rect 40932 -44452 40979 -44388
rect 41043 -44452 41059 -44388
rect 40932 -44468 41059 -44452
rect 40932 -44532 40979 -44468
rect 41043 -44532 41059 -44468
rect 40932 -44548 41059 -44532
rect 40932 -44612 40979 -44548
rect 41043 -44612 41059 -44548
rect 40932 -44628 41059 -44612
rect 40932 -44692 40979 -44628
rect 41043 -44692 41059 -44628
rect 40932 -44708 41059 -44692
rect 40932 -44772 40979 -44708
rect 41043 -44772 41059 -44708
rect 40932 -44788 41059 -44772
rect 40932 -44852 40979 -44788
rect 41043 -44852 41059 -44788
rect 40932 -44868 41059 -44852
rect 40932 -44932 40979 -44868
rect 41043 -44932 41059 -44868
rect 40932 -44948 41059 -44932
rect 40932 -45012 40979 -44948
rect 41043 -45012 41059 -44948
rect 40932 -45028 41059 -45012
rect 40932 -45092 40979 -45028
rect 41043 -45092 41059 -45028
rect 40932 -45108 41059 -45092
rect 40932 -45172 40979 -45108
rect 41043 -45172 41059 -45108
rect 40932 -45188 41059 -45172
rect 40932 -45252 40979 -45188
rect 41043 -45252 41059 -45188
rect 40932 -45268 41059 -45252
rect 40932 -45332 40979 -45268
rect 41043 -45332 41059 -45268
rect 40932 -45348 41059 -45332
rect 40932 -45412 40979 -45348
rect 41043 -45412 41059 -45348
rect 40932 -45428 41059 -45412
rect 40932 -45492 40979 -45428
rect 41043 -45492 41059 -45428
rect 40932 -45508 41059 -45492
rect 40932 -45572 40979 -45508
rect 41043 -45572 41059 -45508
rect 40932 -45588 41059 -45572
rect 40932 -45652 40979 -45588
rect 41043 -45652 41059 -45588
rect 40932 -45668 41059 -45652
rect 40932 -45732 40979 -45668
rect 41043 -45732 41059 -45668
rect 40932 -45748 41059 -45732
rect 40932 -45812 40979 -45748
rect 41043 -45812 41059 -45748
rect 40932 -45828 41059 -45812
rect 40932 -45892 40979 -45828
rect 41043 -45892 41059 -45828
rect 40932 -45908 41059 -45892
rect 40932 -45972 40979 -45908
rect 41043 -45972 41059 -45908
rect 40932 -45988 41059 -45972
rect 40932 -46052 40979 -45988
rect 41043 -46052 41059 -45988
rect 40932 -46068 41059 -46052
rect 40932 -46132 40979 -46068
rect 41043 -46132 41059 -46068
rect 40932 -46148 41059 -46132
rect 40932 -46212 40979 -46148
rect 41043 -46212 41059 -46148
rect 40932 -46228 41059 -46212
rect 40932 -46292 40979 -46228
rect 41043 -46292 41059 -46228
rect 40932 -46308 41059 -46292
rect 40932 -46372 40979 -46308
rect 41043 -46372 41059 -46308
rect 40932 -46388 41059 -46372
rect 40932 -46452 40979 -46388
rect 41043 -46452 41059 -46388
rect 40932 -46468 41059 -46452
rect 40932 -46532 40979 -46468
rect 41043 -46532 41059 -46468
rect 40932 -46548 41059 -46532
rect 40932 -46612 40979 -46548
rect 41043 -46612 41059 -46548
rect 40932 -46628 41059 -46612
rect 40932 -46692 40979 -46628
rect 41043 -46692 41059 -46628
rect 40932 -46708 41059 -46692
rect 40932 -46772 40979 -46708
rect 41043 -46772 41059 -46708
rect 40932 -46788 41059 -46772
rect 40932 -46852 40979 -46788
rect 41043 -46852 41059 -46788
rect 40932 -46868 41059 -46852
rect 40932 -46932 40979 -46868
rect 41043 -46932 41059 -46868
rect 40932 -46948 41059 -46932
rect 40932 -47012 40979 -46948
rect 41043 -47012 41059 -46948
rect 40932 -47028 41059 -47012
rect 34613 -47108 34740 -47092
rect 34613 -47172 34660 -47108
rect 34724 -47172 34740 -47108
rect 34613 -47188 34740 -47172
rect 34613 -47250 34717 -47188
rect 37812 -47250 37916 -47061
rect 40932 -47092 40979 -47028
rect 41043 -47092 41059 -47028
rect 41222 -41148 47144 -41139
rect 41222 -47052 41231 -41148
rect 47135 -47052 47144 -41148
rect 41222 -47061 47144 -47052
rect 47251 -41172 47298 -41108
rect 47362 -41172 47378 -41108
rect 47251 -41188 47378 -41172
rect 47251 -41252 47298 -41188
rect 47362 -41252 47378 -41188
rect 47251 -41268 47378 -41252
rect 47251 -41332 47298 -41268
rect 47362 -41332 47378 -41268
rect 47251 -41348 47378 -41332
rect 47251 -41412 47298 -41348
rect 47362 -41412 47378 -41348
rect 47251 -41428 47378 -41412
rect 47251 -41492 47298 -41428
rect 47362 -41492 47378 -41428
rect 47251 -41508 47378 -41492
rect 47251 -41572 47298 -41508
rect 47362 -41572 47378 -41508
rect 47251 -41588 47378 -41572
rect 47251 -41652 47298 -41588
rect 47362 -41652 47378 -41588
rect 47251 -41668 47378 -41652
rect 47251 -41732 47298 -41668
rect 47362 -41732 47378 -41668
rect 47251 -41748 47378 -41732
rect 47251 -41812 47298 -41748
rect 47362 -41812 47378 -41748
rect 47251 -41828 47378 -41812
rect 47251 -41892 47298 -41828
rect 47362 -41892 47378 -41828
rect 47251 -41908 47378 -41892
rect 47251 -41972 47298 -41908
rect 47362 -41972 47378 -41908
rect 47251 -41988 47378 -41972
rect 47251 -42052 47298 -41988
rect 47362 -42052 47378 -41988
rect 47251 -42068 47378 -42052
rect 47251 -42132 47298 -42068
rect 47362 -42132 47378 -42068
rect 47251 -42148 47378 -42132
rect 47251 -42212 47298 -42148
rect 47362 -42212 47378 -42148
rect 47251 -42228 47378 -42212
rect 47251 -42292 47298 -42228
rect 47362 -42292 47378 -42228
rect 47251 -42308 47378 -42292
rect 47251 -42372 47298 -42308
rect 47362 -42372 47378 -42308
rect 47251 -42388 47378 -42372
rect 47251 -42452 47298 -42388
rect 47362 -42452 47378 -42388
rect 47251 -42468 47378 -42452
rect 47251 -42532 47298 -42468
rect 47362 -42532 47378 -42468
rect 47251 -42548 47378 -42532
rect 47251 -42612 47298 -42548
rect 47362 -42612 47378 -42548
rect 47251 -42628 47378 -42612
rect 47251 -42692 47298 -42628
rect 47362 -42692 47378 -42628
rect 47251 -42708 47378 -42692
rect 47251 -42772 47298 -42708
rect 47362 -42772 47378 -42708
rect 47251 -42788 47378 -42772
rect 47251 -42852 47298 -42788
rect 47362 -42852 47378 -42788
rect 47251 -42868 47378 -42852
rect 47251 -42932 47298 -42868
rect 47362 -42932 47378 -42868
rect 47251 -42948 47378 -42932
rect 47251 -43012 47298 -42948
rect 47362 -43012 47378 -42948
rect 47251 -43028 47378 -43012
rect 47251 -43092 47298 -43028
rect 47362 -43092 47378 -43028
rect 47251 -43108 47378 -43092
rect 47251 -43172 47298 -43108
rect 47362 -43172 47378 -43108
rect 47251 -43188 47378 -43172
rect 47251 -43252 47298 -43188
rect 47362 -43252 47378 -43188
rect 47251 -43268 47378 -43252
rect 47251 -43332 47298 -43268
rect 47362 -43332 47378 -43268
rect 47251 -43348 47378 -43332
rect 47251 -43412 47298 -43348
rect 47362 -43412 47378 -43348
rect 47251 -43428 47378 -43412
rect 47251 -43492 47298 -43428
rect 47362 -43492 47378 -43428
rect 47251 -43508 47378 -43492
rect 47251 -43572 47298 -43508
rect 47362 -43572 47378 -43508
rect 47251 -43588 47378 -43572
rect 47251 -43652 47298 -43588
rect 47362 -43652 47378 -43588
rect 47251 -43668 47378 -43652
rect 47251 -43732 47298 -43668
rect 47362 -43732 47378 -43668
rect 47251 -43748 47378 -43732
rect 47251 -43812 47298 -43748
rect 47362 -43812 47378 -43748
rect 47251 -43828 47378 -43812
rect 47251 -43892 47298 -43828
rect 47362 -43892 47378 -43828
rect 47251 -43908 47378 -43892
rect 47251 -43972 47298 -43908
rect 47362 -43972 47378 -43908
rect 47251 -43988 47378 -43972
rect 47251 -44052 47298 -43988
rect 47362 -44052 47378 -43988
rect 47251 -44068 47378 -44052
rect 47251 -44132 47298 -44068
rect 47362 -44132 47378 -44068
rect 47251 -44148 47378 -44132
rect 47251 -44212 47298 -44148
rect 47362 -44212 47378 -44148
rect 47251 -44228 47378 -44212
rect 47251 -44292 47298 -44228
rect 47362 -44292 47378 -44228
rect 47251 -44308 47378 -44292
rect 47251 -44372 47298 -44308
rect 47362 -44372 47378 -44308
rect 47251 -44388 47378 -44372
rect 47251 -44452 47298 -44388
rect 47362 -44452 47378 -44388
rect 47251 -44468 47378 -44452
rect 47251 -44532 47298 -44468
rect 47362 -44532 47378 -44468
rect 47251 -44548 47378 -44532
rect 47251 -44612 47298 -44548
rect 47362 -44612 47378 -44548
rect 47251 -44628 47378 -44612
rect 47251 -44692 47298 -44628
rect 47362 -44692 47378 -44628
rect 47251 -44708 47378 -44692
rect 47251 -44772 47298 -44708
rect 47362 -44772 47378 -44708
rect 47251 -44788 47378 -44772
rect 47251 -44852 47298 -44788
rect 47362 -44852 47378 -44788
rect 47251 -44868 47378 -44852
rect 47251 -44932 47298 -44868
rect 47362 -44932 47378 -44868
rect 47251 -44948 47378 -44932
rect 47251 -45012 47298 -44948
rect 47362 -45012 47378 -44948
rect 47251 -45028 47378 -45012
rect 47251 -45092 47298 -45028
rect 47362 -45092 47378 -45028
rect 47251 -45108 47378 -45092
rect 47251 -45172 47298 -45108
rect 47362 -45172 47378 -45108
rect 47251 -45188 47378 -45172
rect 47251 -45252 47298 -45188
rect 47362 -45252 47378 -45188
rect 47251 -45268 47378 -45252
rect 47251 -45332 47298 -45268
rect 47362 -45332 47378 -45268
rect 47251 -45348 47378 -45332
rect 47251 -45412 47298 -45348
rect 47362 -45412 47378 -45348
rect 47251 -45428 47378 -45412
rect 47251 -45492 47298 -45428
rect 47362 -45492 47378 -45428
rect 47251 -45508 47378 -45492
rect 47251 -45572 47298 -45508
rect 47362 -45572 47378 -45508
rect 47251 -45588 47378 -45572
rect 47251 -45652 47298 -45588
rect 47362 -45652 47378 -45588
rect 47251 -45668 47378 -45652
rect 47251 -45732 47298 -45668
rect 47362 -45732 47378 -45668
rect 47251 -45748 47378 -45732
rect 47251 -45812 47298 -45748
rect 47362 -45812 47378 -45748
rect 47251 -45828 47378 -45812
rect 47251 -45892 47298 -45828
rect 47362 -45892 47378 -45828
rect 47251 -45908 47378 -45892
rect 47251 -45972 47298 -45908
rect 47362 -45972 47378 -45908
rect 47251 -45988 47378 -45972
rect 47251 -46052 47298 -45988
rect 47362 -46052 47378 -45988
rect 47251 -46068 47378 -46052
rect 47251 -46132 47298 -46068
rect 47362 -46132 47378 -46068
rect 47251 -46148 47378 -46132
rect 47251 -46212 47298 -46148
rect 47362 -46212 47378 -46148
rect 47251 -46228 47378 -46212
rect 47251 -46292 47298 -46228
rect 47362 -46292 47378 -46228
rect 47251 -46308 47378 -46292
rect 47251 -46372 47298 -46308
rect 47362 -46372 47378 -46308
rect 47251 -46388 47378 -46372
rect 47251 -46452 47298 -46388
rect 47362 -46452 47378 -46388
rect 47251 -46468 47378 -46452
rect 47251 -46532 47298 -46468
rect 47362 -46532 47378 -46468
rect 47251 -46548 47378 -46532
rect 47251 -46612 47298 -46548
rect 47362 -46612 47378 -46548
rect 47251 -46628 47378 -46612
rect 47251 -46692 47298 -46628
rect 47362 -46692 47378 -46628
rect 47251 -46708 47378 -46692
rect 47251 -46772 47298 -46708
rect 47362 -46772 47378 -46708
rect 47251 -46788 47378 -46772
rect 47251 -46852 47298 -46788
rect 47362 -46852 47378 -46788
rect 47251 -46868 47378 -46852
rect 47251 -46932 47298 -46868
rect 47362 -46932 47378 -46868
rect 47251 -46948 47378 -46932
rect 47251 -47012 47298 -46948
rect 47362 -47012 47378 -46948
rect 47251 -47028 47378 -47012
rect 40932 -47108 41059 -47092
rect 40932 -47172 40979 -47108
rect 41043 -47172 41059 -47108
rect 40932 -47188 41059 -47172
rect 40932 -47250 41036 -47188
rect 44131 -47250 44235 -47061
rect 47251 -47092 47298 -47028
rect 47362 -47092 47378 -47028
rect 47251 -47108 47378 -47092
rect 47251 -47172 47298 -47108
rect 47362 -47172 47378 -47108
rect 47251 -47188 47378 -47172
rect 47251 -47250 47355 -47188
<< properties >>
string FIXED_BBOX 41083 41000 47283 47200
<< end >>
