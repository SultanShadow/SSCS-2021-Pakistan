magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< error_p >>
rect -31 5081 31 5087
rect -31 5047 -17 5081
rect -31 5041 31 5047
rect -31 -5047 31 -5041
rect -31 -5081 -17 -5047
rect -31 -5087 31 -5081
<< nwell >>
rect -231 -5219 231 5219
<< pmoslvt >>
rect -35 -5000 35 5000
<< pdiff >>
rect -93 4981 -35 5000
rect -93 4947 -81 4981
rect -47 4947 -35 4981
rect -93 4913 -35 4947
rect -93 4879 -81 4913
rect -47 4879 -35 4913
rect -93 4845 -35 4879
rect -93 4811 -81 4845
rect -47 4811 -35 4845
rect -93 4777 -35 4811
rect -93 4743 -81 4777
rect -47 4743 -35 4777
rect -93 4709 -35 4743
rect -93 4675 -81 4709
rect -47 4675 -35 4709
rect -93 4641 -35 4675
rect -93 4607 -81 4641
rect -47 4607 -35 4641
rect -93 4573 -35 4607
rect -93 4539 -81 4573
rect -47 4539 -35 4573
rect -93 4505 -35 4539
rect -93 4471 -81 4505
rect -47 4471 -35 4505
rect -93 4437 -35 4471
rect -93 4403 -81 4437
rect -47 4403 -35 4437
rect -93 4369 -35 4403
rect -93 4335 -81 4369
rect -47 4335 -35 4369
rect -93 4301 -35 4335
rect -93 4267 -81 4301
rect -47 4267 -35 4301
rect -93 4233 -35 4267
rect -93 4199 -81 4233
rect -47 4199 -35 4233
rect -93 4165 -35 4199
rect -93 4131 -81 4165
rect -47 4131 -35 4165
rect -93 4097 -35 4131
rect -93 4063 -81 4097
rect -47 4063 -35 4097
rect -93 4029 -35 4063
rect -93 3995 -81 4029
rect -47 3995 -35 4029
rect -93 3961 -35 3995
rect -93 3927 -81 3961
rect -47 3927 -35 3961
rect -93 3893 -35 3927
rect -93 3859 -81 3893
rect -47 3859 -35 3893
rect -93 3825 -35 3859
rect -93 3791 -81 3825
rect -47 3791 -35 3825
rect -93 3757 -35 3791
rect -93 3723 -81 3757
rect -47 3723 -35 3757
rect -93 3689 -35 3723
rect -93 3655 -81 3689
rect -47 3655 -35 3689
rect -93 3621 -35 3655
rect -93 3587 -81 3621
rect -47 3587 -35 3621
rect -93 3553 -35 3587
rect -93 3519 -81 3553
rect -47 3519 -35 3553
rect -93 3485 -35 3519
rect -93 3451 -81 3485
rect -47 3451 -35 3485
rect -93 3417 -35 3451
rect -93 3383 -81 3417
rect -47 3383 -35 3417
rect -93 3349 -35 3383
rect -93 3315 -81 3349
rect -47 3315 -35 3349
rect -93 3281 -35 3315
rect -93 3247 -81 3281
rect -47 3247 -35 3281
rect -93 3213 -35 3247
rect -93 3179 -81 3213
rect -47 3179 -35 3213
rect -93 3145 -35 3179
rect -93 3111 -81 3145
rect -47 3111 -35 3145
rect -93 3077 -35 3111
rect -93 3043 -81 3077
rect -47 3043 -35 3077
rect -93 3009 -35 3043
rect -93 2975 -81 3009
rect -47 2975 -35 3009
rect -93 2941 -35 2975
rect -93 2907 -81 2941
rect -47 2907 -35 2941
rect -93 2873 -35 2907
rect -93 2839 -81 2873
rect -47 2839 -35 2873
rect -93 2805 -35 2839
rect -93 2771 -81 2805
rect -47 2771 -35 2805
rect -93 2737 -35 2771
rect -93 2703 -81 2737
rect -47 2703 -35 2737
rect -93 2669 -35 2703
rect -93 2635 -81 2669
rect -47 2635 -35 2669
rect -93 2601 -35 2635
rect -93 2567 -81 2601
rect -47 2567 -35 2601
rect -93 2533 -35 2567
rect -93 2499 -81 2533
rect -47 2499 -35 2533
rect -93 2465 -35 2499
rect -93 2431 -81 2465
rect -47 2431 -35 2465
rect -93 2397 -35 2431
rect -93 2363 -81 2397
rect -47 2363 -35 2397
rect -93 2329 -35 2363
rect -93 2295 -81 2329
rect -47 2295 -35 2329
rect -93 2261 -35 2295
rect -93 2227 -81 2261
rect -47 2227 -35 2261
rect -93 2193 -35 2227
rect -93 2159 -81 2193
rect -47 2159 -35 2193
rect -93 2125 -35 2159
rect -93 2091 -81 2125
rect -47 2091 -35 2125
rect -93 2057 -35 2091
rect -93 2023 -81 2057
rect -47 2023 -35 2057
rect -93 1989 -35 2023
rect -93 1955 -81 1989
rect -47 1955 -35 1989
rect -93 1921 -35 1955
rect -93 1887 -81 1921
rect -47 1887 -35 1921
rect -93 1853 -35 1887
rect -93 1819 -81 1853
rect -47 1819 -35 1853
rect -93 1785 -35 1819
rect -93 1751 -81 1785
rect -47 1751 -35 1785
rect -93 1717 -35 1751
rect -93 1683 -81 1717
rect -47 1683 -35 1717
rect -93 1649 -35 1683
rect -93 1615 -81 1649
rect -47 1615 -35 1649
rect -93 1581 -35 1615
rect -93 1547 -81 1581
rect -47 1547 -35 1581
rect -93 1513 -35 1547
rect -93 1479 -81 1513
rect -47 1479 -35 1513
rect -93 1445 -35 1479
rect -93 1411 -81 1445
rect -47 1411 -35 1445
rect -93 1377 -35 1411
rect -93 1343 -81 1377
rect -47 1343 -35 1377
rect -93 1309 -35 1343
rect -93 1275 -81 1309
rect -47 1275 -35 1309
rect -93 1241 -35 1275
rect -93 1207 -81 1241
rect -47 1207 -35 1241
rect -93 1173 -35 1207
rect -93 1139 -81 1173
rect -47 1139 -35 1173
rect -93 1105 -35 1139
rect -93 1071 -81 1105
rect -47 1071 -35 1105
rect -93 1037 -35 1071
rect -93 1003 -81 1037
rect -47 1003 -35 1037
rect -93 969 -35 1003
rect -93 935 -81 969
rect -47 935 -35 969
rect -93 901 -35 935
rect -93 867 -81 901
rect -47 867 -35 901
rect -93 833 -35 867
rect -93 799 -81 833
rect -47 799 -35 833
rect -93 765 -35 799
rect -93 731 -81 765
rect -47 731 -35 765
rect -93 697 -35 731
rect -93 663 -81 697
rect -47 663 -35 697
rect -93 629 -35 663
rect -93 595 -81 629
rect -47 595 -35 629
rect -93 561 -35 595
rect -93 527 -81 561
rect -47 527 -35 561
rect -93 493 -35 527
rect -93 459 -81 493
rect -47 459 -35 493
rect -93 425 -35 459
rect -93 391 -81 425
rect -47 391 -35 425
rect -93 357 -35 391
rect -93 323 -81 357
rect -47 323 -35 357
rect -93 289 -35 323
rect -93 255 -81 289
rect -47 255 -35 289
rect -93 221 -35 255
rect -93 187 -81 221
rect -47 187 -35 221
rect -93 153 -35 187
rect -93 119 -81 153
rect -47 119 -35 153
rect -93 85 -35 119
rect -93 51 -81 85
rect -47 51 -35 85
rect -93 17 -35 51
rect -93 -17 -81 17
rect -47 -17 -35 17
rect -93 -51 -35 -17
rect -93 -85 -81 -51
rect -47 -85 -35 -51
rect -93 -119 -35 -85
rect -93 -153 -81 -119
rect -47 -153 -35 -119
rect -93 -187 -35 -153
rect -93 -221 -81 -187
rect -47 -221 -35 -187
rect -93 -255 -35 -221
rect -93 -289 -81 -255
rect -47 -289 -35 -255
rect -93 -323 -35 -289
rect -93 -357 -81 -323
rect -47 -357 -35 -323
rect -93 -391 -35 -357
rect -93 -425 -81 -391
rect -47 -425 -35 -391
rect -93 -459 -35 -425
rect -93 -493 -81 -459
rect -47 -493 -35 -459
rect -93 -527 -35 -493
rect -93 -561 -81 -527
rect -47 -561 -35 -527
rect -93 -595 -35 -561
rect -93 -629 -81 -595
rect -47 -629 -35 -595
rect -93 -663 -35 -629
rect -93 -697 -81 -663
rect -47 -697 -35 -663
rect -93 -731 -35 -697
rect -93 -765 -81 -731
rect -47 -765 -35 -731
rect -93 -799 -35 -765
rect -93 -833 -81 -799
rect -47 -833 -35 -799
rect -93 -867 -35 -833
rect -93 -901 -81 -867
rect -47 -901 -35 -867
rect -93 -935 -35 -901
rect -93 -969 -81 -935
rect -47 -969 -35 -935
rect -93 -1003 -35 -969
rect -93 -1037 -81 -1003
rect -47 -1037 -35 -1003
rect -93 -1071 -35 -1037
rect -93 -1105 -81 -1071
rect -47 -1105 -35 -1071
rect -93 -1139 -35 -1105
rect -93 -1173 -81 -1139
rect -47 -1173 -35 -1139
rect -93 -1207 -35 -1173
rect -93 -1241 -81 -1207
rect -47 -1241 -35 -1207
rect -93 -1275 -35 -1241
rect -93 -1309 -81 -1275
rect -47 -1309 -35 -1275
rect -93 -1343 -35 -1309
rect -93 -1377 -81 -1343
rect -47 -1377 -35 -1343
rect -93 -1411 -35 -1377
rect -93 -1445 -81 -1411
rect -47 -1445 -35 -1411
rect -93 -1479 -35 -1445
rect -93 -1513 -81 -1479
rect -47 -1513 -35 -1479
rect -93 -1547 -35 -1513
rect -93 -1581 -81 -1547
rect -47 -1581 -35 -1547
rect -93 -1615 -35 -1581
rect -93 -1649 -81 -1615
rect -47 -1649 -35 -1615
rect -93 -1683 -35 -1649
rect -93 -1717 -81 -1683
rect -47 -1717 -35 -1683
rect -93 -1751 -35 -1717
rect -93 -1785 -81 -1751
rect -47 -1785 -35 -1751
rect -93 -1819 -35 -1785
rect -93 -1853 -81 -1819
rect -47 -1853 -35 -1819
rect -93 -1887 -35 -1853
rect -93 -1921 -81 -1887
rect -47 -1921 -35 -1887
rect -93 -1955 -35 -1921
rect -93 -1989 -81 -1955
rect -47 -1989 -35 -1955
rect -93 -2023 -35 -1989
rect -93 -2057 -81 -2023
rect -47 -2057 -35 -2023
rect -93 -2091 -35 -2057
rect -93 -2125 -81 -2091
rect -47 -2125 -35 -2091
rect -93 -2159 -35 -2125
rect -93 -2193 -81 -2159
rect -47 -2193 -35 -2159
rect -93 -2227 -35 -2193
rect -93 -2261 -81 -2227
rect -47 -2261 -35 -2227
rect -93 -2295 -35 -2261
rect -93 -2329 -81 -2295
rect -47 -2329 -35 -2295
rect -93 -2363 -35 -2329
rect -93 -2397 -81 -2363
rect -47 -2397 -35 -2363
rect -93 -2431 -35 -2397
rect -93 -2465 -81 -2431
rect -47 -2465 -35 -2431
rect -93 -2499 -35 -2465
rect -93 -2533 -81 -2499
rect -47 -2533 -35 -2499
rect -93 -2567 -35 -2533
rect -93 -2601 -81 -2567
rect -47 -2601 -35 -2567
rect -93 -2635 -35 -2601
rect -93 -2669 -81 -2635
rect -47 -2669 -35 -2635
rect -93 -2703 -35 -2669
rect -93 -2737 -81 -2703
rect -47 -2737 -35 -2703
rect -93 -2771 -35 -2737
rect -93 -2805 -81 -2771
rect -47 -2805 -35 -2771
rect -93 -2839 -35 -2805
rect -93 -2873 -81 -2839
rect -47 -2873 -35 -2839
rect -93 -2907 -35 -2873
rect -93 -2941 -81 -2907
rect -47 -2941 -35 -2907
rect -93 -2975 -35 -2941
rect -93 -3009 -81 -2975
rect -47 -3009 -35 -2975
rect -93 -3043 -35 -3009
rect -93 -3077 -81 -3043
rect -47 -3077 -35 -3043
rect -93 -3111 -35 -3077
rect -93 -3145 -81 -3111
rect -47 -3145 -35 -3111
rect -93 -3179 -35 -3145
rect -93 -3213 -81 -3179
rect -47 -3213 -35 -3179
rect -93 -3247 -35 -3213
rect -93 -3281 -81 -3247
rect -47 -3281 -35 -3247
rect -93 -3315 -35 -3281
rect -93 -3349 -81 -3315
rect -47 -3349 -35 -3315
rect -93 -3383 -35 -3349
rect -93 -3417 -81 -3383
rect -47 -3417 -35 -3383
rect -93 -3451 -35 -3417
rect -93 -3485 -81 -3451
rect -47 -3485 -35 -3451
rect -93 -3519 -35 -3485
rect -93 -3553 -81 -3519
rect -47 -3553 -35 -3519
rect -93 -3587 -35 -3553
rect -93 -3621 -81 -3587
rect -47 -3621 -35 -3587
rect -93 -3655 -35 -3621
rect -93 -3689 -81 -3655
rect -47 -3689 -35 -3655
rect -93 -3723 -35 -3689
rect -93 -3757 -81 -3723
rect -47 -3757 -35 -3723
rect -93 -3791 -35 -3757
rect -93 -3825 -81 -3791
rect -47 -3825 -35 -3791
rect -93 -3859 -35 -3825
rect -93 -3893 -81 -3859
rect -47 -3893 -35 -3859
rect -93 -3927 -35 -3893
rect -93 -3961 -81 -3927
rect -47 -3961 -35 -3927
rect -93 -3995 -35 -3961
rect -93 -4029 -81 -3995
rect -47 -4029 -35 -3995
rect -93 -4063 -35 -4029
rect -93 -4097 -81 -4063
rect -47 -4097 -35 -4063
rect -93 -4131 -35 -4097
rect -93 -4165 -81 -4131
rect -47 -4165 -35 -4131
rect -93 -4199 -35 -4165
rect -93 -4233 -81 -4199
rect -47 -4233 -35 -4199
rect -93 -4267 -35 -4233
rect -93 -4301 -81 -4267
rect -47 -4301 -35 -4267
rect -93 -4335 -35 -4301
rect -93 -4369 -81 -4335
rect -47 -4369 -35 -4335
rect -93 -4403 -35 -4369
rect -93 -4437 -81 -4403
rect -47 -4437 -35 -4403
rect -93 -4471 -35 -4437
rect -93 -4505 -81 -4471
rect -47 -4505 -35 -4471
rect -93 -4539 -35 -4505
rect -93 -4573 -81 -4539
rect -47 -4573 -35 -4539
rect -93 -4607 -35 -4573
rect -93 -4641 -81 -4607
rect -47 -4641 -35 -4607
rect -93 -4675 -35 -4641
rect -93 -4709 -81 -4675
rect -47 -4709 -35 -4675
rect -93 -4743 -35 -4709
rect -93 -4777 -81 -4743
rect -47 -4777 -35 -4743
rect -93 -4811 -35 -4777
rect -93 -4845 -81 -4811
rect -47 -4845 -35 -4811
rect -93 -4879 -35 -4845
rect -93 -4913 -81 -4879
rect -47 -4913 -35 -4879
rect -93 -4947 -35 -4913
rect -93 -4981 -81 -4947
rect -47 -4981 -35 -4947
rect -93 -5000 -35 -4981
rect 35 4981 93 5000
rect 35 4947 47 4981
rect 81 4947 93 4981
rect 35 4913 93 4947
rect 35 4879 47 4913
rect 81 4879 93 4913
rect 35 4845 93 4879
rect 35 4811 47 4845
rect 81 4811 93 4845
rect 35 4777 93 4811
rect 35 4743 47 4777
rect 81 4743 93 4777
rect 35 4709 93 4743
rect 35 4675 47 4709
rect 81 4675 93 4709
rect 35 4641 93 4675
rect 35 4607 47 4641
rect 81 4607 93 4641
rect 35 4573 93 4607
rect 35 4539 47 4573
rect 81 4539 93 4573
rect 35 4505 93 4539
rect 35 4471 47 4505
rect 81 4471 93 4505
rect 35 4437 93 4471
rect 35 4403 47 4437
rect 81 4403 93 4437
rect 35 4369 93 4403
rect 35 4335 47 4369
rect 81 4335 93 4369
rect 35 4301 93 4335
rect 35 4267 47 4301
rect 81 4267 93 4301
rect 35 4233 93 4267
rect 35 4199 47 4233
rect 81 4199 93 4233
rect 35 4165 93 4199
rect 35 4131 47 4165
rect 81 4131 93 4165
rect 35 4097 93 4131
rect 35 4063 47 4097
rect 81 4063 93 4097
rect 35 4029 93 4063
rect 35 3995 47 4029
rect 81 3995 93 4029
rect 35 3961 93 3995
rect 35 3927 47 3961
rect 81 3927 93 3961
rect 35 3893 93 3927
rect 35 3859 47 3893
rect 81 3859 93 3893
rect 35 3825 93 3859
rect 35 3791 47 3825
rect 81 3791 93 3825
rect 35 3757 93 3791
rect 35 3723 47 3757
rect 81 3723 93 3757
rect 35 3689 93 3723
rect 35 3655 47 3689
rect 81 3655 93 3689
rect 35 3621 93 3655
rect 35 3587 47 3621
rect 81 3587 93 3621
rect 35 3553 93 3587
rect 35 3519 47 3553
rect 81 3519 93 3553
rect 35 3485 93 3519
rect 35 3451 47 3485
rect 81 3451 93 3485
rect 35 3417 93 3451
rect 35 3383 47 3417
rect 81 3383 93 3417
rect 35 3349 93 3383
rect 35 3315 47 3349
rect 81 3315 93 3349
rect 35 3281 93 3315
rect 35 3247 47 3281
rect 81 3247 93 3281
rect 35 3213 93 3247
rect 35 3179 47 3213
rect 81 3179 93 3213
rect 35 3145 93 3179
rect 35 3111 47 3145
rect 81 3111 93 3145
rect 35 3077 93 3111
rect 35 3043 47 3077
rect 81 3043 93 3077
rect 35 3009 93 3043
rect 35 2975 47 3009
rect 81 2975 93 3009
rect 35 2941 93 2975
rect 35 2907 47 2941
rect 81 2907 93 2941
rect 35 2873 93 2907
rect 35 2839 47 2873
rect 81 2839 93 2873
rect 35 2805 93 2839
rect 35 2771 47 2805
rect 81 2771 93 2805
rect 35 2737 93 2771
rect 35 2703 47 2737
rect 81 2703 93 2737
rect 35 2669 93 2703
rect 35 2635 47 2669
rect 81 2635 93 2669
rect 35 2601 93 2635
rect 35 2567 47 2601
rect 81 2567 93 2601
rect 35 2533 93 2567
rect 35 2499 47 2533
rect 81 2499 93 2533
rect 35 2465 93 2499
rect 35 2431 47 2465
rect 81 2431 93 2465
rect 35 2397 93 2431
rect 35 2363 47 2397
rect 81 2363 93 2397
rect 35 2329 93 2363
rect 35 2295 47 2329
rect 81 2295 93 2329
rect 35 2261 93 2295
rect 35 2227 47 2261
rect 81 2227 93 2261
rect 35 2193 93 2227
rect 35 2159 47 2193
rect 81 2159 93 2193
rect 35 2125 93 2159
rect 35 2091 47 2125
rect 81 2091 93 2125
rect 35 2057 93 2091
rect 35 2023 47 2057
rect 81 2023 93 2057
rect 35 1989 93 2023
rect 35 1955 47 1989
rect 81 1955 93 1989
rect 35 1921 93 1955
rect 35 1887 47 1921
rect 81 1887 93 1921
rect 35 1853 93 1887
rect 35 1819 47 1853
rect 81 1819 93 1853
rect 35 1785 93 1819
rect 35 1751 47 1785
rect 81 1751 93 1785
rect 35 1717 93 1751
rect 35 1683 47 1717
rect 81 1683 93 1717
rect 35 1649 93 1683
rect 35 1615 47 1649
rect 81 1615 93 1649
rect 35 1581 93 1615
rect 35 1547 47 1581
rect 81 1547 93 1581
rect 35 1513 93 1547
rect 35 1479 47 1513
rect 81 1479 93 1513
rect 35 1445 93 1479
rect 35 1411 47 1445
rect 81 1411 93 1445
rect 35 1377 93 1411
rect 35 1343 47 1377
rect 81 1343 93 1377
rect 35 1309 93 1343
rect 35 1275 47 1309
rect 81 1275 93 1309
rect 35 1241 93 1275
rect 35 1207 47 1241
rect 81 1207 93 1241
rect 35 1173 93 1207
rect 35 1139 47 1173
rect 81 1139 93 1173
rect 35 1105 93 1139
rect 35 1071 47 1105
rect 81 1071 93 1105
rect 35 1037 93 1071
rect 35 1003 47 1037
rect 81 1003 93 1037
rect 35 969 93 1003
rect 35 935 47 969
rect 81 935 93 969
rect 35 901 93 935
rect 35 867 47 901
rect 81 867 93 901
rect 35 833 93 867
rect 35 799 47 833
rect 81 799 93 833
rect 35 765 93 799
rect 35 731 47 765
rect 81 731 93 765
rect 35 697 93 731
rect 35 663 47 697
rect 81 663 93 697
rect 35 629 93 663
rect 35 595 47 629
rect 81 595 93 629
rect 35 561 93 595
rect 35 527 47 561
rect 81 527 93 561
rect 35 493 93 527
rect 35 459 47 493
rect 81 459 93 493
rect 35 425 93 459
rect 35 391 47 425
rect 81 391 93 425
rect 35 357 93 391
rect 35 323 47 357
rect 81 323 93 357
rect 35 289 93 323
rect 35 255 47 289
rect 81 255 93 289
rect 35 221 93 255
rect 35 187 47 221
rect 81 187 93 221
rect 35 153 93 187
rect 35 119 47 153
rect 81 119 93 153
rect 35 85 93 119
rect 35 51 47 85
rect 81 51 93 85
rect 35 17 93 51
rect 35 -17 47 17
rect 81 -17 93 17
rect 35 -51 93 -17
rect 35 -85 47 -51
rect 81 -85 93 -51
rect 35 -119 93 -85
rect 35 -153 47 -119
rect 81 -153 93 -119
rect 35 -187 93 -153
rect 35 -221 47 -187
rect 81 -221 93 -187
rect 35 -255 93 -221
rect 35 -289 47 -255
rect 81 -289 93 -255
rect 35 -323 93 -289
rect 35 -357 47 -323
rect 81 -357 93 -323
rect 35 -391 93 -357
rect 35 -425 47 -391
rect 81 -425 93 -391
rect 35 -459 93 -425
rect 35 -493 47 -459
rect 81 -493 93 -459
rect 35 -527 93 -493
rect 35 -561 47 -527
rect 81 -561 93 -527
rect 35 -595 93 -561
rect 35 -629 47 -595
rect 81 -629 93 -595
rect 35 -663 93 -629
rect 35 -697 47 -663
rect 81 -697 93 -663
rect 35 -731 93 -697
rect 35 -765 47 -731
rect 81 -765 93 -731
rect 35 -799 93 -765
rect 35 -833 47 -799
rect 81 -833 93 -799
rect 35 -867 93 -833
rect 35 -901 47 -867
rect 81 -901 93 -867
rect 35 -935 93 -901
rect 35 -969 47 -935
rect 81 -969 93 -935
rect 35 -1003 93 -969
rect 35 -1037 47 -1003
rect 81 -1037 93 -1003
rect 35 -1071 93 -1037
rect 35 -1105 47 -1071
rect 81 -1105 93 -1071
rect 35 -1139 93 -1105
rect 35 -1173 47 -1139
rect 81 -1173 93 -1139
rect 35 -1207 93 -1173
rect 35 -1241 47 -1207
rect 81 -1241 93 -1207
rect 35 -1275 93 -1241
rect 35 -1309 47 -1275
rect 81 -1309 93 -1275
rect 35 -1343 93 -1309
rect 35 -1377 47 -1343
rect 81 -1377 93 -1343
rect 35 -1411 93 -1377
rect 35 -1445 47 -1411
rect 81 -1445 93 -1411
rect 35 -1479 93 -1445
rect 35 -1513 47 -1479
rect 81 -1513 93 -1479
rect 35 -1547 93 -1513
rect 35 -1581 47 -1547
rect 81 -1581 93 -1547
rect 35 -1615 93 -1581
rect 35 -1649 47 -1615
rect 81 -1649 93 -1615
rect 35 -1683 93 -1649
rect 35 -1717 47 -1683
rect 81 -1717 93 -1683
rect 35 -1751 93 -1717
rect 35 -1785 47 -1751
rect 81 -1785 93 -1751
rect 35 -1819 93 -1785
rect 35 -1853 47 -1819
rect 81 -1853 93 -1819
rect 35 -1887 93 -1853
rect 35 -1921 47 -1887
rect 81 -1921 93 -1887
rect 35 -1955 93 -1921
rect 35 -1989 47 -1955
rect 81 -1989 93 -1955
rect 35 -2023 93 -1989
rect 35 -2057 47 -2023
rect 81 -2057 93 -2023
rect 35 -2091 93 -2057
rect 35 -2125 47 -2091
rect 81 -2125 93 -2091
rect 35 -2159 93 -2125
rect 35 -2193 47 -2159
rect 81 -2193 93 -2159
rect 35 -2227 93 -2193
rect 35 -2261 47 -2227
rect 81 -2261 93 -2227
rect 35 -2295 93 -2261
rect 35 -2329 47 -2295
rect 81 -2329 93 -2295
rect 35 -2363 93 -2329
rect 35 -2397 47 -2363
rect 81 -2397 93 -2363
rect 35 -2431 93 -2397
rect 35 -2465 47 -2431
rect 81 -2465 93 -2431
rect 35 -2499 93 -2465
rect 35 -2533 47 -2499
rect 81 -2533 93 -2499
rect 35 -2567 93 -2533
rect 35 -2601 47 -2567
rect 81 -2601 93 -2567
rect 35 -2635 93 -2601
rect 35 -2669 47 -2635
rect 81 -2669 93 -2635
rect 35 -2703 93 -2669
rect 35 -2737 47 -2703
rect 81 -2737 93 -2703
rect 35 -2771 93 -2737
rect 35 -2805 47 -2771
rect 81 -2805 93 -2771
rect 35 -2839 93 -2805
rect 35 -2873 47 -2839
rect 81 -2873 93 -2839
rect 35 -2907 93 -2873
rect 35 -2941 47 -2907
rect 81 -2941 93 -2907
rect 35 -2975 93 -2941
rect 35 -3009 47 -2975
rect 81 -3009 93 -2975
rect 35 -3043 93 -3009
rect 35 -3077 47 -3043
rect 81 -3077 93 -3043
rect 35 -3111 93 -3077
rect 35 -3145 47 -3111
rect 81 -3145 93 -3111
rect 35 -3179 93 -3145
rect 35 -3213 47 -3179
rect 81 -3213 93 -3179
rect 35 -3247 93 -3213
rect 35 -3281 47 -3247
rect 81 -3281 93 -3247
rect 35 -3315 93 -3281
rect 35 -3349 47 -3315
rect 81 -3349 93 -3315
rect 35 -3383 93 -3349
rect 35 -3417 47 -3383
rect 81 -3417 93 -3383
rect 35 -3451 93 -3417
rect 35 -3485 47 -3451
rect 81 -3485 93 -3451
rect 35 -3519 93 -3485
rect 35 -3553 47 -3519
rect 81 -3553 93 -3519
rect 35 -3587 93 -3553
rect 35 -3621 47 -3587
rect 81 -3621 93 -3587
rect 35 -3655 93 -3621
rect 35 -3689 47 -3655
rect 81 -3689 93 -3655
rect 35 -3723 93 -3689
rect 35 -3757 47 -3723
rect 81 -3757 93 -3723
rect 35 -3791 93 -3757
rect 35 -3825 47 -3791
rect 81 -3825 93 -3791
rect 35 -3859 93 -3825
rect 35 -3893 47 -3859
rect 81 -3893 93 -3859
rect 35 -3927 93 -3893
rect 35 -3961 47 -3927
rect 81 -3961 93 -3927
rect 35 -3995 93 -3961
rect 35 -4029 47 -3995
rect 81 -4029 93 -3995
rect 35 -4063 93 -4029
rect 35 -4097 47 -4063
rect 81 -4097 93 -4063
rect 35 -4131 93 -4097
rect 35 -4165 47 -4131
rect 81 -4165 93 -4131
rect 35 -4199 93 -4165
rect 35 -4233 47 -4199
rect 81 -4233 93 -4199
rect 35 -4267 93 -4233
rect 35 -4301 47 -4267
rect 81 -4301 93 -4267
rect 35 -4335 93 -4301
rect 35 -4369 47 -4335
rect 81 -4369 93 -4335
rect 35 -4403 93 -4369
rect 35 -4437 47 -4403
rect 81 -4437 93 -4403
rect 35 -4471 93 -4437
rect 35 -4505 47 -4471
rect 81 -4505 93 -4471
rect 35 -4539 93 -4505
rect 35 -4573 47 -4539
rect 81 -4573 93 -4539
rect 35 -4607 93 -4573
rect 35 -4641 47 -4607
rect 81 -4641 93 -4607
rect 35 -4675 93 -4641
rect 35 -4709 47 -4675
rect 81 -4709 93 -4675
rect 35 -4743 93 -4709
rect 35 -4777 47 -4743
rect 81 -4777 93 -4743
rect 35 -4811 93 -4777
rect 35 -4845 47 -4811
rect 81 -4845 93 -4811
rect 35 -4879 93 -4845
rect 35 -4913 47 -4879
rect 81 -4913 93 -4879
rect 35 -4947 93 -4913
rect 35 -4981 47 -4947
rect 81 -4981 93 -4947
rect 35 -5000 93 -4981
<< pdiffc >>
rect -81 4947 -47 4981
rect -81 4879 -47 4913
rect -81 4811 -47 4845
rect -81 4743 -47 4777
rect -81 4675 -47 4709
rect -81 4607 -47 4641
rect -81 4539 -47 4573
rect -81 4471 -47 4505
rect -81 4403 -47 4437
rect -81 4335 -47 4369
rect -81 4267 -47 4301
rect -81 4199 -47 4233
rect -81 4131 -47 4165
rect -81 4063 -47 4097
rect -81 3995 -47 4029
rect -81 3927 -47 3961
rect -81 3859 -47 3893
rect -81 3791 -47 3825
rect -81 3723 -47 3757
rect -81 3655 -47 3689
rect -81 3587 -47 3621
rect -81 3519 -47 3553
rect -81 3451 -47 3485
rect -81 3383 -47 3417
rect -81 3315 -47 3349
rect -81 3247 -47 3281
rect -81 3179 -47 3213
rect -81 3111 -47 3145
rect -81 3043 -47 3077
rect -81 2975 -47 3009
rect -81 2907 -47 2941
rect -81 2839 -47 2873
rect -81 2771 -47 2805
rect -81 2703 -47 2737
rect -81 2635 -47 2669
rect -81 2567 -47 2601
rect -81 2499 -47 2533
rect -81 2431 -47 2465
rect -81 2363 -47 2397
rect -81 2295 -47 2329
rect -81 2227 -47 2261
rect -81 2159 -47 2193
rect -81 2091 -47 2125
rect -81 2023 -47 2057
rect -81 1955 -47 1989
rect -81 1887 -47 1921
rect -81 1819 -47 1853
rect -81 1751 -47 1785
rect -81 1683 -47 1717
rect -81 1615 -47 1649
rect -81 1547 -47 1581
rect -81 1479 -47 1513
rect -81 1411 -47 1445
rect -81 1343 -47 1377
rect -81 1275 -47 1309
rect -81 1207 -47 1241
rect -81 1139 -47 1173
rect -81 1071 -47 1105
rect -81 1003 -47 1037
rect -81 935 -47 969
rect -81 867 -47 901
rect -81 799 -47 833
rect -81 731 -47 765
rect -81 663 -47 697
rect -81 595 -47 629
rect -81 527 -47 561
rect -81 459 -47 493
rect -81 391 -47 425
rect -81 323 -47 357
rect -81 255 -47 289
rect -81 187 -47 221
rect -81 119 -47 153
rect -81 51 -47 85
rect -81 -17 -47 17
rect -81 -85 -47 -51
rect -81 -153 -47 -119
rect -81 -221 -47 -187
rect -81 -289 -47 -255
rect -81 -357 -47 -323
rect -81 -425 -47 -391
rect -81 -493 -47 -459
rect -81 -561 -47 -527
rect -81 -629 -47 -595
rect -81 -697 -47 -663
rect -81 -765 -47 -731
rect -81 -833 -47 -799
rect -81 -901 -47 -867
rect -81 -969 -47 -935
rect -81 -1037 -47 -1003
rect -81 -1105 -47 -1071
rect -81 -1173 -47 -1139
rect -81 -1241 -47 -1207
rect -81 -1309 -47 -1275
rect -81 -1377 -47 -1343
rect -81 -1445 -47 -1411
rect -81 -1513 -47 -1479
rect -81 -1581 -47 -1547
rect -81 -1649 -47 -1615
rect -81 -1717 -47 -1683
rect -81 -1785 -47 -1751
rect -81 -1853 -47 -1819
rect -81 -1921 -47 -1887
rect -81 -1989 -47 -1955
rect -81 -2057 -47 -2023
rect -81 -2125 -47 -2091
rect -81 -2193 -47 -2159
rect -81 -2261 -47 -2227
rect -81 -2329 -47 -2295
rect -81 -2397 -47 -2363
rect -81 -2465 -47 -2431
rect -81 -2533 -47 -2499
rect -81 -2601 -47 -2567
rect -81 -2669 -47 -2635
rect -81 -2737 -47 -2703
rect -81 -2805 -47 -2771
rect -81 -2873 -47 -2839
rect -81 -2941 -47 -2907
rect -81 -3009 -47 -2975
rect -81 -3077 -47 -3043
rect -81 -3145 -47 -3111
rect -81 -3213 -47 -3179
rect -81 -3281 -47 -3247
rect -81 -3349 -47 -3315
rect -81 -3417 -47 -3383
rect -81 -3485 -47 -3451
rect -81 -3553 -47 -3519
rect -81 -3621 -47 -3587
rect -81 -3689 -47 -3655
rect -81 -3757 -47 -3723
rect -81 -3825 -47 -3791
rect -81 -3893 -47 -3859
rect -81 -3961 -47 -3927
rect -81 -4029 -47 -3995
rect -81 -4097 -47 -4063
rect -81 -4165 -47 -4131
rect -81 -4233 -47 -4199
rect -81 -4301 -47 -4267
rect -81 -4369 -47 -4335
rect -81 -4437 -47 -4403
rect -81 -4505 -47 -4471
rect -81 -4573 -47 -4539
rect -81 -4641 -47 -4607
rect -81 -4709 -47 -4675
rect -81 -4777 -47 -4743
rect -81 -4845 -47 -4811
rect -81 -4913 -47 -4879
rect -81 -4981 -47 -4947
rect 47 4947 81 4981
rect 47 4879 81 4913
rect 47 4811 81 4845
rect 47 4743 81 4777
rect 47 4675 81 4709
rect 47 4607 81 4641
rect 47 4539 81 4573
rect 47 4471 81 4505
rect 47 4403 81 4437
rect 47 4335 81 4369
rect 47 4267 81 4301
rect 47 4199 81 4233
rect 47 4131 81 4165
rect 47 4063 81 4097
rect 47 3995 81 4029
rect 47 3927 81 3961
rect 47 3859 81 3893
rect 47 3791 81 3825
rect 47 3723 81 3757
rect 47 3655 81 3689
rect 47 3587 81 3621
rect 47 3519 81 3553
rect 47 3451 81 3485
rect 47 3383 81 3417
rect 47 3315 81 3349
rect 47 3247 81 3281
rect 47 3179 81 3213
rect 47 3111 81 3145
rect 47 3043 81 3077
rect 47 2975 81 3009
rect 47 2907 81 2941
rect 47 2839 81 2873
rect 47 2771 81 2805
rect 47 2703 81 2737
rect 47 2635 81 2669
rect 47 2567 81 2601
rect 47 2499 81 2533
rect 47 2431 81 2465
rect 47 2363 81 2397
rect 47 2295 81 2329
rect 47 2227 81 2261
rect 47 2159 81 2193
rect 47 2091 81 2125
rect 47 2023 81 2057
rect 47 1955 81 1989
rect 47 1887 81 1921
rect 47 1819 81 1853
rect 47 1751 81 1785
rect 47 1683 81 1717
rect 47 1615 81 1649
rect 47 1547 81 1581
rect 47 1479 81 1513
rect 47 1411 81 1445
rect 47 1343 81 1377
rect 47 1275 81 1309
rect 47 1207 81 1241
rect 47 1139 81 1173
rect 47 1071 81 1105
rect 47 1003 81 1037
rect 47 935 81 969
rect 47 867 81 901
rect 47 799 81 833
rect 47 731 81 765
rect 47 663 81 697
rect 47 595 81 629
rect 47 527 81 561
rect 47 459 81 493
rect 47 391 81 425
rect 47 323 81 357
rect 47 255 81 289
rect 47 187 81 221
rect 47 119 81 153
rect 47 51 81 85
rect 47 -17 81 17
rect 47 -85 81 -51
rect 47 -153 81 -119
rect 47 -221 81 -187
rect 47 -289 81 -255
rect 47 -357 81 -323
rect 47 -425 81 -391
rect 47 -493 81 -459
rect 47 -561 81 -527
rect 47 -629 81 -595
rect 47 -697 81 -663
rect 47 -765 81 -731
rect 47 -833 81 -799
rect 47 -901 81 -867
rect 47 -969 81 -935
rect 47 -1037 81 -1003
rect 47 -1105 81 -1071
rect 47 -1173 81 -1139
rect 47 -1241 81 -1207
rect 47 -1309 81 -1275
rect 47 -1377 81 -1343
rect 47 -1445 81 -1411
rect 47 -1513 81 -1479
rect 47 -1581 81 -1547
rect 47 -1649 81 -1615
rect 47 -1717 81 -1683
rect 47 -1785 81 -1751
rect 47 -1853 81 -1819
rect 47 -1921 81 -1887
rect 47 -1989 81 -1955
rect 47 -2057 81 -2023
rect 47 -2125 81 -2091
rect 47 -2193 81 -2159
rect 47 -2261 81 -2227
rect 47 -2329 81 -2295
rect 47 -2397 81 -2363
rect 47 -2465 81 -2431
rect 47 -2533 81 -2499
rect 47 -2601 81 -2567
rect 47 -2669 81 -2635
rect 47 -2737 81 -2703
rect 47 -2805 81 -2771
rect 47 -2873 81 -2839
rect 47 -2941 81 -2907
rect 47 -3009 81 -2975
rect 47 -3077 81 -3043
rect 47 -3145 81 -3111
rect 47 -3213 81 -3179
rect 47 -3281 81 -3247
rect 47 -3349 81 -3315
rect 47 -3417 81 -3383
rect 47 -3485 81 -3451
rect 47 -3553 81 -3519
rect 47 -3621 81 -3587
rect 47 -3689 81 -3655
rect 47 -3757 81 -3723
rect 47 -3825 81 -3791
rect 47 -3893 81 -3859
rect 47 -3961 81 -3927
rect 47 -4029 81 -3995
rect 47 -4097 81 -4063
rect 47 -4165 81 -4131
rect 47 -4233 81 -4199
rect 47 -4301 81 -4267
rect 47 -4369 81 -4335
rect 47 -4437 81 -4403
rect 47 -4505 81 -4471
rect 47 -4573 81 -4539
rect 47 -4641 81 -4607
rect 47 -4709 81 -4675
rect 47 -4777 81 -4743
rect 47 -4845 81 -4811
rect 47 -4913 81 -4879
rect 47 -4981 81 -4947
<< nsubdiff >>
rect -195 5149 -85 5183
rect -51 5149 -17 5183
rect 17 5149 51 5183
rect 85 5149 195 5183
rect -195 5083 -161 5149
rect -195 5015 -161 5049
rect 161 5083 195 5149
rect 161 5015 195 5049
rect -195 4947 -161 4981
rect -195 4879 -161 4913
rect -195 4811 -161 4845
rect -195 4743 -161 4777
rect -195 4675 -161 4709
rect -195 4607 -161 4641
rect -195 4539 -161 4573
rect -195 4471 -161 4505
rect -195 4403 -161 4437
rect -195 4335 -161 4369
rect -195 4267 -161 4301
rect -195 4199 -161 4233
rect -195 4131 -161 4165
rect -195 4063 -161 4097
rect -195 3995 -161 4029
rect -195 3927 -161 3961
rect -195 3859 -161 3893
rect -195 3791 -161 3825
rect -195 3723 -161 3757
rect -195 3655 -161 3689
rect -195 3587 -161 3621
rect -195 3519 -161 3553
rect -195 3451 -161 3485
rect -195 3383 -161 3417
rect -195 3315 -161 3349
rect -195 3247 -161 3281
rect -195 3179 -161 3213
rect -195 3111 -161 3145
rect -195 3043 -161 3077
rect -195 2975 -161 3009
rect -195 2907 -161 2941
rect -195 2839 -161 2873
rect -195 2771 -161 2805
rect -195 2703 -161 2737
rect -195 2635 -161 2669
rect -195 2567 -161 2601
rect -195 2499 -161 2533
rect -195 2431 -161 2465
rect -195 2363 -161 2397
rect -195 2295 -161 2329
rect -195 2227 -161 2261
rect -195 2159 -161 2193
rect -195 2091 -161 2125
rect -195 2023 -161 2057
rect -195 1955 -161 1989
rect -195 1887 -161 1921
rect -195 1819 -161 1853
rect -195 1751 -161 1785
rect -195 1683 -161 1717
rect -195 1615 -161 1649
rect -195 1547 -161 1581
rect -195 1479 -161 1513
rect -195 1411 -161 1445
rect -195 1343 -161 1377
rect -195 1275 -161 1309
rect -195 1207 -161 1241
rect -195 1139 -161 1173
rect -195 1071 -161 1105
rect -195 1003 -161 1037
rect -195 935 -161 969
rect -195 867 -161 901
rect -195 799 -161 833
rect -195 731 -161 765
rect -195 663 -161 697
rect -195 595 -161 629
rect -195 527 -161 561
rect -195 459 -161 493
rect -195 391 -161 425
rect -195 323 -161 357
rect -195 255 -161 289
rect -195 187 -161 221
rect -195 119 -161 153
rect -195 51 -161 85
rect -195 -17 -161 17
rect -195 -85 -161 -51
rect -195 -153 -161 -119
rect -195 -221 -161 -187
rect -195 -289 -161 -255
rect -195 -357 -161 -323
rect -195 -425 -161 -391
rect -195 -493 -161 -459
rect -195 -561 -161 -527
rect -195 -629 -161 -595
rect -195 -697 -161 -663
rect -195 -765 -161 -731
rect -195 -833 -161 -799
rect -195 -901 -161 -867
rect -195 -969 -161 -935
rect -195 -1037 -161 -1003
rect -195 -1105 -161 -1071
rect -195 -1173 -161 -1139
rect -195 -1241 -161 -1207
rect -195 -1309 -161 -1275
rect -195 -1377 -161 -1343
rect -195 -1445 -161 -1411
rect -195 -1513 -161 -1479
rect -195 -1581 -161 -1547
rect -195 -1649 -161 -1615
rect -195 -1717 -161 -1683
rect -195 -1785 -161 -1751
rect -195 -1853 -161 -1819
rect -195 -1921 -161 -1887
rect -195 -1989 -161 -1955
rect -195 -2057 -161 -2023
rect -195 -2125 -161 -2091
rect -195 -2193 -161 -2159
rect -195 -2261 -161 -2227
rect -195 -2329 -161 -2295
rect -195 -2397 -161 -2363
rect -195 -2465 -161 -2431
rect -195 -2533 -161 -2499
rect -195 -2601 -161 -2567
rect -195 -2669 -161 -2635
rect -195 -2737 -161 -2703
rect -195 -2805 -161 -2771
rect -195 -2873 -161 -2839
rect -195 -2941 -161 -2907
rect -195 -3009 -161 -2975
rect -195 -3077 -161 -3043
rect -195 -3145 -161 -3111
rect -195 -3213 -161 -3179
rect -195 -3281 -161 -3247
rect -195 -3349 -161 -3315
rect -195 -3417 -161 -3383
rect -195 -3485 -161 -3451
rect -195 -3553 -161 -3519
rect -195 -3621 -161 -3587
rect -195 -3689 -161 -3655
rect -195 -3757 -161 -3723
rect -195 -3825 -161 -3791
rect -195 -3893 -161 -3859
rect -195 -3961 -161 -3927
rect -195 -4029 -161 -3995
rect -195 -4097 -161 -4063
rect -195 -4165 -161 -4131
rect -195 -4233 -161 -4199
rect -195 -4301 -161 -4267
rect -195 -4369 -161 -4335
rect -195 -4437 -161 -4403
rect -195 -4505 -161 -4471
rect -195 -4573 -161 -4539
rect -195 -4641 -161 -4607
rect -195 -4709 -161 -4675
rect -195 -4777 -161 -4743
rect -195 -4845 -161 -4811
rect -195 -4913 -161 -4879
rect -195 -4981 -161 -4947
rect 161 4947 195 4981
rect 161 4879 195 4913
rect 161 4811 195 4845
rect 161 4743 195 4777
rect 161 4675 195 4709
rect 161 4607 195 4641
rect 161 4539 195 4573
rect 161 4471 195 4505
rect 161 4403 195 4437
rect 161 4335 195 4369
rect 161 4267 195 4301
rect 161 4199 195 4233
rect 161 4131 195 4165
rect 161 4063 195 4097
rect 161 3995 195 4029
rect 161 3927 195 3961
rect 161 3859 195 3893
rect 161 3791 195 3825
rect 161 3723 195 3757
rect 161 3655 195 3689
rect 161 3587 195 3621
rect 161 3519 195 3553
rect 161 3451 195 3485
rect 161 3383 195 3417
rect 161 3315 195 3349
rect 161 3247 195 3281
rect 161 3179 195 3213
rect 161 3111 195 3145
rect 161 3043 195 3077
rect 161 2975 195 3009
rect 161 2907 195 2941
rect 161 2839 195 2873
rect 161 2771 195 2805
rect 161 2703 195 2737
rect 161 2635 195 2669
rect 161 2567 195 2601
rect 161 2499 195 2533
rect 161 2431 195 2465
rect 161 2363 195 2397
rect 161 2295 195 2329
rect 161 2227 195 2261
rect 161 2159 195 2193
rect 161 2091 195 2125
rect 161 2023 195 2057
rect 161 1955 195 1989
rect 161 1887 195 1921
rect 161 1819 195 1853
rect 161 1751 195 1785
rect 161 1683 195 1717
rect 161 1615 195 1649
rect 161 1547 195 1581
rect 161 1479 195 1513
rect 161 1411 195 1445
rect 161 1343 195 1377
rect 161 1275 195 1309
rect 161 1207 195 1241
rect 161 1139 195 1173
rect 161 1071 195 1105
rect 161 1003 195 1037
rect 161 935 195 969
rect 161 867 195 901
rect 161 799 195 833
rect 161 731 195 765
rect 161 663 195 697
rect 161 595 195 629
rect 161 527 195 561
rect 161 459 195 493
rect 161 391 195 425
rect 161 323 195 357
rect 161 255 195 289
rect 161 187 195 221
rect 161 119 195 153
rect 161 51 195 85
rect 161 -17 195 17
rect 161 -85 195 -51
rect 161 -153 195 -119
rect 161 -221 195 -187
rect 161 -289 195 -255
rect 161 -357 195 -323
rect 161 -425 195 -391
rect 161 -493 195 -459
rect 161 -561 195 -527
rect 161 -629 195 -595
rect 161 -697 195 -663
rect 161 -765 195 -731
rect 161 -833 195 -799
rect 161 -901 195 -867
rect 161 -969 195 -935
rect 161 -1037 195 -1003
rect 161 -1105 195 -1071
rect 161 -1173 195 -1139
rect 161 -1241 195 -1207
rect 161 -1309 195 -1275
rect 161 -1377 195 -1343
rect 161 -1445 195 -1411
rect 161 -1513 195 -1479
rect 161 -1581 195 -1547
rect 161 -1649 195 -1615
rect 161 -1717 195 -1683
rect 161 -1785 195 -1751
rect 161 -1853 195 -1819
rect 161 -1921 195 -1887
rect 161 -1989 195 -1955
rect 161 -2057 195 -2023
rect 161 -2125 195 -2091
rect 161 -2193 195 -2159
rect 161 -2261 195 -2227
rect 161 -2329 195 -2295
rect 161 -2397 195 -2363
rect 161 -2465 195 -2431
rect 161 -2533 195 -2499
rect 161 -2601 195 -2567
rect 161 -2669 195 -2635
rect 161 -2737 195 -2703
rect 161 -2805 195 -2771
rect 161 -2873 195 -2839
rect 161 -2941 195 -2907
rect 161 -3009 195 -2975
rect 161 -3077 195 -3043
rect 161 -3145 195 -3111
rect 161 -3213 195 -3179
rect 161 -3281 195 -3247
rect 161 -3349 195 -3315
rect 161 -3417 195 -3383
rect 161 -3485 195 -3451
rect 161 -3553 195 -3519
rect 161 -3621 195 -3587
rect 161 -3689 195 -3655
rect 161 -3757 195 -3723
rect 161 -3825 195 -3791
rect 161 -3893 195 -3859
rect 161 -3961 195 -3927
rect 161 -4029 195 -3995
rect 161 -4097 195 -4063
rect 161 -4165 195 -4131
rect 161 -4233 195 -4199
rect 161 -4301 195 -4267
rect 161 -4369 195 -4335
rect 161 -4437 195 -4403
rect 161 -4505 195 -4471
rect 161 -4573 195 -4539
rect 161 -4641 195 -4607
rect 161 -4709 195 -4675
rect 161 -4777 195 -4743
rect 161 -4845 195 -4811
rect 161 -4913 195 -4879
rect 161 -4981 195 -4947
rect -195 -5049 -161 -5015
rect -195 -5149 -161 -5083
rect 161 -5049 195 -5015
rect 161 -5149 195 -5083
rect -195 -5183 -85 -5149
rect -51 -5183 -17 -5149
rect 17 -5183 51 -5149
rect 85 -5183 195 -5149
<< nsubdiffcont >>
rect -85 5149 -51 5183
rect -17 5149 17 5183
rect 51 5149 85 5183
rect -195 5049 -161 5083
rect -195 4981 -161 5015
rect 161 5049 195 5083
rect -195 4913 -161 4947
rect -195 4845 -161 4879
rect -195 4777 -161 4811
rect -195 4709 -161 4743
rect -195 4641 -161 4675
rect -195 4573 -161 4607
rect -195 4505 -161 4539
rect -195 4437 -161 4471
rect -195 4369 -161 4403
rect -195 4301 -161 4335
rect -195 4233 -161 4267
rect -195 4165 -161 4199
rect -195 4097 -161 4131
rect -195 4029 -161 4063
rect -195 3961 -161 3995
rect -195 3893 -161 3927
rect -195 3825 -161 3859
rect -195 3757 -161 3791
rect -195 3689 -161 3723
rect -195 3621 -161 3655
rect -195 3553 -161 3587
rect -195 3485 -161 3519
rect -195 3417 -161 3451
rect -195 3349 -161 3383
rect -195 3281 -161 3315
rect -195 3213 -161 3247
rect -195 3145 -161 3179
rect -195 3077 -161 3111
rect -195 3009 -161 3043
rect -195 2941 -161 2975
rect -195 2873 -161 2907
rect -195 2805 -161 2839
rect -195 2737 -161 2771
rect -195 2669 -161 2703
rect -195 2601 -161 2635
rect -195 2533 -161 2567
rect -195 2465 -161 2499
rect -195 2397 -161 2431
rect -195 2329 -161 2363
rect -195 2261 -161 2295
rect -195 2193 -161 2227
rect -195 2125 -161 2159
rect -195 2057 -161 2091
rect -195 1989 -161 2023
rect -195 1921 -161 1955
rect -195 1853 -161 1887
rect -195 1785 -161 1819
rect -195 1717 -161 1751
rect -195 1649 -161 1683
rect -195 1581 -161 1615
rect -195 1513 -161 1547
rect -195 1445 -161 1479
rect -195 1377 -161 1411
rect -195 1309 -161 1343
rect -195 1241 -161 1275
rect -195 1173 -161 1207
rect -195 1105 -161 1139
rect -195 1037 -161 1071
rect -195 969 -161 1003
rect -195 901 -161 935
rect -195 833 -161 867
rect -195 765 -161 799
rect -195 697 -161 731
rect -195 629 -161 663
rect -195 561 -161 595
rect -195 493 -161 527
rect -195 425 -161 459
rect -195 357 -161 391
rect -195 289 -161 323
rect -195 221 -161 255
rect -195 153 -161 187
rect -195 85 -161 119
rect -195 17 -161 51
rect -195 -51 -161 -17
rect -195 -119 -161 -85
rect -195 -187 -161 -153
rect -195 -255 -161 -221
rect -195 -323 -161 -289
rect -195 -391 -161 -357
rect -195 -459 -161 -425
rect -195 -527 -161 -493
rect -195 -595 -161 -561
rect -195 -663 -161 -629
rect -195 -731 -161 -697
rect -195 -799 -161 -765
rect -195 -867 -161 -833
rect -195 -935 -161 -901
rect -195 -1003 -161 -969
rect -195 -1071 -161 -1037
rect -195 -1139 -161 -1105
rect -195 -1207 -161 -1173
rect -195 -1275 -161 -1241
rect -195 -1343 -161 -1309
rect -195 -1411 -161 -1377
rect -195 -1479 -161 -1445
rect -195 -1547 -161 -1513
rect -195 -1615 -161 -1581
rect -195 -1683 -161 -1649
rect -195 -1751 -161 -1717
rect -195 -1819 -161 -1785
rect -195 -1887 -161 -1853
rect -195 -1955 -161 -1921
rect -195 -2023 -161 -1989
rect -195 -2091 -161 -2057
rect -195 -2159 -161 -2125
rect -195 -2227 -161 -2193
rect -195 -2295 -161 -2261
rect -195 -2363 -161 -2329
rect -195 -2431 -161 -2397
rect -195 -2499 -161 -2465
rect -195 -2567 -161 -2533
rect -195 -2635 -161 -2601
rect -195 -2703 -161 -2669
rect -195 -2771 -161 -2737
rect -195 -2839 -161 -2805
rect -195 -2907 -161 -2873
rect -195 -2975 -161 -2941
rect -195 -3043 -161 -3009
rect -195 -3111 -161 -3077
rect -195 -3179 -161 -3145
rect -195 -3247 -161 -3213
rect -195 -3315 -161 -3281
rect -195 -3383 -161 -3349
rect -195 -3451 -161 -3417
rect -195 -3519 -161 -3485
rect -195 -3587 -161 -3553
rect -195 -3655 -161 -3621
rect -195 -3723 -161 -3689
rect -195 -3791 -161 -3757
rect -195 -3859 -161 -3825
rect -195 -3927 -161 -3893
rect -195 -3995 -161 -3961
rect -195 -4063 -161 -4029
rect -195 -4131 -161 -4097
rect -195 -4199 -161 -4165
rect -195 -4267 -161 -4233
rect -195 -4335 -161 -4301
rect -195 -4403 -161 -4369
rect -195 -4471 -161 -4437
rect -195 -4539 -161 -4505
rect -195 -4607 -161 -4573
rect -195 -4675 -161 -4641
rect -195 -4743 -161 -4709
rect -195 -4811 -161 -4777
rect -195 -4879 -161 -4845
rect -195 -4947 -161 -4913
rect -195 -5015 -161 -4981
rect 161 4981 195 5015
rect 161 4913 195 4947
rect 161 4845 195 4879
rect 161 4777 195 4811
rect 161 4709 195 4743
rect 161 4641 195 4675
rect 161 4573 195 4607
rect 161 4505 195 4539
rect 161 4437 195 4471
rect 161 4369 195 4403
rect 161 4301 195 4335
rect 161 4233 195 4267
rect 161 4165 195 4199
rect 161 4097 195 4131
rect 161 4029 195 4063
rect 161 3961 195 3995
rect 161 3893 195 3927
rect 161 3825 195 3859
rect 161 3757 195 3791
rect 161 3689 195 3723
rect 161 3621 195 3655
rect 161 3553 195 3587
rect 161 3485 195 3519
rect 161 3417 195 3451
rect 161 3349 195 3383
rect 161 3281 195 3315
rect 161 3213 195 3247
rect 161 3145 195 3179
rect 161 3077 195 3111
rect 161 3009 195 3043
rect 161 2941 195 2975
rect 161 2873 195 2907
rect 161 2805 195 2839
rect 161 2737 195 2771
rect 161 2669 195 2703
rect 161 2601 195 2635
rect 161 2533 195 2567
rect 161 2465 195 2499
rect 161 2397 195 2431
rect 161 2329 195 2363
rect 161 2261 195 2295
rect 161 2193 195 2227
rect 161 2125 195 2159
rect 161 2057 195 2091
rect 161 1989 195 2023
rect 161 1921 195 1955
rect 161 1853 195 1887
rect 161 1785 195 1819
rect 161 1717 195 1751
rect 161 1649 195 1683
rect 161 1581 195 1615
rect 161 1513 195 1547
rect 161 1445 195 1479
rect 161 1377 195 1411
rect 161 1309 195 1343
rect 161 1241 195 1275
rect 161 1173 195 1207
rect 161 1105 195 1139
rect 161 1037 195 1071
rect 161 969 195 1003
rect 161 901 195 935
rect 161 833 195 867
rect 161 765 195 799
rect 161 697 195 731
rect 161 629 195 663
rect 161 561 195 595
rect 161 493 195 527
rect 161 425 195 459
rect 161 357 195 391
rect 161 289 195 323
rect 161 221 195 255
rect 161 153 195 187
rect 161 85 195 119
rect 161 17 195 51
rect 161 -51 195 -17
rect 161 -119 195 -85
rect 161 -187 195 -153
rect 161 -255 195 -221
rect 161 -323 195 -289
rect 161 -391 195 -357
rect 161 -459 195 -425
rect 161 -527 195 -493
rect 161 -595 195 -561
rect 161 -663 195 -629
rect 161 -731 195 -697
rect 161 -799 195 -765
rect 161 -867 195 -833
rect 161 -935 195 -901
rect 161 -1003 195 -969
rect 161 -1071 195 -1037
rect 161 -1139 195 -1105
rect 161 -1207 195 -1173
rect 161 -1275 195 -1241
rect 161 -1343 195 -1309
rect 161 -1411 195 -1377
rect 161 -1479 195 -1445
rect 161 -1547 195 -1513
rect 161 -1615 195 -1581
rect 161 -1683 195 -1649
rect 161 -1751 195 -1717
rect 161 -1819 195 -1785
rect 161 -1887 195 -1853
rect 161 -1955 195 -1921
rect 161 -2023 195 -1989
rect 161 -2091 195 -2057
rect 161 -2159 195 -2125
rect 161 -2227 195 -2193
rect 161 -2295 195 -2261
rect 161 -2363 195 -2329
rect 161 -2431 195 -2397
rect 161 -2499 195 -2465
rect 161 -2567 195 -2533
rect 161 -2635 195 -2601
rect 161 -2703 195 -2669
rect 161 -2771 195 -2737
rect 161 -2839 195 -2805
rect 161 -2907 195 -2873
rect 161 -2975 195 -2941
rect 161 -3043 195 -3009
rect 161 -3111 195 -3077
rect 161 -3179 195 -3145
rect 161 -3247 195 -3213
rect 161 -3315 195 -3281
rect 161 -3383 195 -3349
rect 161 -3451 195 -3417
rect 161 -3519 195 -3485
rect 161 -3587 195 -3553
rect 161 -3655 195 -3621
rect 161 -3723 195 -3689
rect 161 -3791 195 -3757
rect 161 -3859 195 -3825
rect 161 -3927 195 -3893
rect 161 -3995 195 -3961
rect 161 -4063 195 -4029
rect 161 -4131 195 -4097
rect 161 -4199 195 -4165
rect 161 -4267 195 -4233
rect 161 -4335 195 -4301
rect 161 -4403 195 -4369
rect 161 -4471 195 -4437
rect 161 -4539 195 -4505
rect 161 -4607 195 -4573
rect 161 -4675 195 -4641
rect 161 -4743 195 -4709
rect 161 -4811 195 -4777
rect 161 -4879 195 -4845
rect 161 -4947 195 -4913
rect -195 -5083 -161 -5049
rect 161 -5015 195 -4981
rect 161 -5083 195 -5049
rect -85 -5183 -51 -5149
rect -17 -5183 17 -5149
rect 51 -5183 85 -5149
<< poly >>
rect -35 5081 35 5097
rect -35 5047 -17 5081
rect 17 5047 35 5081
rect -35 5000 35 5047
rect -35 -5047 35 -5000
rect -35 -5081 -17 -5047
rect 17 -5081 35 -5047
rect -35 -5097 35 -5081
<< polycont >>
rect -17 5047 17 5081
rect -17 -5081 17 -5047
<< locali >>
rect -195 5149 -85 5183
rect -51 5149 -17 5183
rect 17 5149 51 5183
rect 85 5149 195 5183
rect -195 5083 -161 5149
rect 161 5083 195 5149
rect -195 5015 -161 5049
rect -35 5047 -17 5081
rect 17 5047 35 5081
rect 161 5015 195 5049
rect -195 4947 -161 4981
rect -195 4879 -161 4913
rect -195 4811 -161 4845
rect -195 4743 -161 4777
rect -195 4675 -161 4709
rect -195 4607 -161 4641
rect -195 4539 -161 4573
rect -195 4471 -161 4505
rect -195 4403 -161 4437
rect -195 4335 -161 4369
rect -195 4267 -161 4301
rect -195 4199 -161 4233
rect -195 4131 -161 4165
rect -195 4063 -161 4097
rect -195 3995 -161 4029
rect -195 3927 -161 3961
rect -195 3859 -161 3893
rect -195 3791 -161 3825
rect -195 3723 -161 3757
rect -195 3655 -161 3689
rect -195 3587 -161 3621
rect -195 3519 -161 3553
rect -195 3451 -161 3485
rect -195 3383 -161 3417
rect -195 3315 -161 3349
rect -195 3247 -161 3281
rect -195 3179 -161 3213
rect -195 3111 -161 3145
rect -195 3043 -161 3077
rect -195 2975 -161 3009
rect -195 2907 -161 2941
rect -195 2839 -161 2873
rect -195 2771 -161 2805
rect -195 2703 -161 2737
rect -195 2635 -161 2669
rect -195 2567 -161 2601
rect -195 2499 -161 2533
rect -195 2431 -161 2465
rect -195 2363 -161 2397
rect -195 2295 -161 2329
rect -195 2227 -161 2261
rect -195 2159 -161 2193
rect -195 2091 -161 2125
rect -195 2023 -161 2057
rect -195 1955 -161 1989
rect -195 1887 -161 1921
rect -195 1819 -161 1853
rect -195 1751 -161 1785
rect -195 1683 -161 1717
rect -195 1615 -161 1649
rect -195 1547 -161 1581
rect -195 1479 -161 1513
rect -195 1411 -161 1445
rect -195 1343 -161 1377
rect -195 1275 -161 1309
rect -195 1207 -161 1241
rect -195 1139 -161 1173
rect -195 1071 -161 1105
rect -195 1003 -161 1037
rect -195 935 -161 969
rect -195 867 -161 901
rect -195 799 -161 833
rect -195 731 -161 765
rect -195 663 -161 697
rect -195 595 -161 629
rect -195 527 -161 561
rect -195 459 -161 493
rect -195 391 -161 425
rect -195 323 -161 357
rect -195 255 -161 289
rect -195 187 -161 221
rect -195 119 -161 153
rect -195 51 -161 85
rect -195 -17 -161 17
rect -195 -85 -161 -51
rect -195 -153 -161 -119
rect -195 -221 -161 -187
rect -195 -289 -161 -255
rect -195 -357 -161 -323
rect -195 -425 -161 -391
rect -195 -493 -161 -459
rect -195 -561 -161 -527
rect -195 -629 -161 -595
rect -195 -697 -161 -663
rect -195 -765 -161 -731
rect -195 -833 -161 -799
rect -195 -901 -161 -867
rect -195 -969 -161 -935
rect -195 -1037 -161 -1003
rect -195 -1105 -161 -1071
rect -195 -1173 -161 -1139
rect -195 -1241 -161 -1207
rect -195 -1309 -161 -1275
rect -195 -1377 -161 -1343
rect -195 -1445 -161 -1411
rect -195 -1513 -161 -1479
rect -195 -1581 -161 -1547
rect -195 -1649 -161 -1615
rect -195 -1717 -161 -1683
rect -195 -1785 -161 -1751
rect -195 -1853 -161 -1819
rect -195 -1921 -161 -1887
rect -195 -1989 -161 -1955
rect -195 -2057 -161 -2023
rect -195 -2125 -161 -2091
rect -195 -2193 -161 -2159
rect -195 -2261 -161 -2227
rect -195 -2329 -161 -2295
rect -195 -2397 -161 -2363
rect -195 -2465 -161 -2431
rect -195 -2533 -161 -2499
rect -195 -2601 -161 -2567
rect -195 -2669 -161 -2635
rect -195 -2737 -161 -2703
rect -195 -2805 -161 -2771
rect -195 -2873 -161 -2839
rect -195 -2941 -161 -2907
rect -195 -3009 -161 -2975
rect -195 -3077 -161 -3043
rect -195 -3145 -161 -3111
rect -195 -3213 -161 -3179
rect -195 -3281 -161 -3247
rect -195 -3349 -161 -3315
rect -195 -3417 -161 -3383
rect -195 -3485 -161 -3451
rect -195 -3553 -161 -3519
rect -195 -3621 -161 -3587
rect -195 -3689 -161 -3655
rect -195 -3757 -161 -3723
rect -195 -3825 -161 -3791
rect -195 -3893 -161 -3859
rect -195 -3961 -161 -3927
rect -195 -4029 -161 -3995
rect -195 -4097 -161 -4063
rect -195 -4165 -161 -4131
rect -195 -4233 -161 -4199
rect -195 -4301 -161 -4267
rect -195 -4369 -161 -4335
rect -195 -4437 -161 -4403
rect -195 -4505 -161 -4471
rect -195 -4573 -161 -4539
rect -195 -4641 -161 -4607
rect -195 -4709 -161 -4675
rect -195 -4777 -161 -4743
rect -195 -4845 -161 -4811
rect -195 -4913 -161 -4879
rect -195 -4981 -161 -4947
rect -81 4985 -47 5004
rect -81 4913 -47 4947
rect -81 4845 -47 4879
rect -81 4777 -47 4807
rect -81 4709 -47 4735
rect -81 4641 -47 4663
rect -81 4573 -47 4591
rect -81 4505 -47 4519
rect -81 4437 -47 4447
rect -81 4369 -47 4375
rect -81 4301 -47 4303
rect -81 4265 -47 4267
rect -81 4193 -47 4199
rect -81 4121 -47 4131
rect -81 4049 -47 4063
rect -81 3977 -47 3995
rect -81 3905 -47 3927
rect -81 3833 -47 3859
rect -81 3761 -47 3791
rect -81 3689 -47 3723
rect -81 3621 -47 3655
rect -81 3553 -47 3583
rect -81 3485 -47 3511
rect -81 3417 -47 3439
rect -81 3349 -47 3367
rect -81 3281 -47 3295
rect -81 3213 -47 3223
rect -81 3145 -47 3151
rect -81 3077 -47 3079
rect -81 3041 -47 3043
rect -81 2969 -47 2975
rect -81 2897 -47 2907
rect -81 2825 -47 2839
rect -81 2753 -47 2771
rect -81 2681 -47 2703
rect -81 2609 -47 2635
rect -81 2537 -47 2567
rect -81 2465 -47 2499
rect -81 2397 -47 2431
rect -81 2329 -47 2359
rect -81 2261 -47 2287
rect -81 2193 -47 2215
rect -81 2125 -47 2143
rect -81 2057 -47 2071
rect -81 1989 -47 1999
rect -81 1921 -47 1927
rect -81 1853 -47 1855
rect -81 1817 -47 1819
rect -81 1745 -47 1751
rect -81 1673 -47 1683
rect -81 1601 -47 1615
rect -81 1529 -47 1547
rect -81 1457 -47 1479
rect -81 1385 -47 1411
rect -81 1313 -47 1343
rect -81 1241 -47 1275
rect -81 1173 -47 1207
rect -81 1105 -47 1135
rect -81 1037 -47 1063
rect -81 969 -47 991
rect -81 901 -47 919
rect -81 833 -47 847
rect -81 765 -47 775
rect -81 697 -47 703
rect -81 629 -47 631
rect -81 593 -47 595
rect -81 521 -47 527
rect -81 449 -47 459
rect -81 377 -47 391
rect -81 305 -47 323
rect -81 233 -47 255
rect -81 161 -47 187
rect -81 89 -47 119
rect -81 17 -47 51
rect -81 -51 -47 -17
rect -81 -119 -47 -89
rect -81 -187 -47 -161
rect -81 -255 -47 -233
rect -81 -323 -47 -305
rect -81 -391 -47 -377
rect -81 -459 -47 -449
rect -81 -527 -47 -521
rect -81 -595 -47 -593
rect -81 -631 -47 -629
rect -81 -703 -47 -697
rect -81 -775 -47 -765
rect -81 -847 -47 -833
rect -81 -919 -47 -901
rect -81 -991 -47 -969
rect -81 -1063 -47 -1037
rect -81 -1135 -47 -1105
rect -81 -1207 -47 -1173
rect -81 -1275 -47 -1241
rect -81 -1343 -47 -1313
rect -81 -1411 -47 -1385
rect -81 -1479 -47 -1457
rect -81 -1547 -47 -1529
rect -81 -1615 -47 -1601
rect -81 -1683 -47 -1673
rect -81 -1751 -47 -1745
rect -81 -1819 -47 -1817
rect -81 -1855 -47 -1853
rect -81 -1927 -47 -1921
rect -81 -1999 -47 -1989
rect -81 -2071 -47 -2057
rect -81 -2143 -47 -2125
rect -81 -2215 -47 -2193
rect -81 -2287 -47 -2261
rect -81 -2359 -47 -2329
rect -81 -2431 -47 -2397
rect -81 -2499 -47 -2465
rect -81 -2567 -47 -2537
rect -81 -2635 -47 -2609
rect -81 -2703 -47 -2681
rect -81 -2771 -47 -2753
rect -81 -2839 -47 -2825
rect -81 -2907 -47 -2897
rect -81 -2975 -47 -2969
rect -81 -3043 -47 -3041
rect -81 -3079 -47 -3077
rect -81 -3151 -47 -3145
rect -81 -3223 -47 -3213
rect -81 -3295 -47 -3281
rect -81 -3367 -47 -3349
rect -81 -3439 -47 -3417
rect -81 -3511 -47 -3485
rect -81 -3583 -47 -3553
rect -81 -3655 -47 -3621
rect -81 -3723 -47 -3689
rect -81 -3791 -47 -3761
rect -81 -3859 -47 -3833
rect -81 -3927 -47 -3905
rect -81 -3995 -47 -3977
rect -81 -4063 -47 -4049
rect -81 -4131 -47 -4121
rect -81 -4199 -47 -4193
rect -81 -4267 -47 -4265
rect -81 -4303 -47 -4301
rect -81 -4375 -47 -4369
rect -81 -4447 -47 -4437
rect -81 -4519 -47 -4505
rect -81 -4591 -47 -4573
rect -81 -4663 -47 -4641
rect -81 -4735 -47 -4709
rect -81 -4807 -47 -4777
rect -81 -4879 -47 -4845
rect -81 -4947 -47 -4913
rect -81 -5004 -47 -4985
rect 47 4985 81 5004
rect 47 4913 81 4947
rect 47 4845 81 4879
rect 47 4777 81 4807
rect 47 4709 81 4735
rect 47 4641 81 4663
rect 47 4573 81 4591
rect 47 4505 81 4519
rect 47 4437 81 4447
rect 47 4369 81 4375
rect 47 4301 81 4303
rect 47 4265 81 4267
rect 47 4193 81 4199
rect 47 4121 81 4131
rect 47 4049 81 4063
rect 47 3977 81 3995
rect 47 3905 81 3927
rect 47 3833 81 3859
rect 47 3761 81 3791
rect 47 3689 81 3723
rect 47 3621 81 3655
rect 47 3553 81 3583
rect 47 3485 81 3511
rect 47 3417 81 3439
rect 47 3349 81 3367
rect 47 3281 81 3295
rect 47 3213 81 3223
rect 47 3145 81 3151
rect 47 3077 81 3079
rect 47 3041 81 3043
rect 47 2969 81 2975
rect 47 2897 81 2907
rect 47 2825 81 2839
rect 47 2753 81 2771
rect 47 2681 81 2703
rect 47 2609 81 2635
rect 47 2537 81 2567
rect 47 2465 81 2499
rect 47 2397 81 2431
rect 47 2329 81 2359
rect 47 2261 81 2287
rect 47 2193 81 2215
rect 47 2125 81 2143
rect 47 2057 81 2071
rect 47 1989 81 1999
rect 47 1921 81 1927
rect 47 1853 81 1855
rect 47 1817 81 1819
rect 47 1745 81 1751
rect 47 1673 81 1683
rect 47 1601 81 1615
rect 47 1529 81 1547
rect 47 1457 81 1479
rect 47 1385 81 1411
rect 47 1313 81 1343
rect 47 1241 81 1275
rect 47 1173 81 1207
rect 47 1105 81 1135
rect 47 1037 81 1063
rect 47 969 81 991
rect 47 901 81 919
rect 47 833 81 847
rect 47 765 81 775
rect 47 697 81 703
rect 47 629 81 631
rect 47 593 81 595
rect 47 521 81 527
rect 47 449 81 459
rect 47 377 81 391
rect 47 305 81 323
rect 47 233 81 255
rect 47 161 81 187
rect 47 89 81 119
rect 47 17 81 51
rect 47 -51 81 -17
rect 47 -119 81 -89
rect 47 -187 81 -161
rect 47 -255 81 -233
rect 47 -323 81 -305
rect 47 -391 81 -377
rect 47 -459 81 -449
rect 47 -527 81 -521
rect 47 -595 81 -593
rect 47 -631 81 -629
rect 47 -703 81 -697
rect 47 -775 81 -765
rect 47 -847 81 -833
rect 47 -919 81 -901
rect 47 -991 81 -969
rect 47 -1063 81 -1037
rect 47 -1135 81 -1105
rect 47 -1207 81 -1173
rect 47 -1275 81 -1241
rect 47 -1343 81 -1313
rect 47 -1411 81 -1385
rect 47 -1479 81 -1457
rect 47 -1547 81 -1529
rect 47 -1615 81 -1601
rect 47 -1683 81 -1673
rect 47 -1751 81 -1745
rect 47 -1819 81 -1817
rect 47 -1855 81 -1853
rect 47 -1927 81 -1921
rect 47 -1999 81 -1989
rect 47 -2071 81 -2057
rect 47 -2143 81 -2125
rect 47 -2215 81 -2193
rect 47 -2287 81 -2261
rect 47 -2359 81 -2329
rect 47 -2431 81 -2397
rect 47 -2499 81 -2465
rect 47 -2567 81 -2537
rect 47 -2635 81 -2609
rect 47 -2703 81 -2681
rect 47 -2771 81 -2753
rect 47 -2839 81 -2825
rect 47 -2907 81 -2897
rect 47 -2975 81 -2969
rect 47 -3043 81 -3041
rect 47 -3079 81 -3077
rect 47 -3151 81 -3145
rect 47 -3223 81 -3213
rect 47 -3295 81 -3281
rect 47 -3367 81 -3349
rect 47 -3439 81 -3417
rect 47 -3511 81 -3485
rect 47 -3583 81 -3553
rect 47 -3655 81 -3621
rect 47 -3723 81 -3689
rect 47 -3791 81 -3761
rect 47 -3859 81 -3833
rect 47 -3927 81 -3905
rect 47 -3995 81 -3977
rect 47 -4063 81 -4049
rect 47 -4131 81 -4121
rect 47 -4199 81 -4193
rect 47 -4267 81 -4265
rect 47 -4303 81 -4301
rect 47 -4375 81 -4369
rect 47 -4447 81 -4437
rect 47 -4519 81 -4505
rect 47 -4591 81 -4573
rect 47 -4663 81 -4641
rect 47 -4735 81 -4709
rect 47 -4807 81 -4777
rect 47 -4879 81 -4845
rect 47 -4947 81 -4913
rect 47 -5004 81 -4985
rect 161 4947 195 4981
rect 161 4879 195 4913
rect 161 4811 195 4845
rect 161 4743 195 4777
rect 161 4675 195 4709
rect 161 4607 195 4641
rect 161 4539 195 4573
rect 161 4471 195 4505
rect 161 4403 195 4437
rect 161 4335 195 4369
rect 161 4267 195 4301
rect 161 4199 195 4233
rect 161 4131 195 4165
rect 161 4063 195 4097
rect 161 3995 195 4029
rect 161 3927 195 3961
rect 161 3859 195 3893
rect 161 3791 195 3825
rect 161 3723 195 3757
rect 161 3655 195 3689
rect 161 3587 195 3621
rect 161 3519 195 3553
rect 161 3451 195 3485
rect 161 3383 195 3417
rect 161 3315 195 3349
rect 161 3247 195 3281
rect 161 3179 195 3213
rect 161 3111 195 3145
rect 161 3043 195 3077
rect 161 2975 195 3009
rect 161 2907 195 2941
rect 161 2839 195 2873
rect 161 2771 195 2805
rect 161 2703 195 2737
rect 161 2635 195 2669
rect 161 2567 195 2601
rect 161 2499 195 2533
rect 161 2431 195 2465
rect 161 2363 195 2397
rect 161 2295 195 2329
rect 161 2227 195 2261
rect 161 2159 195 2193
rect 161 2091 195 2125
rect 161 2023 195 2057
rect 161 1955 195 1989
rect 161 1887 195 1921
rect 161 1819 195 1853
rect 161 1751 195 1785
rect 161 1683 195 1717
rect 161 1615 195 1649
rect 161 1547 195 1581
rect 161 1479 195 1513
rect 161 1411 195 1445
rect 161 1343 195 1377
rect 161 1275 195 1309
rect 161 1207 195 1241
rect 161 1139 195 1173
rect 161 1071 195 1105
rect 161 1003 195 1037
rect 161 935 195 969
rect 161 867 195 901
rect 161 799 195 833
rect 161 731 195 765
rect 161 663 195 697
rect 161 595 195 629
rect 161 527 195 561
rect 161 459 195 493
rect 161 391 195 425
rect 161 323 195 357
rect 161 255 195 289
rect 161 187 195 221
rect 161 119 195 153
rect 161 51 195 85
rect 161 -17 195 17
rect 161 -85 195 -51
rect 161 -153 195 -119
rect 161 -221 195 -187
rect 161 -289 195 -255
rect 161 -357 195 -323
rect 161 -425 195 -391
rect 161 -493 195 -459
rect 161 -561 195 -527
rect 161 -629 195 -595
rect 161 -697 195 -663
rect 161 -765 195 -731
rect 161 -833 195 -799
rect 161 -901 195 -867
rect 161 -969 195 -935
rect 161 -1037 195 -1003
rect 161 -1105 195 -1071
rect 161 -1173 195 -1139
rect 161 -1241 195 -1207
rect 161 -1309 195 -1275
rect 161 -1377 195 -1343
rect 161 -1445 195 -1411
rect 161 -1513 195 -1479
rect 161 -1581 195 -1547
rect 161 -1649 195 -1615
rect 161 -1717 195 -1683
rect 161 -1785 195 -1751
rect 161 -1853 195 -1819
rect 161 -1921 195 -1887
rect 161 -1989 195 -1955
rect 161 -2057 195 -2023
rect 161 -2125 195 -2091
rect 161 -2193 195 -2159
rect 161 -2261 195 -2227
rect 161 -2329 195 -2295
rect 161 -2397 195 -2363
rect 161 -2465 195 -2431
rect 161 -2533 195 -2499
rect 161 -2601 195 -2567
rect 161 -2669 195 -2635
rect 161 -2737 195 -2703
rect 161 -2805 195 -2771
rect 161 -2873 195 -2839
rect 161 -2941 195 -2907
rect 161 -3009 195 -2975
rect 161 -3077 195 -3043
rect 161 -3145 195 -3111
rect 161 -3213 195 -3179
rect 161 -3281 195 -3247
rect 161 -3349 195 -3315
rect 161 -3417 195 -3383
rect 161 -3485 195 -3451
rect 161 -3553 195 -3519
rect 161 -3621 195 -3587
rect 161 -3689 195 -3655
rect 161 -3757 195 -3723
rect 161 -3825 195 -3791
rect 161 -3893 195 -3859
rect 161 -3961 195 -3927
rect 161 -4029 195 -3995
rect 161 -4097 195 -4063
rect 161 -4165 195 -4131
rect 161 -4233 195 -4199
rect 161 -4301 195 -4267
rect 161 -4369 195 -4335
rect 161 -4437 195 -4403
rect 161 -4505 195 -4471
rect 161 -4573 195 -4539
rect 161 -4641 195 -4607
rect 161 -4709 195 -4675
rect 161 -4777 195 -4743
rect 161 -4845 195 -4811
rect 161 -4913 195 -4879
rect 161 -4981 195 -4947
rect -195 -5049 -161 -5015
rect -35 -5081 -17 -5047
rect 17 -5081 35 -5047
rect 161 -5049 195 -5015
rect -195 -5149 -161 -5083
rect 161 -5149 195 -5083
rect -195 -5183 -85 -5149
rect -51 -5183 -17 -5149
rect 17 -5183 51 -5149
rect 85 -5183 195 -5149
<< viali >>
rect -17 5047 17 5081
rect -81 4981 -47 4985
rect -81 4951 -47 4981
rect -81 4879 -47 4913
rect -81 4811 -47 4841
rect -81 4807 -47 4811
rect -81 4743 -47 4769
rect -81 4735 -47 4743
rect -81 4675 -47 4697
rect -81 4663 -47 4675
rect -81 4607 -47 4625
rect -81 4591 -47 4607
rect -81 4539 -47 4553
rect -81 4519 -47 4539
rect -81 4471 -47 4481
rect -81 4447 -47 4471
rect -81 4403 -47 4409
rect -81 4375 -47 4403
rect -81 4335 -47 4337
rect -81 4303 -47 4335
rect -81 4233 -47 4265
rect -81 4231 -47 4233
rect -81 4165 -47 4193
rect -81 4159 -47 4165
rect -81 4097 -47 4121
rect -81 4087 -47 4097
rect -81 4029 -47 4049
rect -81 4015 -47 4029
rect -81 3961 -47 3977
rect -81 3943 -47 3961
rect -81 3893 -47 3905
rect -81 3871 -47 3893
rect -81 3825 -47 3833
rect -81 3799 -47 3825
rect -81 3757 -47 3761
rect -81 3727 -47 3757
rect -81 3655 -47 3689
rect -81 3587 -47 3617
rect -81 3583 -47 3587
rect -81 3519 -47 3545
rect -81 3511 -47 3519
rect -81 3451 -47 3473
rect -81 3439 -47 3451
rect -81 3383 -47 3401
rect -81 3367 -47 3383
rect -81 3315 -47 3329
rect -81 3295 -47 3315
rect -81 3247 -47 3257
rect -81 3223 -47 3247
rect -81 3179 -47 3185
rect -81 3151 -47 3179
rect -81 3111 -47 3113
rect -81 3079 -47 3111
rect -81 3009 -47 3041
rect -81 3007 -47 3009
rect -81 2941 -47 2969
rect -81 2935 -47 2941
rect -81 2873 -47 2897
rect -81 2863 -47 2873
rect -81 2805 -47 2825
rect -81 2791 -47 2805
rect -81 2737 -47 2753
rect -81 2719 -47 2737
rect -81 2669 -47 2681
rect -81 2647 -47 2669
rect -81 2601 -47 2609
rect -81 2575 -47 2601
rect -81 2533 -47 2537
rect -81 2503 -47 2533
rect -81 2431 -47 2465
rect -81 2363 -47 2393
rect -81 2359 -47 2363
rect -81 2295 -47 2321
rect -81 2287 -47 2295
rect -81 2227 -47 2249
rect -81 2215 -47 2227
rect -81 2159 -47 2177
rect -81 2143 -47 2159
rect -81 2091 -47 2105
rect -81 2071 -47 2091
rect -81 2023 -47 2033
rect -81 1999 -47 2023
rect -81 1955 -47 1961
rect -81 1927 -47 1955
rect -81 1887 -47 1889
rect -81 1855 -47 1887
rect -81 1785 -47 1817
rect -81 1783 -47 1785
rect -81 1717 -47 1745
rect -81 1711 -47 1717
rect -81 1649 -47 1673
rect -81 1639 -47 1649
rect -81 1581 -47 1601
rect -81 1567 -47 1581
rect -81 1513 -47 1529
rect -81 1495 -47 1513
rect -81 1445 -47 1457
rect -81 1423 -47 1445
rect -81 1377 -47 1385
rect -81 1351 -47 1377
rect -81 1309 -47 1313
rect -81 1279 -47 1309
rect -81 1207 -47 1241
rect -81 1139 -47 1169
rect -81 1135 -47 1139
rect -81 1071 -47 1097
rect -81 1063 -47 1071
rect -81 1003 -47 1025
rect -81 991 -47 1003
rect -81 935 -47 953
rect -81 919 -47 935
rect -81 867 -47 881
rect -81 847 -47 867
rect -81 799 -47 809
rect -81 775 -47 799
rect -81 731 -47 737
rect -81 703 -47 731
rect -81 663 -47 665
rect -81 631 -47 663
rect -81 561 -47 593
rect -81 559 -47 561
rect -81 493 -47 521
rect -81 487 -47 493
rect -81 425 -47 449
rect -81 415 -47 425
rect -81 357 -47 377
rect -81 343 -47 357
rect -81 289 -47 305
rect -81 271 -47 289
rect -81 221 -47 233
rect -81 199 -47 221
rect -81 153 -47 161
rect -81 127 -47 153
rect -81 85 -47 89
rect -81 55 -47 85
rect -81 -17 -47 17
rect -81 -85 -47 -55
rect -81 -89 -47 -85
rect -81 -153 -47 -127
rect -81 -161 -47 -153
rect -81 -221 -47 -199
rect -81 -233 -47 -221
rect -81 -289 -47 -271
rect -81 -305 -47 -289
rect -81 -357 -47 -343
rect -81 -377 -47 -357
rect -81 -425 -47 -415
rect -81 -449 -47 -425
rect -81 -493 -47 -487
rect -81 -521 -47 -493
rect -81 -561 -47 -559
rect -81 -593 -47 -561
rect -81 -663 -47 -631
rect -81 -665 -47 -663
rect -81 -731 -47 -703
rect -81 -737 -47 -731
rect -81 -799 -47 -775
rect -81 -809 -47 -799
rect -81 -867 -47 -847
rect -81 -881 -47 -867
rect -81 -935 -47 -919
rect -81 -953 -47 -935
rect -81 -1003 -47 -991
rect -81 -1025 -47 -1003
rect -81 -1071 -47 -1063
rect -81 -1097 -47 -1071
rect -81 -1139 -47 -1135
rect -81 -1169 -47 -1139
rect -81 -1241 -47 -1207
rect -81 -1309 -47 -1279
rect -81 -1313 -47 -1309
rect -81 -1377 -47 -1351
rect -81 -1385 -47 -1377
rect -81 -1445 -47 -1423
rect -81 -1457 -47 -1445
rect -81 -1513 -47 -1495
rect -81 -1529 -47 -1513
rect -81 -1581 -47 -1567
rect -81 -1601 -47 -1581
rect -81 -1649 -47 -1639
rect -81 -1673 -47 -1649
rect -81 -1717 -47 -1711
rect -81 -1745 -47 -1717
rect -81 -1785 -47 -1783
rect -81 -1817 -47 -1785
rect -81 -1887 -47 -1855
rect -81 -1889 -47 -1887
rect -81 -1955 -47 -1927
rect -81 -1961 -47 -1955
rect -81 -2023 -47 -1999
rect -81 -2033 -47 -2023
rect -81 -2091 -47 -2071
rect -81 -2105 -47 -2091
rect -81 -2159 -47 -2143
rect -81 -2177 -47 -2159
rect -81 -2227 -47 -2215
rect -81 -2249 -47 -2227
rect -81 -2295 -47 -2287
rect -81 -2321 -47 -2295
rect -81 -2363 -47 -2359
rect -81 -2393 -47 -2363
rect -81 -2465 -47 -2431
rect -81 -2533 -47 -2503
rect -81 -2537 -47 -2533
rect -81 -2601 -47 -2575
rect -81 -2609 -47 -2601
rect -81 -2669 -47 -2647
rect -81 -2681 -47 -2669
rect -81 -2737 -47 -2719
rect -81 -2753 -47 -2737
rect -81 -2805 -47 -2791
rect -81 -2825 -47 -2805
rect -81 -2873 -47 -2863
rect -81 -2897 -47 -2873
rect -81 -2941 -47 -2935
rect -81 -2969 -47 -2941
rect -81 -3009 -47 -3007
rect -81 -3041 -47 -3009
rect -81 -3111 -47 -3079
rect -81 -3113 -47 -3111
rect -81 -3179 -47 -3151
rect -81 -3185 -47 -3179
rect -81 -3247 -47 -3223
rect -81 -3257 -47 -3247
rect -81 -3315 -47 -3295
rect -81 -3329 -47 -3315
rect -81 -3383 -47 -3367
rect -81 -3401 -47 -3383
rect -81 -3451 -47 -3439
rect -81 -3473 -47 -3451
rect -81 -3519 -47 -3511
rect -81 -3545 -47 -3519
rect -81 -3587 -47 -3583
rect -81 -3617 -47 -3587
rect -81 -3689 -47 -3655
rect -81 -3757 -47 -3727
rect -81 -3761 -47 -3757
rect -81 -3825 -47 -3799
rect -81 -3833 -47 -3825
rect -81 -3893 -47 -3871
rect -81 -3905 -47 -3893
rect -81 -3961 -47 -3943
rect -81 -3977 -47 -3961
rect -81 -4029 -47 -4015
rect -81 -4049 -47 -4029
rect -81 -4097 -47 -4087
rect -81 -4121 -47 -4097
rect -81 -4165 -47 -4159
rect -81 -4193 -47 -4165
rect -81 -4233 -47 -4231
rect -81 -4265 -47 -4233
rect -81 -4335 -47 -4303
rect -81 -4337 -47 -4335
rect -81 -4403 -47 -4375
rect -81 -4409 -47 -4403
rect -81 -4471 -47 -4447
rect -81 -4481 -47 -4471
rect -81 -4539 -47 -4519
rect -81 -4553 -47 -4539
rect -81 -4607 -47 -4591
rect -81 -4625 -47 -4607
rect -81 -4675 -47 -4663
rect -81 -4697 -47 -4675
rect -81 -4743 -47 -4735
rect -81 -4769 -47 -4743
rect -81 -4811 -47 -4807
rect -81 -4841 -47 -4811
rect -81 -4913 -47 -4879
rect -81 -4981 -47 -4951
rect -81 -4985 -47 -4981
rect 47 4981 81 4985
rect 47 4951 81 4981
rect 47 4879 81 4913
rect 47 4811 81 4841
rect 47 4807 81 4811
rect 47 4743 81 4769
rect 47 4735 81 4743
rect 47 4675 81 4697
rect 47 4663 81 4675
rect 47 4607 81 4625
rect 47 4591 81 4607
rect 47 4539 81 4553
rect 47 4519 81 4539
rect 47 4471 81 4481
rect 47 4447 81 4471
rect 47 4403 81 4409
rect 47 4375 81 4403
rect 47 4335 81 4337
rect 47 4303 81 4335
rect 47 4233 81 4265
rect 47 4231 81 4233
rect 47 4165 81 4193
rect 47 4159 81 4165
rect 47 4097 81 4121
rect 47 4087 81 4097
rect 47 4029 81 4049
rect 47 4015 81 4029
rect 47 3961 81 3977
rect 47 3943 81 3961
rect 47 3893 81 3905
rect 47 3871 81 3893
rect 47 3825 81 3833
rect 47 3799 81 3825
rect 47 3757 81 3761
rect 47 3727 81 3757
rect 47 3655 81 3689
rect 47 3587 81 3617
rect 47 3583 81 3587
rect 47 3519 81 3545
rect 47 3511 81 3519
rect 47 3451 81 3473
rect 47 3439 81 3451
rect 47 3383 81 3401
rect 47 3367 81 3383
rect 47 3315 81 3329
rect 47 3295 81 3315
rect 47 3247 81 3257
rect 47 3223 81 3247
rect 47 3179 81 3185
rect 47 3151 81 3179
rect 47 3111 81 3113
rect 47 3079 81 3111
rect 47 3009 81 3041
rect 47 3007 81 3009
rect 47 2941 81 2969
rect 47 2935 81 2941
rect 47 2873 81 2897
rect 47 2863 81 2873
rect 47 2805 81 2825
rect 47 2791 81 2805
rect 47 2737 81 2753
rect 47 2719 81 2737
rect 47 2669 81 2681
rect 47 2647 81 2669
rect 47 2601 81 2609
rect 47 2575 81 2601
rect 47 2533 81 2537
rect 47 2503 81 2533
rect 47 2431 81 2465
rect 47 2363 81 2393
rect 47 2359 81 2363
rect 47 2295 81 2321
rect 47 2287 81 2295
rect 47 2227 81 2249
rect 47 2215 81 2227
rect 47 2159 81 2177
rect 47 2143 81 2159
rect 47 2091 81 2105
rect 47 2071 81 2091
rect 47 2023 81 2033
rect 47 1999 81 2023
rect 47 1955 81 1961
rect 47 1927 81 1955
rect 47 1887 81 1889
rect 47 1855 81 1887
rect 47 1785 81 1817
rect 47 1783 81 1785
rect 47 1717 81 1745
rect 47 1711 81 1717
rect 47 1649 81 1673
rect 47 1639 81 1649
rect 47 1581 81 1601
rect 47 1567 81 1581
rect 47 1513 81 1529
rect 47 1495 81 1513
rect 47 1445 81 1457
rect 47 1423 81 1445
rect 47 1377 81 1385
rect 47 1351 81 1377
rect 47 1309 81 1313
rect 47 1279 81 1309
rect 47 1207 81 1241
rect 47 1139 81 1169
rect 47 1135 81 1139
rect 47 1071 81 1097
rect 47 1063 81 1071
rect 47 1003 81 1025
rect 47 991 81 1003
rect 47 935 81 953
rect 47 919 81 935
rect 47 867 81 881
rect 47 847 81 867
rect 47 799 81 809
rect 47 775 81 799
rect 47 731 81 737
rect 47 703 81 731
rect 47 663 81 665
rect 47 631 81 663
rect 47 561 81 593
rect 47 559 81 561
rect 47 493 81 521
rect 47 487 81 493
rect 47 425 81 449
rect 47 415 81 425
rect 47 357 81 377
rect 47 343 81 357
rect 47 289 81 305
rect 47 271 81 289
rect 47 221 81 233
rect 47 199 81 221
rect 47 153 81 161
rect 47 127 81 153
rect 47 85 81 89
rect 47 55 81 85
rect 47 -17 81 17
rect 47 -85 81 -55
rect 47 -89 81 -85
rect 47 -153 81 -127
rect 47 -161 81 -153
rect 47 -221 81 -199
rect 47 -233 81 -221
rect 47 -289 81 -271
rect 47 -305 81 -289
rect 47 -357 81 -343
rect 47 -377 81 -357
rect 47 -425 81 -415
rect 47 -449 81 -425
rect 47 -493 81 -487
rect 47 -521 81 -493
rect 47 -561 81 -559
rect 47 -593 81 -561
rect 47 -663 81 -631
rect 47 -665 81 -663
rect 47 -731 81 -703
rect 47 -737 81 -731
rect 47 -799 81 -775
rect 47 -809 81 -799
rect 47 -867 81 -847
rect 47 -881 81 -867
rect 47 -935 81 -919
rect 47 -953 81 -935
rect 47 -1003 81 -991
rect 47 -1025 81 -1003
rect 47 -1071 81 -1063
rect 47 -1097 81 -1071
rect 47 -1139 81 -1135
rect 47 -1169 81 -1139
rect 47 -1241 81 -1207
rect 47 -1309 81 -1279
rect 47 -1313 81 -1309
rect 47 -1377 81 -1351
rect 47 -1385 81 -1377
rect 47 -1445 81 -1423
rect 47 -1457 81 -1445
rect 47 -1513 81 -1495
rect 47 -1529 81 -1513
rect 47 -1581 81 -1567
rect 47 -1601 81 -1581
rect 47 -1649 81 -1639
rect 47 -1673 81 -1649
rect 47 -1717 81 -1711
rect 47 -1745 81 -1717
rect 47 -1785 81 -1783
rect 47 -1817 81 -1785
rect 47 -1887 81 -1855
rect 47 -1889 81 -1887
rect 47 -1955 81 -1927
rect 47 -1961 81 -1955
rect 47 -2023 81 -1999
rect 47 -2033 81 -2023
rect 47 -2091 81 -2071
rect 47 -2105 81 -2091
rect 47 -2159 81 -2143
rect 47 -2177 81 -2159
rect 47 -2227 81 -2215
rect 47 -2249 81 -2227
rect 47 -2295 81 -2287
rect 47 -2321 81 -2295
rect 47 -2363 81 -2359
rect 47 -2393 81 -2363
rect 47 -2465 81 -2431
rect 47 -2533 81 -2503
rect 47 -2537 81 -2533
rect 47 -2601 81 -2575
rect 47 -2609 81 -2601
rect 47 -2669 81 -2647
rect 47 -2681 81 -2669
rect 47 -2737 81 -2719
rect 47 -2753 81 -2737
rect 47 -2805 81 -2791
rect 47 -2825 81 -2805
rect 47 -2873 81 -2863
rect 47 -2897 81 -2873
rect 47 -2941 81 -2935
rect 47 -2969 81 -2941
rect 47 -3009 81 -3007
rect 47 -3041 81 -3009
rect 47 -3111 81 -3079
rect 47 -3113 81 -3111
rect 47 -3179 81 -3151
rect 47 -3185 81 -3179
rect 47 -3247 81 -3223
rect 47 -3257 81 -3247
rect 47 -3315 81 -3295
rect 47 -3329 81 -3315
rect 47 -3383 81 -3367
rect 47 -3401 81 -3383
rect 47 -3451 81 -3439
rect 47 -3473 81 -3451
rect 47 -3519 81 -3511
rect 47 -3545 81 -3519
rect 47 -3587 81 -3583
rect 47 -3617 81 -3587
rect 47 -3689 81 -3655
rect 47 -3757 81 -3727
rect 47 -3761 81 -3757
rect 47 -3825 81 -3799
rect 47 -3833 81 -3825
rect 47 -3893 81 -3871
rect 47 -3905 81 -3893
rect 47 -3961 81 -3943
rect 47 -3977 81 -3961
rect 47 -4029 81 -4015
rect 47 -4049 81 -4029
rect 47 -4097 81 -4087
rect 47 -4121 81 -4097
rect 47 -4165 81 -4159
rect 47 -4193 81 -4165
rect 47 -4233 81 -4231
rect 47 -4265 81 -4233
rect 47 -4335 81 -4303
rect 47 -4337 81 -4335
rect 47 -4403 81 -4375
rect 47 -4409 81 -4403
rect 47 -4471 81 -4447
rect 47 -4481 81 -4471
rect 47 -4539 81 -4519
rect 47 -4553 81 -4539
rect 47 -4607 81 -4591
rect 47 -4625 81 -4607
rect 47 -4675 81 -4663
rect 47 -4697 81 -4675
rect 47 -4743 81 -4735
rect 47 -4769 81 -4743
rect 47 -4811 81 -4807
rect 47 -4841 81 -4811
rect 47 -4913 81 -4879
rect 47 -4981 81 -4951
rect 47 -4985 81 -4981
rect -17 -5081 17 -5047
<< metal1 >>
rect -31 5081 31 5087
rect -31 5047 -17 5081
rect 17 5047 31 5081
rect -31 5041 31 5047
rect -87 4985 -41 5000
rect -87 4951 -81 4985
rect -47 4951 -41 4985
rect -87 4913 -41 4951
rect -87 4879 -81 4913
rect -47 4879 -41 4913
rect -87 4841 -41 4879
rect -87 4807 -81 4841
rect -47 4807 -41 4841
rect -87 4769 -41 4807
rect -87 4735 -81 4769
rect -47 4735 -41 4769
rect -87 4697 -41 4735
rect -87 4663 -81 4697
rect -47 4663 -41 4697
rect -87 4625 -41 4663
rect -87 4591 -81 4625
rect -47 4591 -41 4625
rect -87 4553 -41 4591
rect -87 4519 -81 4553
rect -47 4519 -41 4553
rect -87 4481 -41 4519
rect -87 4447 -81 4481
rect -47 4447 -41 4481
rect -87 4409 -41 4447
rect -87 4375 -81 4409
rect -47 4375 -41 4409
rect -87 4337 -41 4375
rect -87 4303 -81 4337
rect -47 4303 -41 4337
rect -87 4265 -41 4303
rect -87 4231 -81 4265
rect -47 4231 -41 4265
rect -87 4193 -41 4231
rect -87 4159 -81 4193
rect -47 4159 -41 4193
rect -87 4121 -41 4159
rect -87 4087 -81 4121
rect -47 4087 -41 4121
rect -87 4049 -41 4087
rect -87 4015 -81 4049
rect -47 4015 -41 4049
rect -87 3977 -41 4015
rect -87 3943 -81 3977
rect -47 3943 -41 3977
rect -87 3905 -41 3943
rect -87 3871 -81 3905
rect -47 3871 -41 3905
rect -87 3833 -41 3871
rect -87 3799 -81 3833
rect -47 3799 -41 3833
rect -87 3761 -41 3799
rect -87 3727 -81 3761
rect -47 3727 -41 3761
rect -87 3689 -41 3727
rect -87 3655 -81 3689
rect -47 3655 -41 3689
rect -87 3617 -41 3655
rect -87 3583 -81 3617
rect -47 3583 -41 3617
rect -87 3545 -41 3583
rect -87 3511 -81 3545
rect -47 3511 -41 3545
rect -87 3473 -41 3511
rect -87 3439 -81 3473
rect -47 3439 -41 3473
rect -87 3401 -41 3439
rect -87 3367 -81 3401
rect -47 3367 -41 3401
rect -87 3329 -41 3367
rect -87 3295 -81 3329
rect -47 3295 -41 3329
rect -87 3257 -41 3295
rect -87 3223 -81 3257
rect -47 3223 -41 3257
rect -87 3185 -41 3223
rect -87 3151 -81 3185
rect -47 3151 -41 3185
rect -87 3113 -41 3151
rect -87 3079 -81 3113
rect -47 3079 -41 3113
rect -87 3041 -41 3079
rect -87 3007 -81 3041
rect -47 3007 -41 3041
rect -87 2969 -41 3007
rect -87 2935 -81 2969
rect -47 2935 -41 2969
rect -87 2897 -41 2935
rect -87 2863 -81 2897
rect -47 2863 -41 2897
rect -87 2825 -41 2863
rect -87 2791 -81 2825
rect -47 2791 -41 2825
rect -87 2753 -41 2791
rect -87 2719 -81 2753
rect -47 2719 -41 2753
rect -87 2681 -41 2719
rect -87 2647 -81 2681
rect -47 2647 -41 2681
rect -87 2609 -41 2647
rect -87 2575 -81 2609
rect -47 2575 -41 2609
rect -87 2537 -41 2575
rect -87 2503 -81 2537
rect -47 2503 -41 2537
rect -87 2465 -41 2503
rect -87 2431 -81 2465
rect -47 2431 -41 2465
rect -87 2393 -41 2431
rect -87 2359 -81 2393
rect -47 2359 -41 2393
rect -87 2321 -41 2359
rect -87 2287 -81 2321
rect -47 2287 -41 2321
rect -87 2249 -41 2287
rect -87 2215 -81 2249
rect -47 2215 -41 2249
rect -87 2177 -41 2215
rect -87 2143 -81 2177
rect -47 2143 -41 2177
rect -87 2105 -41 2143
rect -87 2071 -81 2105
rect -47 2071 -41 2105
rect -87 2033 -41 2071
rect -87 1999 -81 2033
rect -47 1999 -41 2033
rect -87 1961 -41 1999
rect -87 1927 -81 1961
rect -47 1927 -41 1961
rect -87 1889 -41 1927
rect -87 1855 -81 1889
rect -47 1855 -41 1889
rect -87 1817 -41 1855
rect -87 1783 -81 1817
rect -47 1783 -41 1817
rect -87 1745 -41 1783
rect -87 1711 -81 1745
rect -47 1711 -41 1745
rect -87 1673 -41 1711
rect -87 1639 -81 1673
rect -47 1639 -41 1673
rect -87 1601 -41 1639
rect -87 1567 -81 1601
rect -47 1567 -41 1601
rect -87 1529 -41 1567
rect -87 1495 -81 1529
rect -47 1495 -41 1529
rect -87 1457 -41 1495
rect -87 1423 -81 1457
rect -47 1423 -41 1457
rect -87 1385 -41 1423
rect -87 1351 -81 1385
rect -47 1351 -41 1385
rect -87 1313 -41 1351
rect -87 1279 -81 1313
rect -47 1279 -41 1313
rect -87 1241 -41 1279
rect -87 1207 -81 1241
rect -47 1207 -41 1241
rect -87 1169 -41 1207
rect -87 1135 -81 1169
rect -47 1135 -41 1169
rect -87 1097 -41 1135
rect -87 1063 -81 1097
rect -47 1063 -41 1097
rect -87 1025 -41 1063
rect -87 991 -81 1025
rect -47 991 -41 1025
rect -87 953 -41 991
rect -87 919 -81 953
rect -47 919 -41 953
rect -87 881 -41 919
rect -87 847 -81 881
rect -47 847 -41 881
rect -87 809 -41 847
rect -87 775 -81 809
rect -47 775 -41 809
rect -87 737 -41 775
rect -87 703 -81 737
rect -47 703 -41 737
rect -87 665 -41 703
rect -87 631 -81 665
rect -47 631 -41 665
rect -87 593 -41 631
rect -87 559 -81 593
rect -47 559 -41 593
rect -87 521 -41 559
rect -87 487 -81 521
rect -47 487 -41 521
rect -87 449 -41 487
rect -87 415 -81 449
rect -47 415 -41 449
rect -87 377 -41 415
rect -87 343 -81 377
rect -47 343 -41 377
rect -87 305 -41 343
rect -87 271 -81 305
rect -47 271 -41 305
rect -87 233 -41 271
rect -87 199 -81 233
rect -47 199 -41 233
rect -87 161 -41 199
rect -87 127 -81 161
rect -47 127 -41 161
rect -87 89 -41 127
rect -87 55 -81 89
rect -47 55 -41 89
rect -87 17 -41 55
rect -87 -17 -81 17
rect -47 -17 -41 17
rect -87 -55 -41 -17
rect -87 -89 -81 -55
rect -47 -89 -41 -55
rect -87 -127 -41 -89
rect -87 -161 -81 -127
rect -47 -161 -41 -127
rect -87 -199 -41 -161
rect -87 -233 -81 -199
rect -47 -233 -41 -199
rect -87 -271 -41 -233
rect -87 -305 -81 -271
rect -47 -305 -41 -271
rect -87 -343 -41 -305
rect -87 -377 -81 -343
rect -47 -377 -41 -343
rect -87 -415 -41 -377
rect -87 -449 -81 -415
rect -47 -449 -41 -415
rect -87 -487 -41 -449
rect -87 -521 -81 -487
rect -47 -521 -41 -487
rect -87 -559 -41 -521
rect -87 -593 -81 -559
rect -47 -593 -41 -559
rect -87 -631 -41 -593
rect -87 -665 -81 -631
rect -47 -665 -41 -631
rect -87 -703 -41 -665
rect -87 -737 -81 -703
rect -47 -737 -41 -703
rect -87 -775 -41 -737
rect -87 -809 -81 -775
rect -47 -809 -41 -775
rect -87 -847 -41 -809
rect -87 -881 -81 -847
rect -47 -881 -41 -847
rect -87 -919 -41 -881
rect -87 -953 -81 -919
rect -47 -953 -41 -919
rect -87 -991 -41 -953
rect -87 -1025 -81 -991
rect -47 -1025 -41 -991
rect -87 -1063 -41 -1025
rect -87 -1097 -81 -1063
rect -47 -1097 -41 -1063
rect -87 -1135 -41 -1097
rect -87 -1169 -81 -1135
rect -47 -1169 -41 -1135
rect -87 -1207 -41 -1169
rect -87 -1241 -81 -1207
rect -47 -1241 -41 -1207
rect -87 -1279 -41 -1241
rect -87 -1313 -81 -1279
rect -47 -1313 -41 -1279
rect -87 -1351 -41 -1313
rect -87 -1385 -81 -1351
rect -47 -1385 -41 -1351
rect -87 -1423 -41 -1385
rect -87 -1457 -81 -1423
rect -47 -1457 -41 -1423
rect -87 -1495 -41 -1457
rect -87 -1529 -81 -1495
rect -47 -1529 -41 -1495
rect -87 -1567 -41 -1529
rect -87 -1601 -81 -1567
rect -47 -1601 -41 -1567
rect -87 -1639 -41 -1601
rect -87 -1673 -81 -1639
rect -47 -1673 -41 -1639
rect -87 -1711 -41 -1673
rect -87 -1745 -81 -1711
rect -47 -1745 -41 -1711
rect -87 -1783 -41 -1745
rect -87 -1817 -81 -1783
rect -47 -1817 -41 -1783
rect -87 -1855 -41 -1817
rect -87 -1889 -81 -1855
rect -47 -1889 -41 -1855
rect -87 -1927 -41 -1889
rect -87 -1961 -81 -1927
rect -47 -1961 -41 -1927
rect -87 -1999 -41 -1961
rect -87 -2033 -81 -1999
rect -47 -2033 -41 -1999
rect -87 -2071 -41 -2033
rect -87 -2105 -81 -2071
rect -47 -2105 -41 -2071
rect -87 -2143 -41 -2105
rect -87 -2177 -81 -2143
rect -47 -2177 -41 -2143
rect -87 -2215 -41 -2177
rect -87 -2249 -81 -2215
rect -47 -2249 -41 -2215
rect -87 -2287 -41 -2249
rect -87 -2321 -81 -2287
rect -47 -2321 -41 -2287
rect -87 -2359 -41 -2321
rect -87 -2393 -81 -2359
rect -47 -2393 -41 -2359
rect -87 -2431 -41 -2393
rect -87 -2465 -81 -2431
rect -47 -2465 -41 -2431
rect -87 -2503 -41 -2465
rect -87 -2537 -81 -2503
rect -47 -2537 -41 -2503
rect -87 -2575 -41 -2537
rect -87 -2609 -81 -2575
rect -47 -2609 -41 -2575
rect -87 -2647 -41 -2609
rect -87 -2681 -81 -2647
rect -47 -2681 -41 -2647
rect -87 -2719 -41 -2681
rect -87 -2753 -81 -2719
rect -47 -2753 -41 -2719
rect -87 -2791 -41 -2753
rect -87 -2825 -81 -2791
rect -47 -2825 -41 -2791
rect -87 -2863 -41 -2825
rect -87 -2897 -81 -2863
rect -47 -2897 -41 -2863
rect -87 -2935 -41 -2897
rect -87 -2969 -81 -2935
rect -47 -2969 -41 -2935
rect -87 -3007 -41 -2969
rect -87 -3041 -81 -3007
rect -47 -3041 -41 -3007
rect -87 -3079 -41 -3041
rect -87 -3113 -81 -3079
rect -47 -3113 -41 -3079
rect -87 -3151 -41 -3113
rect -87 -3185 -81 -3151
rect -47 -3185 -41 -3151
rect -87 -3223 -41 -3185
rect -87 -3257 -81 -3223
rect -47 -3257 -41 -3223
rect -87 -3295 -41 -3257
rect -87 -3329 -81 -3295
rect -47 -3329 -41 -3295
rect -87 -3367 -41 -3329
rect -87 -3401 -81 -3367
rect -47 -3401 -41 -3367
rect -87 -3439 -41 -3401
rect -87 -3473 -81 -3439
rect -47 -3473 -41 -3439
rect -87 -3511 -41 -3473
rect -87 -3545 -81 -3511
rect -47 -3545 -41 -3511
rect -87 -3583 -41 -3545
rect -87 -3617 -81 -3583
rect -47 -3617 -41 -3583
rect -87 -3655 -41 -3617
rect -87 -3689 -81 -3655
rect -47 -3689 -41 -3655
rect -87 -3727 -41 -3689
rect -87 -3761 -81 -3727
rect -47 -3761 -41 -3727
rect -87 -3799 -41 -3761
rect -87 -3833 -81 -3799
rect -47 -3833 -41 -3799
rect -87 -3871 -41 -3833
rect -87 -3905 -81 -3871
rect -47 -3905 -41 -3871
rect -87 -3943 -41 -3905
rect -87 -3977 -81 -3943
rect -47 -3977 -41 -3943
rect -87 -4015 -41 -3977
rect -87 -4049 -81 -4015
rect -47 -4049 -41 -4015
rect -87 -4087 -41 -4049
rect -87 -4121 -81 -4087
rect -47 -4121 -41 -4087
rect -87 -4159 -41 -4121
rect -87 -4193 -81 -4159
rect -47 -4193 -41 -4159
rect -87 -4231 -41 -4193
rect -87 -4265 -81 -4231
rect -47 -4265 -41 -4231
rect -87 -4303 -41 -4265
rect -87 -4337 -81 -4303
rect -47 -4337 -41 -4303
rect -87 -4375 -41 -4337
rect -87 -4409 -81 -4375
rect -47 -4409 -41 -4375
rect -87 -4447 -41 -4409
rect -87 -4481 -81 -4447
rect -47 -4481 -41 -4447
rect -87 -4519 -41 -4481
rect -87 -4553 -81 -4519
rect -47 -4553 -41 -4519
rect -87 -4591 -41 -4553
rect -87 -4625 -81 -4591
rect -47 -4625 -41 -4591
rect -87 -4663 -41 -4625
rect -87 -4697 -81 -4663
rect -47 -4697 -41 -4663
rect -87 -4735 -41 -4697
rect -87 -4769 -81 -4735
rect -47 -4769 -41 -4735
rect -87 -4807 -41 -4769
rect -87 -4841 -81 -4807
rect -47 -4841 -41 -4807
rect -87 -4879 -41 -4841
rect -87 -4913 -81 -4879
rect -47 -4913 -41 -4879
rect -87 -4951 -41 -4913
rect -87 -4985 -81 -4951
rect -47 -4985 -41 -4951
rect -87 -5000 -41 -4985
rect 41 4985 87 5000
rect 41 4951 47 4985
rect 81 4951 87 4985
rect 41 4913 87 4951
rect 41 4879 47 4913
rect 81 4879 87 4913
rect 41 4841 87 4879
rect 41 4807 47 4841
rect 81 4807 87 4841
rect 41 4769 87 4807
rect 41 4735 47 4769
rect 81 4735 87 4769
rect 41 4697 87 4735
rect 41 4663 47 4697
rect 81 4663 87 4697
rect 41 4625 87 4663
rect 41 4591 47 4625
rect 81 4591 87 4625
rect 41 4553 87 4591
rect 41 4519 47 4553
rect 81 4519 87 4553
rect 41 4481 87 4519
rect 41 4447 47 4481
rect 81 4447 87 4481
rect 41 4409 87 4447
rect 41 4375 47 4409
rect 81 4375 87 4409
rect 41 4337 87 4375
rect 41 4303 47 4337
rect 81 4303 87 4337
rect 41 4265 87 4303
rect 41 4231 47 4265
rect 81 4231 87 4265
rect 41 4193 87 4231
rect 41 4159 47 4193
rect 81 4159 87 4193
rect 41 4121 87 4159
rect 41 4087 47 4121
rect 81 4087 87 4121
rect 41 4049 87 4087
rect 41 4015 47 4049
rect 81 4015 87 4049
rect 41 3977 87 4015
rect 41 3943 47 3977
rect 81 3943 87 3977
rect 41 3905 87 3943
rect 41 3871 47 3905
rect 81 3871 87 3905
rect 41 3833 87 3871
rect 41 3799 47 3833
rect 81 3799 87 3833
rect 41 3761 87 3799
rect 41 3727 47 3761
rect 81 3727 87 3761
rect 41 3689 87 3727
rect 41 3655 47 3689
rect 81 3655 87 3689
rect 41 3617 87 3655
rect 41 3583 47 3617
rect 81 3583 87 3617
rect 41 3545 87 3583
rect 41 3511 47 3545
rect 81 3511 87 3545
rect 41 3473 87 3511
rect 41 3439 47 3473
rect 81 3439 87 3473
rect 41 3401 87 3439
rect 41 3367 47 3401
rect 81 3367 87 3401
rect 41 3329 87 3367
rect 41 3295 47 3329
rect 81 3295 87 3329
rect 41 3257 87 3295
rect 41 3223 47 3257
rect 81 3223 87 3257
rect 41 3185 87 3223
rect 41 3151 47 3185
rect 81 3151 87 3185
rect 41 3113 87 3151
rect 41 3079 47 3113
rect 81 3079 87 3113
rect 41 3041 87 3079
rect 41 3007 47 3041
rect 81 3007 87 3041
rect 41 2969 87 3007
rect 41 2935 47 2969
rect 81 2935 87 2969
rect 41 2897 87 2935
rect 41 2863 47 2897
rect 81 2863 87 2897
rect 41 2825 87 2863
rect 41 2791 47 2825
rect 81 2791 87 2825
rect 41 2753 87 2791
rect 41 2719 47 2753
rect 81 2719 87 2753
rect 41 2681 87 2719
rect 41 2647 47 2681
rect 81 2647 87 2681
rect 41 2609 87 2647
rect 41 2575 47 2609
rect 81 2575 87 2609
rect 41 2537 87 2575
rect 41 2503 47 2537
rect 81 2503 87 2537
rect 41 2465 87 2503
rect 41 2431 47 2465
rect 81 2431 87 2465
rect 41 2393 87 2431
rect 41 2359 47 2393
rect 81 2359 87 2393
rect 41 2321 87 2359
rect 41 2287 47 2321
rect 81 2287 87 2321
rect 41 2249 87 2287
rect 41 2215 47 2249
rect 81 2215 87 2249
rect 41 2177 87 2215
rect 41 2143 47 2177
rect 81 2143 87 2177
rect 41 2105 87 2143
rect 41 2071 47 2105
rect 81 2071 87 2105
rect 41 2033 87 2071
rect 41 1999 47 2033
rect 81 1999 87 2033
rect 41 1961 87 1999
rect 41 1927 47 1961
rect 81 1927 87 1961
rect 41 1889 87 1927
rect 41 1855 47 1889
rect 81 1855 87 1889
rect 41 1817 87 1855
rect 41 1783 47 1817
rect 81 1783 87 1817
rect 41 1745 87 1783
rect 41 1711 47 1745
rect 81 1711 87 1745
rect 41 1673 87 1711
rect 41 1639 47 1673
rect 81 1639 87 1673
rect 41 1601 87 1639
rect 41 1567 47 1601
rect 81 1567 87 1601
rect 41 1529 87 1567
rect 41 1495 47 1529
rect 81 1495 87 1529
rect 41 1457 87 1495
rect 41 1423 47 1457
rect 81 1423 87 1457
rect 41 1385 87 1423
rect 41 1351 47 1385
rect 81 1351 87 1385
rect 41 1313 87 1351
rect 41 1279 47 1313
rect 81 1279 87 1313
rect 41 1241 87 1279
rect 41 1207 47 1241
rect 81 1207 87 1241
rect 41 1169 87 1207
rect 41 1135 47 1169
rect 81 1135 87 1169
rect 41 1097 87 1135
rect 41 1063 47 1097
rect 81 1063 87 1097
rect 41 1025 87 1063
rect 41 991 47 1025
rect 81 991 87 1025
rect 41 953 87 991
rect 41 919 47 953
rect 81 919 87 953
rect 41 881 87 919
rect 41 847 47 881
rect 81 847 87 881
rect 41 809 87 847
rect 41 775 47 809
rect 81 775 87 809
rect 41 737 87 775
rect 41 703 47 737
rect 81 703 87 737
rect 41 665 87 703
rect 41 631 47 665
rect 81 631 87 665
rect 41 593 87 631
rect 41 559 47 593
rect 81 559 87 593
rect 41 521 87 559
rect 41 487 47 521
rect 81 487 87 521
rect 41 449 87 487
rect 41 415 47 449
rect 81 415 87 449
rect 41 377 87 415
rect 41 343 47 377
rect 81 343 87 377
rect 41 305 87 343
rect 41 271 47 305
rect 81 271 87 305
rect 41 233 87 271
rect 41 199 47 233
rect 81 199 87 233
rect 41 161 87 199
rect 41 127 47 161
rect 81 127 87 161
rect 41 89 87 127
rect 41 55 47 89
rect 81 55 87 89
rect 41 17 87 55
rect 41 -17 47 17
rect 81 -17 87 17
rect 41 -55 87 -17
rect 41 -89 47 -55
rect 81 -89 87 -55
rect 41 -127 87 -89
rect 41 -161 47 -127
rect 81 -161 87 -127
rect 41 -199 87 -161
rect 41 -233 47 -199
rect 81 -233 87 -199
rect 41 -271 87 -233
rect 41 -305 47 -271
rect 81 -305 87 -271
rect 41 -343 87 -305
rect 41 -377 47 -343
rect 81 -377 87 -343
rect 41 -415 87 -377
rect 41 -449 47 -415
rect 81 -449 87 -415
rect 41 -487 87 -449
rect 41 -521 47 -487
rect 81 -521 87 -487
rect 41 -559 87 -521
rect 41 -593 47 -559
rect 81 -593 87 -559
rect 41 -631 87 -593
rect 41 -665 47 -631
rect 81 -665 87 -631
rect 41 -703 87 -665
rect 41 -737 47 -703
rect 81 -737 87 -703
rect 41 -775 87 -737
rect 41 -809 47 -775
rect 81 -809 87 -775
rect 41 -847 87 -809
rect 41 -881 47 -847
rect 81 -881 87 -847
rect 41 -919 87 -881
rect 41 -953 47 -919
rect 81 -953 87 -919
rect 41 -991 87 -953
rect 41 -1025 47 -991
rect 81 -1025 87 -991
rect 41 -1063 87 -1025
rect 41 -1097 47 -1063
rect 81 -1097 87 -1063
rect 41 -1135 87 -1097
rect 41 -1169 47 -1135
rect 81 -1169 87 -1135
rect 41 -1207 87 -1169
rect 41 -1241 47 -1207
rect 81 -1241 87 -1207
rect 41 -1279 87 -1241
rect 41 -1313 47 -1279
rect 81 -1313 87 -1279
rect 41 -1351 87 -1313
rect 41 -1385 47 -1351
rect 81 -1385 87 -1351
rect 41 -1423 87 -1385
rect 41 -1457 47 -1423
rect 81 -1457 87 -1423
rect 41 -1495 87 -1457
rect 41 -1529 47 -1495
rect 81 -1529 87 -1495
rect 41 -1567 87 -1529
rect 41 -1601 47 -1567
rect 81 -1601 87 -1567
rect 41 -1639 87 -1601
rect 41 -1673 47 -1639
rect 81 -1673 87 -1639
rect 41 -1711 87 -1673
rect 41 -1745 47 -1711
rect 81 -1745 87 -1711
rect 41 -1783 87 -1745
rect 41 -1817 47 -1783
rect 81 -1817 87 -1783
rect 41 -1855 87 -1817
rect 41 -1889 47 -1855
rect 81 -1889 87 -1855
rect 41 -1927 87 -1889
rect 41 -1961 47 -1927
rect 81 -1961 87 -1927
rect 41 -1999 87 -1961
rect 41 -2033 47 -1999
rect 81 -2033 87 -1999
rect 41 -2071 87 -2033
rect 41 -2105 47 -2071
rect 81 -2105 87 -2071
rect 41 -2143 87 -2105
rect 41 -2177 47 -2143
rect 81 -2177 87 -2143
rect 41 -2215 87 -2177
rect 41 -2249 47 -2215
rect 81 -2249 87 -2215
rect 41 -2287 87 -2249
rect 41 -2321 47 -2287
rect 81 -2321 87 -2287
rect 41 -2359 87 -2321
rect 41 -2393 47 -2359
rect 81 -2393 87 -2359
rect 41 -2431 87 -2393
rect 41 -2465 47 -2431
rect 81 -2465 87 -2431
rect 41 -2503 87 -2465
rect 41 -2537 47 -2503
rect 81 -2537 87 -2503
rect 41 -2575 87 -2537
rect 41 -2609 47 -2575
rect 81 -2609 87 -2575
rect 41 -2647 87 -2609
rect 41 -2681 47 -2647
rect 81 -2681 87 -2647
rect 41 -2719 87 -2681
rect 41 -2753 47 -2719
rect 81 -2753 87 -2719
rect 41 -2791 87 -2753
rect 41 -2825 47 -2791
rect 81 -2825 87 -2791
rect 41 -2863 87 -2825
rect 41 -2897 47 -2863
rect 81 -2897 87 -2863
rect 41 -2935 87 -2897
rect 41 -2969 47 -2935
rect 81 -2969 87 -2935
rect 41 -3007 87 -2969
rect 41 -3041 47 -3007
rect 81 -3041 87 -3007
rect 41 -3079 87 -3041
rect 41 -3113 47 -3079
rect 81 -3113 87 -3079
rect 41 -3151 87 -3113
rect 41 -3185 47 -3151
rect 81 -3185 87 -3151
rect 41 -3223 87 -3185
rect 41 -3257 47 -3223
rect 81 -3257 87 -3223
rect 41 -3295 87 -3257
rect 41 -3329 47 -3295
rect 81 -3329 87 -3295
rect 41 -3367 87 -3329
rect 41 -3401 47 -3367
rect 81 -3401 87 -3367
rect 41 -3439 87 -3401
rect 41 -3473 47 -3439
rect 81 -3473 87 -3439
rect 41 -3511 87 -3473
rect 41 -3545 47 -3511
rect 81 -3545 87 -3511
rect 41 -3583 87 -3545
rect 41 -3617 47 -3583
rect 81 -3617 87 -3583
rect 41 -3655 87 -3617
rect 41 -3689 47 -3655
rect 81 -3689 87 -3655
rect 41 -3727 87 -3689
rect 41 -3761 47 -3727
rect 81 -3761 87 -3727
rect 41 -3799 87 -3761
rect 41 -3833 47 -3799
rect 81 -3833 87 -3799
rect 41 -3871 87 -3833
rect 41 -3905 47 -3871
rect 81 -3905 87 -3871
rect 41 -3943 87 -3905
rect 41 -3977 47 -3943
rect 81 -3977 87 -3943
rect 41 -4015 87 -3977
rect 41 -4049 47 -4015
rect 81 -4049 87 -4015
rect 41 -4087 87 -4049
rect 41 -4121 47 -4087
rect 81 -4121 87 -4087
rect 41 -4159 87 -4121
rect 41 -4193 47 -4159
rect 81 -4193 87 -4159
rect 41 -4231 87 -4193
rect 41 -4265 47 -4231
rect 81 -4265 87 -4231
rect 41 -4303 87 -4265
rect 41 -4337 47 -4303
rect 81 -4337 87 -4303
rect 41 -4375 87 -4337
rect 41 -4409 47 -4375
rect 81 -4409 87 -4375
rect 41 -4447 87 -4409
rect 41 -4481 47 -4447
rect 81 -4481 87 -4447
rect 41 -4519 87 -4481
rect 41 -4553 47 -4519
rect 81 -4553 87 -4519
rect 41 -4591 87 -4553
rect 41 -4625 47 -4591
rect 81 -4625 87 -4591
rect 41 -4663 87 -4625
rect 41 -4697 47 -4663
rect 81 -4697 87 -4663
rect 41 -4735 87 -4697
rect 41 -4769 47 -4735
rect 81 -4769 87 -4735
rect 41 -4807 87 -4769
rect 41 -4841 47 -4807
rect 81 -4841 87 -4807
rect 41 -4879 87 -4841
rect 41 -4913 47 -4879
rect 81 -4913 87 -4879
rect 41 -4951 87 -4913
rect 41 -4985 47 -4951
rect 81 -4985 87 -4951
rect 41 -5000 87 -4985
rect -31 -5047 31 -5041
rect -31 -5081 -17 -5047
rect 17 -5081 31 -5047
rect -31 -5087 31 -5081
<< properties >>
string FIXED_BBOX -178 -5166 178 5166
<< end >>
