magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< error_p >>
rect -73 -400 -15 400
rect 15 -400 73 400
<< pwell >>
rect -99 -426 99 426
<< nmoslvt >>
rect -15 -400 15 400
<< ndiff >>
rect -73 357 -15 400
rect -73 323 -61 357
rect -27 323 -15 357
rect -73 289 -15 323
rect -73 255 -61 289
rect -27 255 -15 289
rect -73 221 -15 255
rect -73 187 -61 221
rect -27 187 -15 221
rect -73 153 -15 187
rect -73 119 -61 153
rect -27 119 -15 153
rect -73 85 -15 119
rect -73 51 -61 85
rect -27 51 -15 85
rect -73 17 -15 51
rect -73 -17 -61 17
rect -27 -17 -15 17
rect -73 -51 -15 -17
rect -73 -85 -61 -51
rect -27 -85 -15 -51
rect -73 -119 -15 -85
rect -73 -153 -61 -119
rect -27 -153 -15 -119
rect -73 -187 -15 -153
rect -73 -221 -61 -187
rect -27 -221 -15 -187
rect -73 -255 -15 -221
rect -73 -289 -61 -255
rect -27 -289 -15 -255
rect -73 -323 -15 -289
rect -73 -357 -61 -323
rect -27 -357 -15 -323
rect -73 -400 -15 -357
rect 15 357 73 400
rect 15 323 27 357
rect 61 323 73 357
rect 15 289 73 323
rect 15 255 27 289
rect 61 255 73 289
rect 15 221 73 255
rect 15 187 27 221
rect 61 187 73 221
rect 15 153 73 187
rect 15 119 27 153
rect 61 119 73 153
rect 15 85 73 119
rect 15 51 27 85
rect 61 51 73 85
rect 15 17 73 51
rect 15 -17 27 17
rect 61 -17 73 17
rect 15 -51 73 -17
rect 15 -85 27 -51
rect 61 -85 73 -51
rect 15 -119 73 -85
rect 15 -153 27 -119
rect 61 -153 73 -119
rect 15 -187 73 -153
rect 15 -221 27 -187
rect 61 -221 73 -187
rect 15 -255 73 -221
rect 15 -289 27 -255
rect 61 -289 73 -255
rect 15 -323 73 -289
rect 15 -357 27 -323
rect 61 -357 73 -323
rect 15 -400 73 -357
<< ndiffc >>
rect -61 323 -27 357
rect -61 255 -27 289
rect -61 187 -27 221
rect -61 119 -27 153
rect -61 51 -27 85
rect -61 -17 -27 17
rect -61 -85 -27 -51
rect -61 -153 -27 -119
rect -61 -221 -27 -187
rect -61 -289 -27 -255
rect -61 -357 -27 -323
rect 27 323 61 357
rect 27 255 61 289
rect 27 187 61 221
rect 27 119 61 153
rect 27 51 61 85
rect 27 -17 61 17
rect 27 -85 61 -51
rect 27 -153 61 -119
rect 27 -221 61 -187
rect 27 -289 61 -255
rect 27 -357 61 -323
<< poly >>
rect -15 400 15 426
rect -15 -426 15 -400
<< locali >>
rect -61 377 -27 404
rect -61 305 -27 323
rect -61 233 -27 255
rect -61 161 -27 187
rect -61 89 -27 119
rect -61 17 -27 51
rect -61 -51 -27 -17
rect -61 -119 -27 -89
rect -61 -187 -27 -161
rect -61 -255 -27 -233
rect -61 -323 -27 -305
rect -61 -404 -27 -377
rect 27 377 61 404
rect 27 305 61 323
rect 27 233 61 255
rect 27 161 61 187
rect 27 89 61 119
rect 27 17 61 51
rect 27 -51 61 -17
rect 27 -119 61 -89
rect 27 -187 61 -161
rect 27 -255 61 -233
rect 27 -323 61 -305
rect 27 -404 61 -377
<< viali >>
rect -61 357 -27 377
rect -61 343 -27 357
rect -61 289 -27 305
rect -61 271 -27 289
rect -61 221 -27 233
rect -61 199 -27 221
rect -61 153 -27 161
rect -61 127 -27 153
rect -61 85 -27 89
rect -61 55 -27 85
rect -61 -17 -27 17
rect -61 -85 -27 -55
rect -61 -89 -27 -85
rect -61 -153 -27 -127
rect -61 -161 -27 -153
rect -61 -221 -27 -199
rect -61 -233 -27 -221
rect -61 -289 -27 -271
rect -61 -305 -27 -289
rect -61 -357 -27 -343
rect -61 -377 -27 -357
rect 27 357 61 377
rect 27 343 61 357
rect 27 289 61 305
rect 27 271 61 289
rect 27 221 61 233
rect 27 199 61 221
rect 27 153 61 161
rect 27 127 61 153
rect 27 85 61 89
rect 27 55 61 85
rect 27 -17 61 17
rect 27 -85 61 -55
rect 27 -89 61 -85
rect 27 -153 61 -127
rect 27 -161 61 -153
rect 27 -221 61 -199
rect 27 -233 61 -221
rect 27 -289 61 -271
rect 27 -305 61 -289
rect 27 -357 61 -343
rect 27 -377 61 -357
<< metal1 >>
rect -67 377 -21 400
rect -67 343 -61 377
rect -27 343 -21 377
rect -67 305 -21 343
rect -67 271 -61 305
rect -27 271 -21 305
rect -67 233 -21 271
rect -67 199 -61 233
rect -27 199 -21 233
rect -67 161 -21 199
rect -67 127 -61 161
rect -27 127 -21 161
rect -67 89 -21 127
rect -67 55 -61 89
rect -27 55 -21 89
rect -67 17 -21 55
rect -67 -17 -61 17
rect -27 -17 -21 17
rect -67 -55 -21 -17
rect -67 -89 -61 -55
rect -27 -89 -21 -55
rect -67 -127 -21 -89
rect -67 -161 -61 -127
rect -27 -161 -21 -127
rect -67 -199 -21 -161
rect -67 -233 -61 -199
rect -27 -233 -21 -199
rect -67 -271 -21 -233
rect -67 -305 -61 -271
rect -27 -305 -21 -271
rect -67 -343 -21 -305
rect -67 -377 -61 -343
rect -27 -377 -21 -343
rect -67 -400 -21 -377
rect 21 377 67 400
rect 21 343 27 377
rect 61 343 67 377
rect 21 305 67 343
rect 21 271 27 305
rect 61 271 67 305
rect 21 233 67 271
rect 21 199 27 233
rect 61 199 67 233
rect 21 161 67 199
rect 21 127 27 161
rect 61 127 67 161
rect 21 89 67 127
rect 21 55 27 89
rect 61 55 67 89
rect 21 17 67 55
rect 21 -17 27 17
rect 61 -17 67 17
rect 21 -55 67 -17
rect 21 -89 27 -55
rect 61 -89 67 -55
rect 21 -127 67 -89
rect 21 -161 27 -127
rect 61 -161 67 -127
rect 21 -199 67 -161
rect 21 -233 27 -199
rect 61 -233 67 -199
rect 21 -271 67 -233
rect 21 -305 27 -271
rect 61 -305 67 -271
rect 21 -343 67 -305
rect 21 -377 27 -343
rect 61 -377 67 -343
rect 21 -400 67 -377
<< end >>
