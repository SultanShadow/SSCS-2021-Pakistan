magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< nwell >>
rect 4063 236 5520 3108
<< pwell >>
rect 3117 3362 3781 3484
<< pmos >>
rect 4336 591 4366 2591
rect 4424 591 4454 2591
rect 4512 591 4542 2591
rect 4600 591 4630 2591
rect 4688 591 4718 2591
rect 4776 591 4806 2591
rect 4864 591 4894 2591
rect 4952 591 4982 2591
rect 5040 591 5070 2591
rect 5128 591 5158 2591
rect 5216 591 5246 2591
<< pdiff >>
rect 4278 2560 4336 2591
rect 4278 2526 4290 2560
rect 4324 2526 4336 2560
rect 4278 2492 4336 2526
rect 4278 2458 4290 2492
rect 4324 2458 4336 2492
rect 4278 2424 4336 2458
rect 4278 2390 4290 2424
rect 4324 2390 4336 2424
rect 4278 2356 4336 2390
rect 4278 2322 4290 2356
rect 4324 2322 4336 2356
rect 4278 2288 4336 2322
rect 4278 2254 4290 2288
rect 4324 2254 4336 2288
rect 4278 2220 4336 2254
rect 4278 2186 4290 2220
rect 4324 2186 4336 2220
rect 4278 2152 4336 2186
rect 4278 2118 4290 2152
rect 4324 2118 4336 2152
rect 4278 2084 4336 2118
rect 4278 2050 4290 2084
rect 4324 2050 4336 2084
rect 4278 2016 4336 2050
rect 4278 1982 4290 2016
rect 4324 1982 4336 2016
rect 4278 1948 4336 1982
rect 4278 1914 4290 1948
rect 4324 1914 4336 1948
rect 4278 1880 4336 1914
rect 4278 1846 4290 1880
rect 4324 1846 4336 1880
rect 4278 1812 4336 1846
rect 4278 1778 4290 1812
rect 4324 1778 4336 1812
rect 4278 1744 4336 1778
rect 4278 1710 4290 1744
rect 4324 1710 4336 1744
rect 4278 1676 4336 1710
rect 4278 1642 4290 1676
rect 4324 1642 4336 1676
rect 4278 1608 4336 1642
rect 4278 1574 4290 1608
rect 4324 1574 4336 1608
rect 4278 1540 4336 1574
rect 4278 1506 4290 1540
rect 4324 1506 4336 1540
rect 4278 1472 4336 1506
rect 4278 1438 4290 1472
rect 4324 1438 4336 1472
rect 4278 1404 4336 1438
rect 4278 1370 4290 1404
rect 4324 1370 4336 1404
rect 4278 1336 4336 1370
rect 4278 1302 4290 1336
rect 4324 1302 4336 1336
rect 4278 1268 4336 1302
rect 4278 1234 4290 1268
rect 4324 1234 4336 1268
rect 4278 1200 4336 1234
rect 4278 1166 4290 1200
rect 4324 1166 4336 1200
rect 4278 1132 4336 1166
rect 4278 1098 4290 1132
rect 4324 1098 4336 1132
rect 4278 1064 4336 1098
rect 4278 1030 4290 1064
rect 4324 1030 4336 1064
rect 4278 996 4336 1030
rect 4278 962 4290 996
rect 4324 962 4336 996
rect 4278 928 4336 962
rect 4278 894 4290 928
rect 4324 894 4336 928
rect 4278 860 4336 894
rect 4278 826 4290 860
rect 4324 826 4336 860
rect 4278 792 4336 826
rect 4278 758 4290 792
rect 4324 758 4336 792
rect 4278 724 4336 758
rect 4278 690 4290 724
rect 4324 690 4336 724
rect 4278 656 4336 690
rect 4278 622 4290 656
rect 4324 622 4336 656
rect 4278 591 4336 622
rect 4366 2560 4424 2591
rect 4366 2526 4378 2560
rect 4412 2526 4424 2560
rect 4366 2492 4424 2526
rect 4366 2458 4378 2492
rect 4412 2458 4424 2492
rect 4366 2424 4424 2458
rect 4366 2390 4378 2424
rect 4412 2390 4424 2424
rect 4366 2356 4424 2390
rect 4366 2322 4378 2356
rect 4412 2322 4424 2356
rect 4366 2288 4424 2322
rect 4366 2254 4378 2288
rect 4412 2254 4424 2288
rect 4366 2220 4424 2254
rect 4366 2186 4378 2220
rect 4412 2186 4424 2220
rect 4366 2152 4424 2186
rect 4366 2118 4378 2152
rect 4412 2118 4424 2152
rect 4366 2084 4424 2118
rect 4366 2050 4378 2084
rect 4412 2050 4424 2084
rect 4366 2016 4424 2050
rect 4366 1982 4378 2016
rect 4412 1982 4424 2016
rect 4366 1948 4424 1982
rect 4366 1914 4378 1948
rect 4412 1914 4424 1948
rect 4366 1880 4424 1914
rect 4366 1846 4378 1880
rect 4412 1846 4424 1880
rect 4366 1812 4424 1846
rect 4366 1778 4378 1812
rect 4412 1778 4424 1812
rect 4366 1744 4424 1778
rect 4366 1710 4378 1744
rect 4412 1710 4424 1744
rect 4366 1676 4424 1710
rect 4366 1642 4378 1676
rect 4412 1642 4424 1676
rect 4366 1608 4424 1642
rect 4366 1574 4378 1608
rect 4412 1574 4424 1608
rect 4366 1540 4424 1574
rect 4366 1506 4378 1540
rect 4412 1506 4424 1540
rect 4366 1472 4424 1506
rect 4366 1438 4378 1472
rect 4412 1438 4424 1472
rect 4366 1404 4424 1438
rect 4366 1370 4378 1404
rect 4412 1370 4424 1404
rect 4366 1336 4424 1370
rect 4366 1302 4378 1336
rect 4412 1302 4424 1336
rect 4366 1268 4424 1302
rect 4366 1234 4378 1268
rect 4412 1234 4424 1268
rect 4366 1200 4424 1234
rect 4366 1166 4378 1200
rect 4412 1166 4424 1200
rect 4366 1132 4424 1166
rect 4366 1098 4378 1132
rect 4412 1098 4424 1132
rect 4366 1064 4424 1098
rect 4366 1030 4378 1064
rect 4412 1030 4424 1064
rect 4366 996 4424 1030
rect 4366 962 4378 996
rect 4412 962 4424 996
rect 4366 928 4424 962
rect 4366 894 4378 928
rect 4412 894 4424 928
rect 4366 860 4424 894
rect 4366 826 4378 860
rect 4412 826 4424 860
rect 4366 792 4424 826
rect 4366 758 4378 792
rect 4412 758 4424 792
rect 4366 724 4424 758
rect 4366 690 4378 724
rect 4412 690 4424 724
rect 4366 656 4424 690
rect 4366 622 4378 656
rect 4412 622 4424 656
rect 4366 591 4424 622
rect 4454 2560 4512 2591
rect 4454 2526 4466 2560
rect 4500 2526 4512 2560
rect 4454 2492 4512 2526
rect 4454 2458 4466 2492
rect 4500 2458 4512 2492
rect 4454 2424 4512 2458
rect 4454 2390 4466 2424
rect 4500 2390 4512 2424
rect 4454 2356 4512 2390
rect 4454 2322 4466 2356
rect 4500 2322 4512 2356
rect 4454 2288 4512 2322
rect 4454 2254 4466 2288
rect 4500 2254 4512 2288
rect 4454 2220 4512 2254
rect 4454 2186 4466 2220
rect 4500 2186 4512 2220
rect 4454 2152 4512 2186
rect 4454 2118 4466 2152
rect 4500 2118 4512 2152
rect 4454 2084 4512 2118
rect 4454 2050 4466 2084
rect 4500 2050 4512 2084
rect 4454 2016 4512 2050
rect 4454 1982 4466 2016
rect 4500 1982 4512 2016
rect 4454 1948 4512 1982
rect 4454 1914 4466 1948
rect 4500 1914 4512 1948
rect 4454 1880 4512 1914
rect 4454 1846 4466 1880
rect 4500 1846 4512 1880
rect 4454 1812 4512 1846
rect 4454 1778 4466 1812
rect 4500 1778 4512 1812
rect 4454 1744 4512 1778
rect 4454 1710 4466 1744
rect 4500 1710 4512 1744
rect 4454 1676 4512 1710
rect 4454 1642 4466 1676
rect 4500 1642 4512 1676
rect 4454 1608 4512 1642
rect 4454 1574 4466 1608
rect 4500 1574 4512 1608
rect 4454 1540 4512 1574
rect 4454 1506 4466 1540
rect 4500 1506 4512 1540
rect 4454 1472 4512 1506
rect 4454 1438 4466 1472
rect 4500 1438 4512 1472
rect 4454 1404 4512 1438
rect 4454 1370 4466 1404
rect 4500 1370 4512 1404
rect 4454 1336 4512 1370
rect 4454 1302 4466 1336
rect 4500 1302 4512 1336
rect 4454 1268 4512 1302
rect 4454 1234 4466 1268
rect 4500 1234 4512 1268
rect 4454 1200 4512 1234
rect 4454 1166 4466 1200
rect 4500 1166 4512 1200
rect 4454 1132 4512 1166
rect 4454 1098 4466 1132
rect 4500 1098 4512 1132
rect 4454 1064 4512 1098
rect 4454 1030 4466 1064
rect 4500 1030 4512 1064
rect 4454 996 4512 1030
rect 4454 962 4466 996
rect 4500 962 4512 996
rect 4454 928 4512 962
rect 4454 894 4466 928
rect 4500 894 4512 928
rect 4454 860 4512 894
rect 4454 826 4466 860
rect 4500 826 4512 860
rect 4454 792 4512 826
rect 4454 758 4466 792
rect 4500 758 4512 792
rect 4454 724 4512 758
rect 4454 690 4466 724
rect 4500 690 4512 724
rect 4454 656 4512 690
rect 4454 622 4466 656
rect 4500 622 4512 656
rect 4454 591 4512 622
rect 4542 2560 4600 2591
rect 4542 2526 4554 2560
rect 4588 2526 4600 2560
rect 4542 2492 4600 2526
rect 4542 2458 4554 2492
rect 4588 2458 4600 2492
rect 4542 2424 4600 2458
rect 4542 2390 4554 2424
rect 4588 2390 4600 2424
rect 4542 2356 4600 2390
rect 4542 2322 4554 2356
rect 4588 2322 4600 2356
rect 4542 2288 4600 2322
rect 4542 2254 4554 2288
rect 4588 2254 4600 2288
rect 4542 2220 4600 2254
rect 4542 2186 4554 2220
rect 4588 2186 4600 2220
rect 4542 2152 4600 2186
rect 4542 2118 4554 2152
rect 4588 2118 4600 2152
rect 4542 2084 4600 2118
rect 4542 2050 4554 2084
rect 4588 2050 4600 2084
rect 4542 2016 4600 2050
rect 4542 1982 4554 2016
rect 4588 1982 4600 2016
rect 4542 1948 4600 1982
rect 4542 1914 4554 1948
rect 4588 1914 4600 1948
rect 4542 1880 4600 1914
rect 4542 1846 4554 1880
rect 4588 1846 4600 1880
rect 4542 1812 4600 1846
rect 4542 1778 4554 1812
rect 4588 1778 4600 1812
rect 4542 1744 4600 1778
rect 4542 1710 4554 1744
rect 4588 1710 4600 1744
rect 4542 1676 4600 1710
rect 4542 1642 4554 1676
rect 4588 1642 4600 1676
rect 4542 1608 4600 1642
rect 4542 1574 4554 1608
rect 4588 1574 4600 1608
rect 4542 1540 4600 1574
rect 4542 1506 4554 1540
rect 4588 1506 4600 1540
rect 4542 1472 4600 1506
rect 4542 1438 4554 1472
rect 4588 1438 4600 1472
rect 4542 1404 4600 1438
rect 4542 1370 4554 1404
rect 4588 1370 4600 1404
rect 4542 1336 4600 1370
rect 4542 1302 4554 1336
rect 4588 1302 4600 1336
rect 4542 1268 4600 1302
rect 4542 1234 4554 1268
rect 4588 1234 4600 1268
rect 4542 1200 4600 1234
rect 4542 1166 4554 1200
rect 4588 1166 4600 1200
rect 4542 1132 4600 1166
rect 4542 1098 4554 1132
rect 4588 1098 4600 1132
rect 4542 1064 4600 1098
rect 4542 1030 4554 1064
rect 4588 1030 4600 1064
rect 4542 996 4600 1030
rect 4542 962 4554 996
rect 4588 962 4600 996
rect 4542 928 4600 962
rect 4542 894 4554 928
rect 4588 894 4600 928
rect 4542 860 4600 894
rect 4542 826 4554 860
rect 4588 826 4600 860
rect 4542 792 4600 826
rect 4542 758 4554 792
rect 4588 758 4600 792
rect 4542 724 4600 758
rect 4542 690 4554 724
rect 4588 690 4600 724
rect 4542 656 4600 690
rect 4542 622 4554 656
rect 4588 622 4600 656
rect 4542 591 4600 622
rect 4630 2560 4688 2591
rect 4630 2526 4642 2560
rect 4676 2526 4688 2560
rect 4630 2492 4688 2526
rect 4630 2458 4642 2492
rect 4676 2458 4688 2492
rect 4630 2424 4688 2458
rect 4630 2390 4642 2424
rect 4676 2390 4688 2424
rect 4630 2356 4688 2390
rect 4630 2322 4642 2356
rect 4676 2322 4688 2356
rect 4630 2288 4688 2322
rect 4630 2254 4642 2288
rect 4676 2254 4688 2288
rect 4630 2220 4688 2254
rect 4630 2186 4642 2220
rect 4676 2186 4688 2220
rect 4630 2152 4688 2186
rect 4630 2118 4642 2152
rect 4676 2118 4688 2152
rect 4630 2084 4688 2118
rect 4630 2050 4642 2084
rect 4676 2050 4688 2084
rect 4630 2016 4688 2050
rect 4630 1982 4642 2016
rect 4676 1982 4688 2016
rect 4630 1948 4688 1982
rect 4630 1914 4642 1948
rect 4676 1914 4688 1948
rect 4630 1880 4688 1914
rect 4630 1846 4642 1880
rect 4676 1846 4688 1880
rect 4630 1812 4688 1846
rect 4630 1778 4642 1812
rect 4676 1778 4688 1812
rect 4630 1744 4688 1778
rect 4630 1710 4642 1744
rect 4676 1710 4688 1744
rect 4630 1676 4688 1710
rect 4630 1642 4642 1676
rect 4676 1642 4688 1676
rect 4630 1608 4688 1642
rect 4630 1574 4642 1608
rect 4676 1574 4688 1608
rect 4630 1540 4688 1574
rect 4630 1506 4642 1540
rect 4676 1506 4688 1540
rect 4630 1472 4688 1506
rect 4630 1438 4642 1472
rect 4676 1438 4688 1472
rect 4630 1404 4688 1438
rect 4630 1370 4642 1404
rect 4676 1370 4688 1404
rect 4630 1336 4688 1370
rect 4630 1302 4642 1336
rect 4676 1302 4688 1336
rect 4630 1268 4688 1302
rect 4630 1234 4642 1268
rect 4676 1234 4688 1268
rect 4630 1200 4688 1234
rect 4630 1166 4642 1200
rect 4676 1166 4688 1200
rect 4630 1132 4688 1166
rect 4630 1098 4642 1132
rect 4676 1098 4688 1132
rect 4630 1064 4688 1098
rect 4630 1030 4642 1064
rect 4676 1030 4688 1064
rect 4630 996 4688 1030
rect 4630 962 4642 996
rect 4676 962 4688 996
rect 4630 928 4688 962
rect 4630 894 4642 928
rect 4676 894 4688 928
rect 4630 860 4688 894
rect 4630 826 4642 860
rect 4676 826 4688 860
rect 4630 792 4688 826
rect 4630 758 4642 792
rect 4676 758 4688 792
rect 4630 724 4688 758
rect 4630 690 4642 724
rect 4676 690 4688 724
rect 4630 656 4688 690
rect 4630 622 4642 656
rect 4676 622 4688 656
rect 4630 591 4688 622
rect 4718 2560 4776 2591
rect 4718 2526 4730 2560
rect 4764 2526 4776 2560
rect 4718 2492 4776 2526
rect 4718 2458 4730 2492
rect 4764 2458 4776 2492
rect 4718 2424 4776 2458
rect 4718 2390 4730 2424
rect 4764 2390 4776 2424
rect 4718 2356 4776 2390
rect 4718 2322 4730 2356
rect 4764 2322 4776 2356
rect 4718 2288 4776 2322
rect 4718 2254 4730 2288
rect 4764 2254 4776 2288
rect 4718 2220 4776 2254
rect 4718 2186 4730 2220
rect 4764 2186 4776 2220
rect 4718 2152 4776 2186
rect 4718 2118 4730 2152
rect 4764 2118 4776 2152
rect 4718 2084 4776 2118
rect 4718 2050 4730 2084
rect 4764 2050 4776 2084
rect 4718 2016 4776 2050
rect 4718 1982 4730 2016
rect 4764 1982 4776 2016
rect 4718 1948 4776 1982
rect 4718 1914 4730 1948
rect 4764 1914 4776 1948
rect 4718 1880 4776 1914
rect 4718 1846 4730 1880
rect 4764 1846 4776 1880
rect 4718 1812 4776 1846
rect 4718 1778 4730 1812
rect 4764 1778 4776 1812
rect 4718 1744 4776 1778
rect 4718 1710 4730 1744
rect 4764 1710 4776 1744
rect 4718 1676 4776 1710
rect 4718 1642 4730 1676
rect 4764 1642 4776 1676
rect 4718 1608 4776 1642
rect 4718 1574 4730 1608
rect 4764 1574 4776 1608
rect 4718 1540 4776 1574
rect 4718 1506 4730 1540
rect 4764 1506 4776 1540
rect 4718 1472 4776 1506
rect 4718 1438 4730 1472
rect 4764 1438 4776 1472
rect 4718 1404 4776 1438
rect 4718 1370 4730 1404
rect 4764 1370 4776 1404
rect 4718 1336 4776 1370
rect 4718 1302 4730 1336
rect 4764 1302 4776 1336
rect 4718 1268 4776 1302
rect 4718 1234 4730 1268
rect 4764 1234 4776 1268
rect 4718 1200 4776 1234
rect 4718 1166 4730 1200
rect 4764 1166 4776 1200
rect 4718 1132 4776 1166
rect 4718 1098 4730 1132
rect 4764 1098 4776 1132
rect 4718 1064 4776 1098
rect 4718 1030 4730 1064
rect 4764 1030 4776 1064
rect 4718 996 4776 1030
rect 4718 962 4730 996
rect 4764 962 4776 996
rect 4718 928 4776 962
rect 4718 894 4730 928
rect 4764 894 4776 928
rect 4718 860 4776 894
rect 4718 826 4730 860
rect 4764 826 4776 860
rect 4718 792 4776 826
rect 4718 758 4730 792
rect 4764 758 4776 792
rect 4718 724 4776 758
rect 4718 690 4730 724
rect 4764 690 4776 724
rect 4718 656 4776 690
rect 4718 622 4730 656
rect 4764 622 4776 656
rect 4718 591 4776 622
rect 4806 2560 4864 2591
rect 4806 2526 4818 2560
rect 4852 2526 4864 2560
rect 4806 2492 4864 2526
rect 4806 2458 4818 2492
rect 4852 2458 4864 2492
rect 4806 2424 4864 2458
rect 4806 2390 4818 2424
rect 4852 2390 4864 2424
rect 4806 2356 4864 2390
rect 4806 2322 4818 2356
rect 4852 2322 4864 2356
rect 4806 2288 4864 2322
rect 4806 2254 4818 2288
rect 4852 2254 4864 2288
rect 4806 2220 4864 2254
rect 4806 2186 4818 2220
rect 4852 2186 4864 2220
rect 4806 2152 4864 2186
rect 4806 2118 4818 2152
rect 4852 2118 4864 2152
rect 4806 2084 4864 2118
rect 4806 2050 4818 2084
rect 4852 2050 4864 2084
rect 4806 2016 4864 2050
rect 4806 1982 4818 2016
rect 4852 1982 4864 2016
rect 4806 1948 4864 1982
rect 4806 1914 4818 1948
rect 4852 1914 4864 1948
rect 4806 1880 4864 1914
rect 4806 1846 4818 1880
rect 4852 1846 4864 1880
rect 4806 1812 4864 1846
rect 4806 1778 4818 1812
rect 4852 1778 4864 1812
rect 4806 1744 4864 1778
rect 4806 1710 4818 1744
rect 4852 1710 4864 1744
rect 4806 1676 4864 1710
rect 4806 1642 4818 1676
rect 4852 1642 4864 1676
rect 4806 1608 4864 1642
rect 4806 1574 4818 1608
rect 4852 1574 4864 1608
rect 4806 1540 4864 1574
rect 4806 1506 4818 1540
rect 4852 1506 4864 1540
rect 4806 1472 4864 1506
rect 4806 1438 4818 1472
rect 4852 1438 4864 1472
rect 4806 1404 4864 1438
rect 4806 1370 4818 1404
rect 4852 1370 4864 1404
rect 4806 1336 4864 1370
rect 4806 1302 4818 1336
rect 4852 1302 4864 1336
rect 4806 1268 4864 1302
rect 4806 1234 4818 1268
rect 4852 1234 4864 1268
rect 4806 1200 4864 1234
rect 4806 1166 4818 1200
rect 4852 1166 4864 1200
rect 4806 1132 4864 1166
rect 4806 1098 4818 1132
rect 4852 1098 4864 1132
rect 4806 1064 4864 1098
rect 4806 1030 4818 1064
rect 4852 1030 4864 1064
rect 4806 996 4864 1030
rect 4806 962 4818 996
rect 4852 962 4864 996
rect 4806 928 4864 962
rect 4806 894 4818 928
rect 4852 894 4864 928
rect 4806 860 4864 894
rect 4806 826 4818 860
rect 4852 826 4864 860
rect 4806 792 4864 826
rect 4806 758 4818 792
rect 4852 758 4864 792
rect 4806 724 4864 758
rect 4806 690 4818 724
rect 4852 690 4864 724
rect 4806 656 4864 690
rect 4806 622 4818 656
rect 4852 622 4864 656
rect 4806 591 4864 622
rect 4894 2560 4952 2591
rect 4894 2526 4906 2560
rect 4940 2526 4952 2560
rect 4894 2492 4952 2526
rect 4894 2458 4906 2492
rect 4940 2458 4952 2492
rect 4894 2424 4952 2458
rect 4894 2390 4906 2424
rect 4940 2390 4952 2424
rect 4894 2356 4952 2390
rect 4894 2322 4906 2356
rect 4940 2322 4952 2356
rect 4894 2288 4952 2322
rect 4894 2254 4906 2288
rect 4940 2254 4952 2288
rect 4894 2220 4952 2254
rect 4894 2186 4906 2220
rect 4940 2186 4952 2220
rect 4894 2152 4952 2186
rect 4894 2118 4906 2152
rect 4940 2118 4952 2152
rect 4894 2084 4952 2118
rect 4894 2050 4906 2084
rect 4940 2050 4952 2084
rect 4894 2016 4952 2050
rect 4894 1982 4906 2016
rect 4940 1982 4952 2016
rect 4894 1948 4952 1982
rect 4894 1914 4906 1948
rect 4940 1914 4952 1948
rect 4894 1880 4952 1914
rect 4894 1846 4906 1880
rect 4940 1846 4952 1880
rect 4894 1812 4952 1846
rect 4894 1778 4906 1812
rect 4940 1778 4952 1812
rect 4894 1744 4952 1778
rect 4894 1710 4906 1744
rect 4940 1710 4952 1744
rect 4894 1676 4952 1710
rect 4894 1642 4906 1676
rect 4940 1642 4952 1676
rect 4894 1608 4952 1642
rect 4894 1574 4906 1608
rect 4940 1574 4952 1608
rect 4894 1540 4952 1574
rect 4894 1506 4906 1540
rect 4940 1506 4952 1540
rect 4894 1472 4952 1506
rect 4894 1438 4906 1472
rect 4940 1438 4952 1472
rect 4894 1404 4952 1438
rect 4894 1370 4906 1404
rect 4940 1370 4952 1404
rect 4894 1336 4952 1370
rect 4894 1302 4906 1336
rect 4940 1302 4952 1336
rect 4894 1268 4952 1302
rect 4894 1234 4906 1268
rect 4940 1234 4952 1268
rect 4894 1200 4952 1234
rect 4894 1166 4906 1200
rect 4940 1166 4952 1200
rect 4894 1132 4952 1166
rect 4894 1098 4906 1132
rect 4940 1098 4952 1132
rect 4894 1064 4952 1098
rect 4894 1030 4906 1064
rect 4940 1030 4952 1064
rect 4894 996 4952 1030
rect 4894 962 4906 996
rect 4940 962 4952 996
rect 4894 928 4952 962
rect 4894 894 4906 928
rect 4940 894 4952 928
rect 4894 860 4952 894
rect 4894 826 4906 860
rect 4940 826 4952 860
rect 4894 792 4952 826
rect 4894 758 4906 792
rect 4940 758 4952 792
rect 4894 724 4952 758
rect 4894 690 4906 724
rect 4940 690 4952 724
rect 4894 656 4952 690
rect 4894 622 4906 656
rect 4940 622 4952 656
rect 4894 591 4952 622
rect 4982 2560 5040 2591
rect 4982 2526 4994 2560
rect 5028 2526 5040 2560
rect 4982 2492 5040 2526
rect 4982 2458 4994 2492
rect 5028 2458 5040 2492
rect 4982 2424 5040 2458
rect 4982 2390 4994 2424
rect 5028 2390 5040 2424
rect 4982 2356 5040 2390
rect 4982 2322 4994 2356
rect 5028 2322 5040 2356
rect 4982 2288 5040 2322
rect 4982 2254 4994 2288
rect 5028 2254 5040 2288
rect 4982 2220 5040 2254
rect 4982 2186 4994 2220
rect 5028 2186 5040 2220
rect 4982 2152 5040 2186
rect 4982 2118 4994 2152
rect 5028 2118 5040 2152
rect 4982 2084 5040 2118
rect 4982 2050 4994 2084
rect 5028 2050 5040 2084
rect 4982 2016 5040 2050
rect 4982 1982 4994 2016
rect 5028 1982 5040 2016
rect 4982 1948 5040 1982
rect 4982 1914 4994 1948
rect 5028 1914 5040 1948
rect 4982 1880 5040 1914
rect 4982 1846 4994 1880
rect 5028 1846 5040 1880
rect 4982 1812 5040 1846
rect 4982 1778 4994 1812
rect 5028 1778 5040 1812
rect 4982 1744 5040 1778
rect 4982 1710 4994 1744
rect 5028 1710 5040 1744
rect 4982 1676 5040 1710
rect 4982 1642 4994 1676
rect 5028 1642 5040 1676
rect 4982 1608 5040 1642
rect 4982 1574 4994 1608
rect 5028 1574 5040 1608
rect 4982 1540 5040 1574
rect 4982 1506 4994 1540
rect 5028 1506 5040 1540
rect 4982 1472 5040 1506
rect 4982 1438 4994 1472
rect 5028 1438 5040 1472
rect 4982 1404 5040 1438
rect 4982 1370 4994 1404
rect 5028 1370 5040 1404
rect 4982 1336 5040 1370
rect 4982 1302 4994 1336
rect 5028 1302 5040 1336
rect 4982 1268 5040 1302
rect 4982 1234 4994 1268
rect 5028 1234 5040 1268
rect 4982 1200 5040 1234
rect 4982 1166 4994 1200
rect 5028 1166 5040 1200
rect 4982 1132 5040 1166
rect 4982 1098 4994 1132
rect 5028 1098 5040 1132
rect 4982 1064 5040 1098
rect 4982 1030 4994 1064
rect 5028 1030 5040 1064
rect 4982 996 5040 1030
rect 4982 962 4994 996
rect 5028 962 5040 996
rect 4982 928 5040 962
rect 4982 894 4994 928
rect 5028 894 5040 928
rect 4982 860 5040 894
rect 4982 826 4994 860
rect 5028 826 5040 860
rect 4982 792 5040 826
rect 4982 758 4994 792
rect 5028 758 5040 792
rect 4982 724 5040 758
rect 4982 690 4994 724
rect 5028 690 5040 724
rect 4982 656 5040 690
rect 4982 622 4994 656
rect 5028 622 5040 656
rect 4982 591 5040 622
rect 5070 2560 5128 2591
rect 5070 2526 5082 2560
rect 5116 2526 5128 2560
rect 5070 2492 5128 2526
rect 5070 2458 5082 2492
rect 5116 2458 5128 2492
rect 5070 2424 5128 2458
rect 5070 2390 5082 2424
rect 5116 2390 5128 2424
rect 5070 2356 5128 2390
rect 5070 2322 5082 2356
rect 5116 2322 5128 2356
rect 5070 2288 5128 2322
rect 5070 2254 5082 2288
rect 5116 2254 5128 2288
rect 5070 2220 5128 2254
rect 5070 2186 5082 2220
rect 5116 2186 5128 2220
rect 5070 2152 5128 2186
rect 5070 2118 5082 2152
rect 5116 2118 5128 2152
rect 5070 2084 5128 2118
rect 5070 2050 5082 2084
rect 5116 2050 5128 2084
rect 5070 2016 5128 2050
rect 5070 1982 5082 2016
rect 5116 1982 5128 2016
rect 5070 1948 5128 1982
rect 5070 1914 5082 1948
rect 5116 1914 5128 1948
rect 5070 1880 5128 1914
rect 5070 1846 5082 1880
rect 5116 1846 5128 1880
rect 5070 1812 5128 1846
rect 5070 1778 5082 1812
rect 5116 1778 5128 1812
rect 5070 1744 5128 1778
rect 5070 1710 5082 1744
rect 5116 1710 5128 1744
rect 5070 1676 5128 1710
rect 5070 1642 5082 1676
rect 5116 1642 5128 1676
rect 5070 1608 5128 1642
rect 5070 1574 5082 1608
rect 5116 1574 5128 1608
rect 5070 1540 5128 1574
rect 5070 1506 5082 1540
rect 5116 1506 5128 1540
rect 5070 1472 5128 1506
rect 5070 1438 5082 1472
rect 5116 1438 5128 1472
rect 5070 1404 5128 1438
rect 5070 1370 5082 1404
rect 5116 1370 5128 1404
rect 5070 1336 5128 1370
rect 5070 1302 5082 1336
rect 5116 1302 5128 1336
rect 5070 1268 5128 1302
rect 5070 1234 5082 1268
rect 5116 1234 5128 1268
rect 5070 1200 5128 1234
rect 5070 1166 5082 1200
rect 5116 1166 5128 1200
rect 5070 1132 5128 1166
rect 5070 1098 5082 1132
rect 5116 1098 5128 1132
rect 5070 1064 5128 1098
rect 5070 1030 5082 1064
rect 5116 1030 5128 1064
rect 5070 996 5128 1030
rect 5070 962 5082 996
rect 5116 962 5128 996
rect 5070 928 5128 962
rect 5070 894 5082 928
rect 5116 894 5128 928
rect 5070 860 5128 894
rect 5070 826 5082 860
rect 5116 826 5128 860
rect 5070 792 5128 826
rect 5070 758 5082 792
rect 5116 758 5128 792
rect 5070 724 5128 758
rect 5070 690 5082 724
rect 5116 690 5128 724
rect 5070 656 5128 690
rect 5070 622 5082 656
rect 5116 622 5128 656
rect 5070 591 5128 622
rect 5158 2560 5216 2591
rect 5158 2526 5170 2560
rect 5204 2526 5216 2560
rect 5158 2492 5216 2526
rect 5158 2458 5170 2492
rect 5204 2458 5216 2492
rect 5158 2424 5216 2458
rect 5158 2390 5170 2424
rect 5204 2390 5216 2424
rect 5158 2356 5216 2390
rect 5158 2322 5170 2356
rect 5204 2322 5216 2356
rect 5158 2288 5216 2322
rect 5158 2254 5170 2288
rect 5204 2254 5216 2288
rect 5158 2220 5216 2254
rect 5158 2186 5170 2220
rect 5204 2186 5216 2220
rect 5158 2152 5216 2186
rect 5158 2118 5170 2152
rect 5204 2118 5216 2152
rect 5158 2084 5216 2118
rect 5158 2050 5170 2084
rect 5204 2050 5216 2084
rect 5158 2016 5216 2050
rect 5158 1982 5170 2016
rect 5204 1982 5216 2016
rect 5158 1948 5216 1982
rect 5158 1914 5170 1948
rect 5204 1914 5216 1948
rect 5158 1880 5216 1914
rect 5158 1846 5170 1880
rect 5204 1846 5216 1880
rect 5158 1812 5216 1846
rect 5158 1778 5170 1812
rect 5204 1778 5216 1812
rect 5158 1744 5216 1778
rect 5158 1710 5170 1744
rect 5204 1710 5216 1744
rect 5158 1676 5216 1710
rect 5158 1642 5170 1676
rect 5204 1642 5216 1676
rect 5158 1608 5216 1642
rect 5158 1574 5170 1608
rect 5204 1574 5216 1608
rect 5158 1540 5216 1574
rect 5158 1506 5170 1540
rect 5204 1506 5216 1540
rect 5158 1472 5216 1506
rect 5158 1438 5170 1472
rect 5204 1438 5216 1472
rect 5158 1404 5216 1438
rect 5158 1370 5170 1404
rect 5204 1370 5216 1404
rect 5158 1336 5216 1370
rect 5158 1302 5170 1336
rect 5204 1302 5216 1336
rect 5158 1268 5216 1302
rect 5158 1234 5170 1268
rect 5204 1234 5216 1268
rect 5158 1200 5216 1234
rect 5158 1166 5170 1200
rect 5204 1166 5216 1200
rect 5158 1132 5216 1166
rect 5158 1098 5170 1132
rect 5204 1098 5216 1132
rect 5158 1064 5216 1098
rect 5158 1030 5170 1064
rect 5204 1030 5216 1064
rect 5158 996 5216 1030
rect 5158 962 5170 996
rect 5204 962 5216 996
rect 5158 928 5216 962
rect 5158 894 5170 928
rect 5204 894 5216 928
rect 5158 860 5216 894
rect 5158 826 5170 860
rect 5204 826 5216 860
rect 5158 792 5216 826
rect 5158 758 5170 792
rect 5204 758 5216 792
rect 5158 724 5216 758
rect 5158 690 5170 724
rect 5204 690 5216 724
rect 5158 656 5216 690
rect 5158 622 5170 656
rect 5204 622 5216 656
rect 5158 591 5216 622
rect 5246 2560 5304 2591
rect 5246 2526 5258 2560
rect 5292 2526 5304 2560
rect 5246 2492 5304 2526
rect 5246 2458 5258 2492
rect 5292 2458 5304 2492
rect 5246 2424 5304 2458
rect 5246 2390 5258 2424
rect 5292 2390 5304 2424
rect 5246 2356 5304 2390
rect 5246 2322 5258 2356
rect 5292 2322 5304 2356
rect 5246 2288 5304 2322
rect 5246 2254 5258 2288
rect 5292 2254 5304 2288
rect 5246 2220 5304 2254
rect 5246 2186 5258 2220
rect 5292 2186 5304 2220
rect 5246 2152 5304 2186
rect 5246 2118 5258 2152
rect 5292 2118 5304 2152
rect 5246 2084 5304 2118
rect 5246 2050 5258 2084
rect 5292 2050 5304 2084
rect 5246 2016 5304 2050
rect 5246 1982 5258 2016
rect 5292 1982 5304 2016
rect 5246 1948 5304 1982
rect 5246 1914 5258 1948
rect 5292 1914 5304 1948
rect 5246 1880 5304 1914
rect 5246 1846 5258 1880
rect 5292 1846 5304 1880
rect 5246 1812 5304 1846
rect 5246 1778 5258 1812
rect 5292 1778 5304 1812
rect 5246 1744 5304 1778
rect 5246 1710 5258 1744
rect 5292 1710 5304 1744
rect 5246 1676 5304 1710
rect 5246 1642 5258 1676
rect 5292 1642 5304 1676
rect 5246 1608 5304 1642
rect 5246 1574 5258 1608
rect 5292 1574 5304 1608
rect 5246 1540 5304 1574
rect 5246 1506 5258 1540
rect 5292 1506 5304 1540
rect 5246 1472 5304 1506
rect 5246 1438 5258 1472
rect 5292 1438 5304 1472
rect 5246 1404 5304 1438
rect 5246 1370 5258 1404
rect 5292 1370 5304 1404
rect 5246 1336 5304 1370
rect 5246 1302 5258 1336
rect 5292 1302 5304 1336
rect 5246 1268 5304 1302
rect 5246 1234 5258 1268
rect 5292 1234 5304 1268
rect 5246 1200 5304 1234
rect 5246 1166 5258 1200
rect 5292 1166 5304 1200
rect 5246 1132 5304 1166
rect 5246 1098 5258 1132
rect 5292 1098 5304 1132
rect 5246 1064 5304 1098
rect 5246 1030 5258 1064
rect 5292 1030 5304 1064
rect 5246 996 5304 1030
rect 5246 962 5258 996
rect 5292 962 5304 996
rect 5246 928 5304 962
rect 5246 894 5258 928
rect 5292 894 5304 928
rect 5246 860 5304 894
rect 5246 826 5258 860
rect 5292 826 5304 860
rect 5246 792 5304 826
rect 5246 758 5258 792
rect 5292 758 5304 792
rect 5246 724 5304 758
rect 5246 690 5258 724
rect 5292 690 5304 724
rect 5246 656 5304 690
rect 5246 622 5258 656
rect 5292 622 5304 656
rect 5246 591 5304 622
<< pdiffc >>
rect 4290 2526 4324 2560
rect 4290 2458 4324 2492
rect 4290 2390 4324 2424
rect 4290 2322 4324 2356
rect 4290 2254 4324 2288
rect 4290 2186 4324 2220
rect 4290 2118 4324 2152
rect 4290 2050 4324 2084
rect 4290 1982 4324 2016
rect 4290 1914 4324 1948
rect 4290 1846 4324 1880
rect 4290 1778 4324 1812
rect 4290 1710 4324 1744
rect 4290 1642 4324 1676
rect 4290 1574 4324 1608
rect 4290 1506 4324 1540
rect 4290 1438 4324 1472
rect 4290 1370 4324 1404
rect 4290 1302 4324 1336
rect 4290 1234 4324 1268
rect 4290 1166 4324 1200
rect 4290 1098 4324 1132
rect 4290 1030 4324 1064
rect 4290 962 4324 996
rect 4290 894 4324 928
rect 4290 826 4324 860
rect 4290 758 4324 792
rect 4290 690 4324 724
rect 4290 622 4324 656
rect 4378 2526 4412 2560
rect 4378 2458 4412 2492
rect 4378 2390 4412 2424
rect 4378 2322 4412 2356
rect 4378 2254 4412 2288
rect 4378 2186 4412 2220
rect 4378 2118 4412 2152
rect 4378 2050 4412 2084
rect 4378 1982 4412 2016
rect 4378 1914 4412 1948
rect 4378 1846 4412 1880
rect 4378 1778 4412 1812
rect 4378 1710 4412 1744
rect 4378 1642 4412 1676
rect 4378 1574 4412 1608
rect 4378 1506 4412 1540
rect 4378 1438 4412 1472
rect 4378 1370 4412 1404
rect 4378 1302 4412 1336
rect 4378 1234 4412 1268
rect 4378 1166 4412 1200
rect 4378 1098 4412 1132
rect 4378 1030 4412 1064
rect 4378 962 4412 996
rect 4378 894 4412 928
rect 4378 826 4412 860
rect 4378 758 4412 792
rect 4378 690 4412 724
rect 4378 622 4412 656
rect 4466 2526 4500 2560
rect 4466 2458 4500 2492
rect 4466 2390 4500 2424
rect 4466 2322 4500 2356
rect 4466 2254 4500 2288
rect 4466 2186 4500 2220
rect 4466 2118 4500 2152
rect 4466 2050 4500 2084
rect 4466 1982 4500 2016
rect 4466 1914 4500 1948
rect 4466 1846 4500 1880
rect 4466 1778 4500 1812
rect 4466 1710 4500 1744
rect 4466 1642 4500 1676
rect 4466 1574 4500 1608
rect 4466 1506 4500 1540
rect 4466 1438 4500 1472
rect 4466 1370 4500 1404
rect 4466 1302 4500 1336
rect 4466 1234 4500 1268
rect 4466 1166 4500 1200
rect 4466 1098 4500 1132
rect 4466 1030 4500 1064
rect 4466 962 4500 996
rect 4466 894 4500 928
rect 4466 826 4500 860
rect 4466 758 4500 792
rect 4466 690 4500 724
rect 4466 622 4500 656
rect 4554 2526 4588 2560
rect 4554 2458 4588 2492
rect 4554 2390 4588 2424
rect 4554 2322 4588 2356
rect 4554 2254 4588 2288
rect 4554 2186 4588 2220
rect 4554 2118 4588 2152
rect 4554 2050 4588 2084
rect 4554 1982 4588 2016
rect 4554 1914 4588 1948
rect 4554 1846 4588 1880
rect 4554 1778 4588 1812
rect 4554 1710 4588 1744
rect 4554 1642 4588 1676
rect 4554 1574 4588 1608
rect 4554 1506 4588 1540
rect 4554 1438 4588 1472
rect 4554 1370 4588 1404
rect 4554 1302 4588 1336
rect 4554 1234 4588 1268
rect 4554 1166 4588 1200
rect 4554 1098 4588 1132
rect 4554 1030 4588 1064
rect 4554 962 4588 996
rect 4554 894 4588 928
rect 4554 826 4588 860
rect 4554 758 4588 792
rect 4554 690 4588 724
rect 4554 622 4588 656
rect 4642 2526 4676 2560
rect 4642 2458 4676 2492
rect 4642 2390 4676 2424
rect 4642 2322 4676 2356
rect 4642 2254 4676 2288
rect 4642 2186 4676 2220
rect 4642 2118 4676 2152
rect 4642 2050 4676 2084
rect 4642 1982 4676 2016
rect 4642 1914 4676 1948
rect 4642 1846 4676 1880
rect 4642 1778 4676 1812
rect 4642 1710 4676 1744
rect 4642 1642 4676 1676
rect 4642 1574 4676 1608
rect 4642 1506 4676 1540
rect 4642 1438 4676 1472
rect 4642 1370 4676 1404
rect 4642 1302 4676 1336
rect 4642 1234 4676 1268
rect 4642 1166 4676 1200
rect 4642 1098 4676 1132
rect 4642 1030 4676 1064
rect 4642 962 4676 996
rect 4642 894 4676 928
rect 4642 826 4676 860
rect 4642 758 4676 792
rect 4642 690 4676 724
rect 4642 622 4676 656
rect 4730 2526 4764 2560
rect 4730 2458 4764 2492
rect 4730 2390 4764 2424
rect 4730 2322 4764 2356
rect 4730 2254 4764 2288
rect 4730 2186 4764 2220
rect 4730 2118 4764 2152
rect 4730 2050 4764 2084
rect 4730 1982 4764 2016
rect 4730 1914 4764 1948
rect 4730 1846 4764 1880
rect 4730 1778 4764 1812
rect 4730 1710 4764 1744
rect 4730 1642 4764 1676
rect 4730 1574 4764 1608
rect 4730 1506 4764 1540
rect 4730 1438 4764 1472
rect 4730 1370 4764 1404
rect 4730 1302 4764 1336
rect 4730 1234 4764 1268
rect 4730 1166 4764 1200
rect 4730 1098 4764 1132
rect 4730 1030 4764 1064
rect 4730 962 4764 996
rect 4730 894 4764 928
rect 4730 826 4764 860
rect 4730 758 4764 792
rect 4730 690 4764 724
rect 4730 622 4764 656
rect 4818 2526 4852 2560
rect 4818 2458 4852 2492
rect 4818 2390 4852 2424
rect 4818 2322 4852 2356
rect 4818 2254 4852 2288
rect 4818 2186 4852 2220
rect 4818 2118 4852 2152
rect 4818 2050 4852 2084
rect 4818 1982 4852 2016
rect 4818 1914 4852 1948
rect 4818 1846 4852 1880
rect 4818 1778 4852 1812
rect 4818 1710 4852 1744
rect 4818 1642 4852 1676
rect 4818 1574 4852 1608
rect 4818 1506 4852 1540
rect 4818 1438 4852 1472
rect 4818 1370 4852 1404
rect 4818 1302 4852 1336
rect 4818 1234 4852 1268
rect 4818 1166 4852 1200
rect 4818 1098 4852 1132
rect 4818 1030 4852 1064
rect 4818 962 4852 996
rect 4818 894 4852 928
rect 4818 826 4852 860
rect 4818 758 4852 792
rect 4818 690 4852 724
rect 4818 622 4852 656
rect 4906 2526 4940 2560
rect 4906 2458 4940 2492
rect 4906 2390 4940 2424
rect 4906 2322 4940 2356
rect 4906 2254 4940 2288
rect 4906 2186 4940 2220
rect 4906 2118 4940 2152
rect 4906 2050 4940 2084
rect 4906 1982 4940 2016
rect 4906 1914 4940 1948
rect 4906 1846 4940 1880
rect 4906 1778 4940 1812
rect 4906 1710 4940 1744
rect 4906 1642 4940 1676
rect 4906 1574 4940 1608
rect 4906 1506 4940 1540
rect 4906 1438 4940 1472
rect 4906 1370 4940 1404
rect 4906 1302 4940 1336
rect 4906 1234 4940 1268
rect 4906 1166 4940 1200
rect 4906 1098 4940 1132
rect 4906 1030 4940 1064
rect 4906 962 4940 996
rect 4906 894 4940 928
rect 4906 826 4940 860
rect 4906 758 4940 792
rect 4906 690 4940 724
rect 4906 622 4940 656
rect 4994 2526 5028 2560
rect 4994 2458 5028 2492
rect 4994 2390 5028 2424
rect 4994 2322 5028 2356
rect 4994 2254 5028 2288
rect 4994 2186 5028 2220
rect 4994 2118 5028 2152
rect 4994 2050 5028 2084
rect 4994 1982 5028 2016
rect 4994 1914 5028 1948
rect 4994 1846 5028 1880
rect 4994 1778 5028 1812
rect 4994 1710 5028 1744
rect 4994 1642 5028 1676
rect 4994 1574 5028 1608
rect 4994 1506 5028 1540
rect 4994 1438 5028 1472
rect 4994 1370 5028 1404
rect 4994 1302 5028 1336
rect 4994 1234 5028 1268
rect 4994 1166 5028 1200
rect 4994 1098 5028 1132
rect 4994 1030 5028 1064
rect 4994 962 5028 996
rect 4994 894 5028 928
rect 4994 826 5028 860
rect 4994 758 5028 792
rect 4994 690 5028 724
rect 4994 622 5028 656
rect 5082 2526 5116 2560
rect 5082 2458 5116 2492
rect 5082 2390 5116 2424
rect 5082 2322 5116 2356
rect 5082 2254 5116 2288
rect 5082 2186 5116 2220
rect 5082 2118 5116 2152
rect 5082 2050 5116 2084
rect 5082 1982 5116 2016
rect 5082 1914 5116 1948
rect 5082 1846 5116 1880
rect 5082 1778 5116 1812
rect 5082 1710 5116 1744
rect 5082 1642 5116 1676
rect 5082 1574 5116 1608
rect 5082 1506 5116 1540
rect 5082 1438 5116 1472
rect 5082 1370 5116 1404
rect 5082 1302 5116 1336
rect 5082 1234 5116 1268
rect 5082 1166 5116 1200
rect 5082 1098 5116 1132
rect 5082 1030 5116 1064
rect 5082 962 5116 996
rect 5082 894 5116 928
rect 5082 826 5116 860
rect 5082 758 5116 792
rect 5082 690 5116 724
rect 5082 622 5116 656
rect 5170 2526 5204 2560
rect 5170 2458 5204 2492
rect 5170 2390 5204 2424
rect 5170 2322 5204 2356
rect 5170 2254 5204 2288
rect 5170 2186 5204 2220
rect 5170 2118 5204 2152
rect 5170 2050 5204 2084
rect 5170 1982 5204 2016
rect 5170 1914 5204 1948
rect 5170 1846 5204 1880
rect 5170 1778 5204 1812
rect 5170 1710 5204 1744
rect 5170 1642 5204 1676
rect 5170 1574 5204 1608
rect 5170 1506 5204 1540
rect 5170 1438 5204 1472
rect 5170 1370 5204 1404
rect 5170 1302 5204 1336
rect 5170 1234 5204 1268
rect 5170 1166 5204 1200
rect 5170 1098 5204 1132
rect 5170 1030 5204 1064
rect 5170 962 5204 996
rect 5170 894 5204 928
rect 5170 826 5204 860
rect 5170 758 5204 792
rect 5170 690 5204 724
rect 5170 622 5204 656
rect 5258 2526 5292 2560
rect 5258 2458 5292 2492
rect 5258 2390 5292 2424
rect 5258 2322 5292 2356
rect 5258 2254 5292 2288
rect 5258 2186 5292 2220
rect 5258 2118 5292 2152
rect 5258 2050 5292 2084
rect 5258 1982 5292 2016
rect 5258 1914 5292 1948
rect 5258 1846 5292 1880
rect 5258 1778 5292 1812
rect 5258 1710 5292 1744
rect 5258 1642 5292 1676
rect 5258 1574 5292 1608
rect 5258 1506 5292 1540
rect 5258 1438 5292 1472
rect 5258 1370 5292 1404
rect 5258 1302 5292 1336
rect 5258 1234 5292 1268
rect 5258 1166 5292 1200
rect 5258 1098 5292 1132
rect 5258 1030 5292 1064
rect 5258 962 5292 996
rect 5258 894 5292 928
rect 5258 826 5292 860
rect 5258 758 5292 792
rect 5258 690 5292 724
rect 5258 622 5292 656
<< psubdiff >>
rect 3143 3388 3755 3458
<< nsubdiff >>
rect 4130 3004 5420 3005
rect 4130 2970 4364 3004
rect 4398 2970 4432 3004
rect 4466 2970 4500 3004
rect 4534 2970 4568 3004
rect 4602 2970 4636 3004
rect 4670 2970 4704 3004
rect 4738 2970 4772 3004
rect 4806 2970 4840 3004
rect 4874 2970 4908 3004
rect 4942 2970 4976 3004
rect 5010 2970 5044 3004
rect 5078 2970 5112 3004
rect 5146 2970 5180 3004
rect 5214 2970 5420 3004
rect 4130 2969 5420 2970
rect 4130 2559 4164 2969
rect 4130 2491 4164 2525
rect 4130 2423 4164 2457
rect 4130 2355 4164 2389
rect 4130 2287 4164 2321
rect 4130 2219 4164 2253
rect 4130 2151 4164 2185
rect 4130 2083 4164 2117
rect 4130 2015 4164 2049
rect 4130 1947 4164 1981
rect 4130 1879 4164 1913
rect 4130 1811 4164 1845
rect 4130 1743 4164 1777
rect 4130 1675 4164 1709
rect 4130 1607 4164 1641
rect 4130 1539 4164 1573
rect 4130 1471 4164 1505
rect 4130 1403 4164 1437
rect 4130 1335 4164 1369
rect 4130 1267 4164 1301
rect 4130 1199 4164 1233
rect 4130 1131 4164 1165
rect 4130 1063 4164 1097
rect 4130 995 4164 1029
rect 4130 927 4164 961
rect 4130 859 4164 893
rect 4130 791 4164 825
rect 4130 723 4164 757
rect 4130 655 4164 689
rect 4130 325 4164 621
rect 5386 2555 5420 2969
rect 5386 2487 5420 2521
rect 5386 2419 5420 2453
rect 5386 2351 5420 2385
rect 5386 2283 5420 2317
rect 5386 2215 5420 2249
rect 5386 2147 5420 2181
rect 5386 2079 5420 2113
rect 5386 2011 5420 2045
rect 5386 1943 5420 1977
rect 5386 1875 5420 1909
rect 5386 1807 5420 1841
rect 5386 1739 5420 1773
rect 5386 1671 5420 1705
rect 5386 1603 5420 1637
rect 5386 1535 5420 1569
rect 5386 1467 5420 1501
rect 5386 1399 5420 1433
rect 5386 1331 5420 1365
rect 5386 1263 5420 1297
rect 5386 1195 5420 1229
rect 5386 1127 5420 1161
rect 5386 1059 5420 1093
rect 5386 991 5420 1025
rect 5386 923 5420 957
rect 5386 855 5420 889
rect 5386 787 5420 821
rect 5386 719 5420 753
rect 5386 651 5420 685
rect 5386 325 5420 617
rect 4130 324 5420 325
rect 4130 290 4364 324
rect 4398 290 4432 324
rect 4466 290 4500 324
rect 4534 290 4568 324
rect 4602 290 4636 324
rect 4670 290 4704 324
rect 4738 290 4772 324
rect 4806 290 4840 324
rect 4874 290 4908 324
rect 4942 290 4976 324
rect 5010 290 5044 324
rect 5078 290 5112 324
rect 5146 290 5180 324
rect 5214 290 5420 324
rect 4130 289 5420 290
<< nsubdiffcont >>
rect 4364 2970 4398 3004
rect 4432 2970 4466 3004
rect 4500 2970 4534 3004
rect 4568 2970 4602 3004
rect 4636 2970 4670 3004
rect 4704 2970 4738 3004
rect 4772 2970 4806 3004
rect 4840 2970 4874 3004
rect 4908 2970 4942 3004
rect 4976 2970 5010 3004
rect 5044 2970 5078 3004
rect 5112 2970 5146 3004
rect 5180 2970 5214 3004
rect 4130 2525 4164 2559
rect 4130 2457 4164 2491
rect 4130 2389 4164 2423
rect 4130 2321 4164 2355
rect 4130 2253 4164 2287
rect 4130 2185 4164 2219
rect 4130 2117 4164 2151
rect 4130 2049 4164 2083
rect 4130 1981 4164 2015
rect 4130 1913 4164 1947
rect 4130 1845 4164 1879
rect 4130 1777 4164 1811
rect 4130 1709 4164 1743
rect 4130 1641 4164 1675
rect 4130 1573 4164 1607
rect 4130 1505 4164 1539
rect 4130 1437 4164 1471
rect 4130 1369 4164 1403
rect 4130 1301 4164 1335
rect 4130 1233 4164 1267
rect 4130 1165 4164 1199
rect 4130 1097 4164 1131
rect 4130 1029 4164 1063
rect 4130 961 4164 995
rect 4130 893 4164 927
rect 4130 825 4164 859
rect 4130 757 4164 791
rect 4130 689 4164 723
rect 4130 621 4164 655
rect 5386 2521 5420 2555
rect 5386 2453 5420 2487
rect 5386 2385 5420 2419
rect 5386 2317 5420 2351
rect 5386 2249 5420 2283
rect 5386 2181 5420 2215
rect 5386 2113 5420 2147
rect 5386 2045 5420 2079
rect 5386 1977 5420 2011
rect 5386 1909 5420 1943
rect 5386 1841 5420 1875
rect 5386 1773 5420 1807
rect 5386 1705 5420 1739
rect 5386 1637 5420 1671
rect 5386 1569 5420 1603
rect 5386 1501 5420 1535
rect 5386 1433 5420 1467
rect 5386 1365 5420 1399
rect 5386 1297 5420 1331
rect 5386 1229 5420 1263
rect 5386 1161 5420 1195
rect 5386 1093 5420 1127
rect 5386 1025 5420 1059
rect 5386 957 5420 991
rect 5386 889 5420 923
rect 5386 821 5420 855
rect 5386 753 5420 787
rect 5386 685 5420 719
rect 5386 617 5420 651
rect 4364 290 4398 324
rect 4432 290 4466 324
rect 4500 290 4534 324
rect 4568 290 4602 324
rect 4636 290 4670 324
rect 4704 290 4738 324
rect 4772 290 4806 324
rect 4840 290 4874 324
rect 4908 290 4942 324
rect 4976 290 5010 324
rect 5044 290 5078 324
rect 5112 290 5146 324
rect 5180 290 5214 324
<< poly >>
rect 4336 2591 4366 2617
rect 4424 2591 4454 2617
rect 4512 2591 4542 2617
rect 4600 2591 4630 2617
rect 4688 2591 4718 2617
rect 4776 2591 4806 2617
rect 4864 2591 4894 2617
rect 4952 2591 4982 2617
rect 5040 2591 5070 2617
rect 5128 2591 5158 2617
rect 5216 2591 5246 2617
rect 4336 553 4366 591
rect 4424 553 4454 591
rect 4336 524 4454 553
rect 4336 490 4378 524
rect 4412 490 4454 524
rect 4336 461 4454 490
rect 4512 553 4542 591
rect 4600 553 4630 591
rect 4512 524 4630 553
rect 4512 490 4554 524
rect 4588 490 4630 524
rect 4512 461 4630 490
rect 4688 553 4718 591
rect 4776 553 4806 591
rect 4688 524 4806 553
rect 4688 490 4730 524
rect 4764 490 4806 524
rect 4688 461 4806 490
rect 4864 553 4894 591
rect 4952 553 4982 591
rect 4864 524 4982 553
rect 4864 490 4906 524
rect 4940 490 4982 524
rect 4864 461 4982 490
rect 5040 553 5070 591
rect 5128 553 5158 591
rect 5216 553 5246 591
rect 5040 524 5246 553
rect 5040 490 5082 524
rect 5116 490 5246 524
rect 5040 461 5246 490
<< polycont >>
rect 4378 490 4412 524
rect 4554 490 4588 524
rect 4730 490 4764 524
rect 4906 490 4940 524
rect 5082 490 5116 524
<< locali >>
rect 680 3440 752 3458
rect 680 3406 699 3440
rect 733 3406 752 3440
rect 680 3010 752 3406
rect 280 2992 352 3010
rect 280 2958 299 2992
rect 333 2958 352 2992
rect 280 2940 352 2958
rect 392 2940 752 3010
rect 856 3440 928 3458
rect 856 3406 875 3440
rect 909 3406 928 3440
rect 856 2940 928 3406
rect 1032 3440 1104 3458
rect 1032 3406 1051 3440
rect 1085 3406 1104 3440
rect 1032 2940 1104 3406
rect 1208 3388 1280 3458
rect 1384 2940 1456 3458
rect 1560 3388 1632 3458
rect 1736 2940 1808 3458
rect 1912 3388 1984 3458
rect 2088 2940 2160 3458
rect 2264 3388 2336 3458
rect 2440 2940 2512 3458
rect 2616 3388 2688 3458
rect 2792 3440 2864 3458
rect 2792 3406 2811 3440
rect 2845 3406 2864 3440
rect 2792 2940 2864 3406
rect 2968 3440 3040 3458
rect 2968 3406 2987 3440
rect 3021 3406 3040 3440
rect 2968 2940 3040 3406
rect 3143 3440 3755 3458
rect 3143 3406 3163 3440
rect 3197 3406 3755 3440
rect 3143 3388 3755 3406
rect 3144 3010 3216 3388
rect 3144 2992 3740 3010
rect 3144 2958 3687 2992
rect 3721 2958 3740 2992
rect 3144 2940 3740 2958
rect 4130 3004 5420 3005
rect 4130 2970 4364 3004
rect 4398 2970 4432 3004
rect 4466 2970 4500 3004
rect 4534 2970 4568 3004
rect 4602 2970 4636 3004
rect 4670 2970 4704 3004
rect 4738 2970 4772 3004
rect 4806 2970 4840 3004
rect 4874 2970 4908 3004
rect 4942 2970 4976 3004
rect 5010 2970 5044 3004
rect 5078 2970 5112 3004
rect 5146 2970 5180 3004
rect 5214 2970 5420 3004
rect 4130 2969 5420 2970
rect 4130 2721 4164 2969
rect 4269 2877 5311 2906
rect 4269 2843 4290 2877
rect 4324 2843 4466 2877
rect 4500 2843 4642 2877
rect 4676 2843 4818 2877
rect 4852 2843 4994 2877
rect 5028 2843 5170 2877
rect 5204 2843 5311 2877
rect 4269 2807 5311 2843
rect 4269 2773 4378 2807
rect 4412 2773 4554 2807
rect 4588 2773 4730 2807
rect 4764 2773 4906 2807
rect 4940 2773 5082 2807
rect 5116 2773 5258 2807
rect 5292 2773 5311 2807
rect 4269 2755 5311 2773
rect 4130 2703 4343 2721
rect 4130 2702 4290 2703
rect 4130 2668 4149 2702
rect 4183 2669 4290 2702
rect 4324 2669 4343 2703
rect 4183 2668 4343 2669
rect 4130 2651 4343 2668
rect 4130 2650 4324 2651
rect 4130 2559 4164 2650
rect 4130 2491 4164 2525
rect 4130 2423 4164 2457
rect 4130 2355 4164 2389
rect 4130 2287 4164 2321
rect 4130 2219 4164 2253
rect 4130 2151 4164 2185
rect 4130 2083 4164 2117
rect 4130 2015 4164 2049
rect 4130 1947 4164 1981
rect 4130 1879 4164 1913
rect 4130 1811 4164 1845
rect 4130 1743 4164 1777
rect 4130 1675 4164 1709
rect 4130 1607 4164 1641
rect 4130 1539 4164 1573
rect 4130 1471 4164 1505
rect 4130 1403 4164 1437
rect 4130 1335 4164 1369
rect 4130 1267 4164 1301
rect 4130 1199 4164 1233
rect 4130 1131 4164 1165
rect 4130 1063 4164 1097
rect 4130 995 4164 1029
rect 4130 927 4164 961
rect 4130 859 4164 893
rect 4130 791 4164 825
rect 4130 723 4164 757
rect 4130 655 4164 689
rect 4130 325 4164 621
rect 4290 2560 4324 2650
rect 4290 2492 4324 2510
rect 4290 2424 4324 2438
rect 4290 2356 4324 2366
rect 4290 2288 4324 2294
rect 4290 2220 4324 2222
rect 4290 2184 4324 2186
rect 4290 2112 4324 2118
rect 4290 2040 4324 2050
rect 4290 1968 4324 1982
rect 4290 1896 4324 1914
rect 4290 1824 4324 1846
rect 4290 1752 4324 1778
rect 4290 1680 4324 1710
rect 4290 1608 4324 1642
rect 4290 1540 4324 1574
rect 4290 1472 4324 1502
rect 4290 1404 4324 1430
rect 4290 1336 4324 1358
rect 4290 1268 4324 1286
rect 4290 1200 4324 1214
rect 4290 1132 4324 1142
rect 4290 1064 4324 1070
rect 4290 996 4324 998
rect 4290 960 4324 962
rect 4290 888 4324 894
rect 4290 816 4324 826
rect 4290 744 4324 758
rect 4290 672 4324 690
rect 4290 587 4324 622
rect 4378 2560 4412 2755
rect 4447 2703 4519 2721
rect 4447 2669 4466 2703
rect 4500 2669 4519 2703
rect 4447 2651 4519 2669
rect 4378 2492 4412 2510
rect 4378 2424 4412 2438
rect 4378 2356 4412 2366
rect 4378 2288 4412 2294
rect 4378 2220 4412 2222
rect 4378 2184 4412 2186
rect 4378 2112 4412 2118
rect 4378 2040 4412 2050
rect 4378 1968 4412 1982
rect 4378 1896 4412 1914
rect 4378 1824 4412 1846
rect 4378 1752 4412 1778
rect 4378 1680 4412 1710
rect 4378 1608 4412 1642
rect 4378 1540 4412 1574
rect 4378 1472 4412 1502
rect 4378 1404 4412 1430
rect 4378 1336 4412 1358
rect 4378 1268 4412 1286
rect 4378 1200 4412 1214
rect 4378 1132 4412 1142
rect 4378 1064 4412 1070
rect 4378 996 4412 998
rect 4378 960 4412 962
rect 4378 888 4412 894
rect 4378 816 4412 826
rect 4378 744 4412 758
rect 4378 672 4412 690
rect 4378 587 4412 622
rect 4466 2560 4500 2651
rect 4466 2492 4500 2510
rect 4466 2424 4500 2438
rect 4466 2356 4500 2366
rect 4466 2288 4500 2294
rect 4466 2220 4500 2222
rect 4466 2184 4500 2186
rect 4466 2112 4500 2118
rect 4466 2040 4500 2050
rect 4466 1968 4500 1982
rect 4466 1896 4500 1914
rect 4466 1824 4500 1846
rect 4466 1752 4500 1778
rect 4466 1680 4500 1710
rect 4466 1608 4500 1642
rect 4466 1540 4500 1574
rect 4466 1472 4500 1502
rect 4466 1404 4500 1430
rect 4466 1336 4500 1358
rect 4466 1268 4500 1286
rect 4466 1200 4500 1214
rect 4466 1132 4500 1142
rect 4466 1064 4500 1070
rect 4466 996 4500 998
rect 4466 960 4500 962
rect 4466 888 4500 894
rect 4466 816 4500 826
rect 4466 744 4500 758
rect 4466 672 4500 690
rect 4466 587 4500 622
rect 4554 2560 4588 2755
rect 4623 2703 4695 2721
rect 4623 2669 4642 2703
rect 4676 2669 4695 2703
rect 4623 2651 4695 2669
rect 4554 2492 4588 2510
rect 4554 2424 4588 2438
rect 4554 2356 4588 2366
rect 4554 2288 4588 2294
rect 4554 2220 4588 2222
rect 4554 2184 4588 2186
rect 4554 2112 4588 2118
rect 4554 2040 4588 2050
rect 4554 1968 4588 1982
rect 4554 1896 4588 1914
rect 4554 1824 4588 1846
rect 4554 1752 4588 1778
rect 4554 1680 4588 1710
rect 4554 1608 4588 1642
rect 4554 1540 4588 1574
rect 4554 1472 4588 1502
rect 4554 1404 4588 1430
rect 4554 1336 4588 1358
rect 4554 1268 4588 1286
rect 4554 1200 4588 1214
rect 4554 1132 4588 1142
rect 4554 1064 4588 1070
rect 4554 996 4588 998
rect 4554 960 4588 962
rect 4554 888 4588 894
rect 4554 816 4588 826
rect 4554 744 4588 758
rect 4554 672 4588 690
rect 4554 587 4588 622
rect 4642 2560 4676 2651
rect 4642 2492 4676 2510
rect 4642 2424 4676 2438
rect 4642 2356 4676 2366
rect 4642 2288 4676 2294
rect 4642 2220 4676 2222
rect 4642 2184 4676 2186
rect 4642 2112 4676 2118
rect 4642 2040 4676 2050
rect 4642 1968 4676 1982
rect 4642 1896 4676 1914
rect 4642 1824 4676 1846
rect 4642 1752 4676 1778
rect 4642 1680 4676 1710
rect 4642 1608 4676 1642
rect 4642 1540 4676 1574
rect 4642 1472 4676 1502
rect 4642 1404 4676 1430
rect 4642 1336 4676 1358
rect 4642 1268 4676 1286
rect 4642 1200 4676 1214
rect 4642 1132 4676 1142
rect 4642 1064 4676 1070
rect 4642 996 4676 998
rect 4642 960 4676 962
rect 4642 888 4676 894
rect 4642 816 4676 826
rect 4642 744 4676 758
rect 4642 672 4676 690
rect 4642 587 4676 622
rect 4730 2560 4764 2755
rect 4799 2703 4871 2721
rect 4799 2669 4818 2703
rect 4852 2669 4871 2703
rect 4799 2651 4871 2669
rect 4730 2492 4764 2510
rect 4730 2424 4764 2438
rect 4730 2356 4764 2366
rect 4730 2288 4764 2294
rect 4730 2220 4764 2222
rect 4730 2184 4764 2186
rect 4730 2112 4764 2118
rect 4730 2040 4764 2050
rect 4730 1968 4764 1982
rect 4730 1896 4764 1914
rect 4730 1824 4764 1846
rect 4730 1752 4764 1778
rect 4730 1680 4764 1710
rect 4730 1608 4764 1642
rect 4730 1540 4764 1574
rect 4730 1472 4764 1502
rect 4730 1404 4764 1430
rect 4730 1336 4764 1358
rect 4730 1268 4764 1286
rect 4730 1200 4764 1214
rect 4730 1132 4764 1142
rect 4730 1064 4764 1070
rect 4730 996 4764 998
rect 4730 960 4764 962
rect 4730 888 4764 894
rect 4730 816 4764 826
rect 4730 744 4764 758
rect 4730 672 4764 690
rect 4730 587 4764 622
rect 4818 2560 4852 2651
rect 4818 2492 4852 2510
rect 4818 2424 4852 2438
rect 4818 2356 4852 2366
rect 4818 2288 4852 2294
rect 4818 2220 4852 2222
rect 4818 2184 4852 2186
rect 4818 2112 4852 2118
rect 4818 2040 4852 2050
rect 4818 1968 4852 1982
rect 4818 1896 4852 1914
rect 4818 1824 4852 1846
rect 4818 1752 4852 1778
rect 4818 1680 4852 1710
rect 4818 1608 4852 1642
rect 4818 1540 4852 1574
rect 4818 1472 4852 1502
rect 4818 1404 4852 1430
rect 4818 1336 4852 1358
rect 4818 1268 4852 1286
rect 4818 1200 4852 1214
rect 4818 1132 4852 1142
rect 4818 1064 4852 1070
rect 4818 996 4852 998
rect 4818 960 4852 962
rect 4818 888 4852 894
rect 4818 816 4852 826
rect 4818 744 4852 758
rect 4818 672 4852 690
rect 4818 587 4852 622
rect 4906 2560 4940 2755
rect 4975 2703 5047 2721
rect 4975 2669 4994 2703
rect 5028 2669 5047 2703
rect 4975 2651 5047 2669
rect 4906 2492 4940 2510
rect 4906 2424 4940 2438
rect 4906 2356 4940 2366
rect 4906 2288 4940 2294
rect 4906 2220 4940 2222
rect 4906 2184 4940 2186
rect 4906 2112 4940 2118
rect 4906 2040 4940 2050
rect 4906 1968 4940 1982
rect 4906 1896 4940 1914
rect 4906 1824 4940 1846
rect 4906 1752 4940 1778
rect 4906 1680 4940 1710
rect 4906 1608 4940 1642
rect 4906 1540 4940 1574
rect 4906 1472 4940 1502
rect 4906 1404 4940 1430
rect 4906 1336 4940 1358
rect 4906 1268 4940 1286
rect 4906 1200 4940 1214
rect 4906 1132 4940 1142
rect 4906 1064 4940 1070
rect 4906 996 4940 998
rect 4906 960 4940 962
rect 4906 888 4940 894
rect 4906 816 4940 826
rect 4906 744 4940 758
rect 4906 672 4940 690
rect 4906 587 4940 622
rect 4994 2560 5028 2651
rect 4994 2492 5028 2510
rect 4994 2424 5028 2438
rect 4994 2356 5028 2366
rect 4994 2288 5028 2294
rect 4994 2220 5028 2222
rect 4994 2184 5028 2186
rect 4994 2112 5028 2118
rect 4994 2040 5028 2050
rect 4994 1968 5028 1982
rect 4994 1896 5028 1914
rect 4994 1824 5028 1846
rect 4994 1752 5028 1778
rect 4994 1680 5028 1710
rect 4994 1608 5028 1642
rect 4994 1540 5028 1574
rect 4994 1472 5028 1502
rect 4994 1404 5028 1430
rect 4994 1336 5028 1358
rect 4994 1268 5028 1286
rect 4994 1200 5028 1214
rect 4994 1132 5028 1142
rect 4994 1064 5028 1070
rect 4994 996 5028 998
rect 4994 960 5028 962
rect 4994 888 5028 894
rect 4994 816 5028 826
rect 4994 744 5028 758
rect 4994 672 5028 690
rect 4994 587 5028 622
rect 5082 2560 5116 2755
rect 5151 2703 5223 2721
rect 5151 2669 5170 2703
rect 5204 2669 5223 2703
rect 5151 2651 5223 2669
rect 5082 2492 5116 2510
rect 5082 2424 5116 2438
rect 5082 2356 5116 2366
rect 5082 2288 5116 2294
rect 5082 2220 5116 2222
rect 5082 2184 5116 2186
rect 5082 2112 5116 2118
rect 5082 2040 5116 2050
rect 5082 1968 5116 1982
rect 5082 1896 5116 1914
rect 5082 1824 5116 1846
rect 5082 1752 5116 1778
rect 5082 1680 5116 1710
rect 5082 1608 5116 1642
rect 5082 1540 5116 1574
rect 5082 1472 5116 1502
rect 5082 1404 5116 1430
rect 5082 1336 5116 1358
rect 5082 1268 5116 1286
rect 5082 1200 5116 1214
rect 5082 1132 5116 1142
rect 5082 1064 5116 1070
rect 5082 996 5116 998
rect 5082 960 5116 962
rect 5082 888 5116 894
rect 5082 816 5116 826
rect 5082 744 5116 758
rect 5082 672 5116 690
rect 5082 587 5116 622
rect 5170 2560 5204 2651
rect 5170 2492 5204 2510
rect 5170 2424 5204 2438
rect 5170 2356 5204 2366
rect 5170 2288 5204 2294
rect 5170 2220 5204 2222
rect 5170 2184 5204 2186
rect 5170 2112 5204 2118
rect 5170 2040 5204 2050
rect 5170 1968 5204 1982
rect 5170 1896 5204 1914
rect 5170 1824 5204 1846
rect 5170 1752 5204 1778
rect 5170 1680 5204 1710
rect 5170 1608 5204 1642
rect 5170 1540 5204 1574
rect 5170 1472 5204 1502
rect 5170 1404 5204 1430
rect 5170 1336 5204 1358
rect 5170 1268 5204 1286
rect 5170 1200 5204 1214
rect 5170 1132 5204 1142
rect 5170 1064 5204 1070
rect 5170 996 5204 998
rect 5170 960 5204 962
rect 5170 888 5204 894
rect 5170 816 5204 826
rect 5170 744 5204 758
rect 5170 672 5204 690
rect 5170 587 5204 622
rect 5258 2560 5292 2755
rect 5386 2721 5420 2969
rect 5348 2703 5420 2721
rect 5348 2669 5367 2703
rect 5401 2669 5420 2703
rect 5348 2651 5420 2669
rect 5258 2492 5292 2510
rect 5258 2424 5292 2438
rect 5258 2356 5292 2366
rect 5258 2288 5292 2294
rect 5258 2220 5292 2222
rect 5258 2184 5292 2186
rect 5258 2112 5292 2118
rect 5258 2040 5292 2050
rect 5258 1968 5292 1982
rect 5258 1896 5292 1914
rect 5258 1824 5292 1846
rect 5258 1752 5292 1778
rect 5258 1680 5292 1710
rect 5258 1608 5292 1642
rect 5258 1540 5292 1574
rect 5258 1472 5292 1502
rect 5258 1404 5292 1430
rect 5258 1336 5292 1358
rect 5258 1268 5292 1286
rect 5258 1200 5292 1214
rect 5258 1132 5292 1142
rect 5258 1064 5292 1070
rect 5258 996 5292 998
rect 5258 960 5292 962
rect 5258 888 5292 894
rect 5258 816 5292 826
rect 5258 744 5292 758
rect 5258 672 5292 690
rect 5258 587 5292 622
rect 5386 2555 5420 2651
rect 5386 2487 5420 2521
rect 5386 2419 5420 2453
rect 5386 2351 5420 2385
rect 5386 2283 5420 2317
rect 5386 2215 5420 2249
rect 5386 2147 5420 2181
rect 5386 2079 5420 2113
rect 5386 2011 5420 2045
rect 5386 1943 5420 1977
rect 5386 1875 5420 1909
rect 5386 1807 5420 1841
rect 5386 1739 5420 1773
rect 5386 1671 5420 1705
rect 5386 1603 5420 1637
rect 5386 1535 5420 1569
rect 5386 1467 5420 1501
rect 5386 1399 5420 1433
rect 5386 1331 5420 1365
rect 5386 1263 5420 1297
rect 5386 1195 5420 1229
rect 5386 1127 5420 1161
rect 5386 1059 5420 1093
rect 5386 991 5420 1025
rect 5386 923 5420 957
rect 5386 855 5420 889
rect 5386 787 5420 821
rect 5386 719 5420 753
rect 5386 651 5420 685
rect 4336 524 5159 553
rect 4336 475 4378 524
rect 4412 475 4554 524
rect 4588 475 4730 524
rect 4764 475 4906 524
rect 4940 475 5082 524
rect 5116 475 5159 524
rect 4336 418 5159 475
rect 5386 325 5420 617
rect 4130 324 5420 325
rect 4130 290 4364 324
rect 4398 290 4432 324
rect 4466 290 4500 324
rect 4534 290 4568 324
rect 4602 290 4636 324
rect 4670 290 4704 324
rect 4738 290 4772 324
rect 4806 290 4840 324
rect 4874 290 4908 324
rect 4942 290 4976 324
rect 5010 290 5044 324
rect 5078 290 5112 324
rect 5146 290 5180 324
rect 5214 290 5420 324
rect 4130 289 5420 290
<< viali >>
rect 699 3406 733 3440
rect 299 2958 333 2992
rect 875 3406 909 3440
rect 1051 3406 1085 3440
rect 2811 3406 2845 3440
rect 2987 3406 3021 3440
rect 3163 3406 3197 3440
rect 3687 2958 3721 2992
rect 4290 2843 4324 2877
rect 4466 2843 4500 2877
rect 4642 2843 4676 2877
rect 4818 2843 4852 2877
rect 4994 2843 5028 2877
rect 5170 2843 5204 2877
rect 4378 2773 4412 2807
rect 4554 2773 4588 2807
rect 4730 2773 4764 2807
rect 4906 2773 4940 2807
rect 5082 2773 5116 2807
rect 5258 2773 5292 2807
rect 4149 2668 4183 2702
rect 4290 2669 4324 2703
rect 4290 2526 4324 2544
rect 4290 2510 4324 2526
rect 4290 2458 4324 2472
rect 4290 2438 4324 2458
rect 4290 2390 4324 2400
rect 4290 2366 4324 2390
rect 4290 2322 4324 2328
rect 4290 2294 4324 2322
rect 4290 2254 4324 2256
rect 4290 2222 4324 2254
rect 4290 2152 4324 2184
rect 4290 2150 4324 2152
rect 4290 2084 4324 2112
rect 4290 2078 4324 2084
rect 4290 2016 4324 2040
rect 4290 2006 4324 2016
rect 4290 1948 4324 1968
rect 4290 1934 4324 1948
rect 4290 1880 4324 1896
rect 4290 1862 4324 1880
rect 4290 1812 4324 1824
rect 4290 1790 4324 1812
rect 4290 1744 4324 1752
rect 4290 1718 4324 1744
rect 4290 1676 4324 1680
rect 4290 1646 4324 1676
rect 4290 1574 4324 1608
rect 4290 1506 4324 1536
rect 4290 1502 4324 1506
rect 4290 1438 4324 1464
rect 4290 1430 4324 1438
rect 4290 1370 4324 1392
rect 4290 1358 4324 1370
rect 4290 1302 4324 1320
rect 4290 1286 4324 1302
rect 4290 1234 4324 1248
rect 4290 1214 4324 1234
rect 4290 1166 4324 1176
rect 4290 1142 4324 1166
rect 4290 1098 4324 1104
rect 4290 1070 4324 1098
rect 4290 1030 4324 1032
rect 4290 998 4324 1030
rect 4290 928 4324 960
rect 4290 926 4324 928
rect 4290 860 4324 888
rect 4290 854 4324 860
rect 4290 792 4324 816
rect 4290 782 4324 792
rect 4290 724 4324 744
rect 4290 710 4324 724
rect 4290 656 4324 672
rect 4290 638 4324 656
rect 4466 2669 4500 2703
rect 4378 2526 4412 2544
rect 4378 2510 4412 2526
rect 4378 2458 4412 2472
rect 4378 2438 4412 2458
rect 4378 2390 4412 2400
rect 4378 2366 4412 2390
rect 4378 2322 4412 2328
rect 4378 2294 4412 2322
rect 4378 2254 4412 2256
rect 4378 2222 4412 2254
rect 4378 2152 4412 2184
rect 4378 2150 4412 2152
rect 4378 2084 4412 2112
rect 4378 2078 4412 2084
rect 4378 2016 4412 2040
rect 4378 2006 4412 2016
rect 4378 1948 4412 1968
rect 4378 1934 4412 1948
rect 4378 1880 4412 1896
rect 4378 1862 4412 1880
rect 4378 1812 4412 1824
rect 4378 1790 4412 1812
rect 4378 1744 4412 1752
rect 4378 1718 4412 1744
rect 4378 1676 4412 1680
rect 4378 1646 4412 1676
rect 4378 1574 4412 1608
rect 4378 1506 4412 1536
rect 4378 1502 4412 1506
rect 4378 1438 4412 1464
rect 4378 1430 4412 1438
rect 4378 1370 4412 1392
rect 4378 1358 4412 1370
rect 4378 1302 4412 1320
rect 4378 1286 4412 1302
rect 4378 1234 4412 1248
rect 4378 1214 4412 1234
rect 4378 1166 4412 1176
rect 4378 1142 4412 1166
rect 4378 1098 4412 1104
rect 4378 1070 4412 1098
rect 4378 1030 4412 1032
rect 4378 998 4412 1030
rect 4378 928 4412 960
rect 4378 926 4412 928
rect 4378 860 4412 888
rect 4378 854 4412 860
rect 4378 792 4412 816
rect 4378 782 4412 792
rect 4378 724 4412 744
rect 4378 710 4412 724
rect 4378 656 4412 672
rect 4378 638 4412 656
rect 4466 2526 4500 2544
rect 4466 2510 4500 2526
rect 4466 2458 4500 2472
rect 4466 2438 4500 2458
rect 4466 2390 4500 2400
rect 4466 2366 4500 2390
rect 4466 2322 4500 2328
rect 4466 2294 4500 2322
rect 4466 2254 4500 2256
rect 4466 2222 4500 2254
rect 4466 2152 4500 2184
rect 4466 2150 4500 2152
rect 4466 2084 4500 2112
rect 4466 2078 4500 2084
rect 4466 2016 4500 2040
rect 4466 2006 4500 2016
rect 4466 1948 4500 1968
rect 4466 1934 4500 1948
rect 4466 1880 4500 1896
rect 4466 1862 4500 1880
rect 4466 1812 4500 1824
rect 4466 1790 4500 1812
rect 4466 1744 4500 1752
rect 4466 1718 4500 1744
rect 4466 1676 4500 1680
rect 4466 1646 4500 1676
rect 4466 1574 4500 1608
rect 4466 1506 4500 1536
rect 4466 1502 4500 1506
rect 4466 1438 4500 1464
rect 4466 1430 4500 1438
rect 4466 1370 4500 1392
rect 4466 1358 4500 1370
rect 4466 1302 4500 1320
rect 4466 1286 4500 1302
rect 4466 1234 4500 1248
rect 4466 1214 4500 1234
rect 4466 1166 4500 1176
rect 4466 1142 4500 1166
rect 4466 1098 4500 1104
rect 4466 1070 4500 1098
rect 4466 1030 4500 1032
rect 4466 998 4500 1030
rect 4466 928 4500 960
rect 4466 926 4500 928
rect 4466 860 4500 888
rect 4466 854 4500 860
rect 4466 792 4500 816
rect 4466 782 4500 792
rect 4466 724 4500 744
rect 4466 710 4500 724
rect 4466 656 4500 672
rect 4466 638 4500 656
rect 4642 2669 4676 2703
rect 4554 2526 4588 2544
rect 4554 2510 4588 2526
rect 4554 2458 4588 2472
rect 4554 2438 4588 2458
rect 4554 2390 4588 2400
rect 4554 2366 4588 2390
rect 4554 2322 4588 2328
rect 4554 2294 4588 2322
rect 4554 2254 4588 2256
rect 4554 2222 4588 2254
rect 4554 2152 4588 2184
rect 4554 2150 4588 2152
rect 4554 2084 4588 2112
rect 4554 2078 4588 2084
rect 4554 2016 4588 2040
rect 4554 2006 4588 2016
rect 4554 1948 4588 1968
rect 4554 1934 4588 1948
rect 4554 1880 4588 1896
rect 4554 1862 4588 1880
rect 4554 1812 4588 1824
rect 4554 1790 4588 1812
rect 4554 1744 4588 1752
rect 4554 1718 4588 1744
rect 4554 1676 4588 1680
rect 4554 1646 4588 1676
rect 4554 1574 4588 1608
rect 4554 1506 4588 1536
rect 4554 1502 4588 1506
rect 4554 1438 4588 1464
rect 4554 1430 4588 1438
rect 4554 1370 4588 1392
rect 4554 1358 4588 1370
rect 4554 1302 4588 1320
rect 4554 1286 4588 1302
rect 4554 1234 4588 1248
rect 4554 1214 4588 1234
rect 4554 1166 4588 1176
rect 4554 1142 4588 1166
rect 4554 1098 4588 1104
rect 4554 1070 4588 1098
rect 4554 1030 4588 1032
rect 4554 998 4588 1030
rect 4554 928 4588 960
rect 4554 926 4588 928
rect 4554 860 4588 888
rect 4554 854 4588 860
rect 4554 792 4588 816
rect 4554 782 4588 792
rect 4554 724 4588 744
rect 4554 710 4588 724
rect 4554 656 4588 672
rect 4554 638 4588 656
rect 4642 2526 4676 2544
rect 4642 2510 4676 2526
rect 4642 2458 4676 2472
rect 4642 2438 4676 2458
rect 4642 2390 4676 2400
rect 4642 2366 4676 2390
rect 4642 2322 4676 2328
rect 4642 2294 4676 2322
rect 4642 2254 4676 2256
rect 4642 2222 4676 2254
rect 4642 2152 4676 2184
rect 4642 2150 4676 2152
rect 4642 2084 4676 2112
rect 4642 2078 4676 2084
rect 4642 2016 4676 2040
rect 4642 2006 4676 2016
rect 4642 1948 4676 1968
rect 4642 1934 4676 1948
rect 4642 1880 4676 1896
rect 4642 1862 4676 1880
rect 4642 1812 4676 1824
rect 4642 1790 4676 1812
rect 4642 1744 4676 1752
rect 4642 1718 4676 1744
rect 4642 1676 4676 1680
rect 4642 1646 4676 1676
rect 4642 1574 4676 1608
rect 4642 1506 4676 1536
rect 4642 1502 4676 1506
rect 4642 1438 4676 1464
rect 4642 1430 4676 1438
rect 4642 1370 4676 1392
rect 4642 1358 4676 1370
rect 4642 1302 4676 1320
rect 4642 1286 4676 1302
rect 4642 1234 4676 1248
rect 4642 1214 4676 1234
rect 4642 1166 4676 1176
rect 4642 1142 4676 1166
rect 4642 1098 4676 1104
rect 4642 1070 4676 1098
rect 4642 1030 4676 1032
rect 4642 998 4676 1030
rect 4642 928 4676 960
rect 4642 926 4676 928
rect 4642 860 4676 888
rect 4642 854 4676 860
rect 4642 792 4676 816
rect 4642 782 4676 792
rect 4642 724 4676 744
rect 4642 710 4676 724
rect 4642 656 4676 672
rect 4642 638 4676 656
rect 4818 2669 4852 2703
rect 4730 2526 4764 2544
rect 4730 2510 4764 2526
rect 4730 2458 4764 2472
rect 4730 2438 4764 2458
rect 4730 2390 4764 2400
rect 4730 2366 4764 2390
rect 4730 2322 4764 2328
rect 4730 2294 4764 2322
rect 4730 2254 4764 2256
rect 4730 2222 4764 2254
rect 4730 2152 4764 2184
rect 4730 2150 4764 2152
rect 4730 2084 4764 2112
rect 4730 2078 4764 2084
rect 4730 2016 4764 2040
rect 4730 2006 4764 2016
rect 4730 1948 4764 1968
rect 4730 1934 4764 1948
rect 4730 1880 4764 1896
rect 4730 1862 4764 1880
rect 4730 1812 4764 1824
rect 4730 1790 4764 1812
rect 4730 1744 4764 1752
rect 4730 1718 4764 1744
rect 4730 1676 4764 1680
rect 4730 1646 4764 1676
rect 4730 1574 4764 1608
rect 4730 1506 4764 1536
rect 4730 1502 4764 1506
rect 4730 1438 4764 1464
rect 4730 1430 4764 1438
rect 4730 1370 4764 1392
rect 4730 1358 4764 1370
rect 4730 1302 4764 1320
rect 4730 1286 4764 1302
rect 4730 1234 4764 1248
rect 4730 1214 4764 1234
rect 4730 1166 4764 1176
rect 4730 1142 4764 1166
rect 4730 1098 4764 1104
rect 4730 1070 4764 1098
rect 4730 1030 4764 1032
rect 4730 998 4764 1030
rect 4730 928 4764 960
rect 4730 926 4764 928
rect 4730 860 4764 888
rect 4730 854 4764 860
rect 4730 792 4764 816
rect 4730 782 4764 792
rect 4730 724 4764 744
rect 4730 710 4764 724
rect 4730 656 4764 672
rect 4730 638 4764 656
rect 4818 2526 4852 2544
rect 4818 2510 4852 2526
rect 4818 2458 4852 2472
rect 4818 2438 4852 2458
rect 4818 2390 4852 2400
rect 4818 2366 4852 2390
rect 4818 2322 4852 2328
rect 4818 2294 4852 2322
rect 4818 2254 4852 2256
rect 4818 2222 4852 2254
rect 4818 2152 4852 2184
rect 4818 2150 4852 2152
rect 4818 2084 4852 2112
rect 4818 2078 4852 2084
rect 4818 2016 4852 2040
rect 4818 2006 4852 2016
rect 4818 1948 4852 1968
rect 4818 1934 4852 1948
rect 4818 1880 4852 1896
rect 4818 1862 4852 1880
rect 4818 1812 4852 1824
rect 4818 1790 4852 1812
rect 4818 1744 4852 1752
rect 4818 1718 4852 1744
rect 4818 1676 4852 1680
rect 4818 1646 4852 1676
rect 4818 1574 4852 1608
rect 4818 1506 4852 1536
rect 4818 1502 4852 1506
rect 4818 1438 4852 1464
rect 4818 1430 4852 1438
rect 4818 1370 4852 1392
rect 4818 1358 4852 1370
rect 4818 1302 4852 1320
rect 4818 1286 4852 1302
rect 4818 1234 4852 1248
rect 4818 1214 4852 1234
rect 4818 1166 4852 1176
rect 4818 1142 4852 1166
rect 4818 1098 4852 1104
rect 4818 1070 4852 1098
rect 4818 1030 4852 1032
rect 4818 998 4852 1030
rect 4818 928 4852 960
rect 4818 926 4852 928
rect 4818 860 4852 888
rect 4818 854 4852 860
rect 4818 792 4852 816
rect 4818 782 4852 792
rect 4818 724 4852 744
rect 4818 710 4852 724
rect 4818 656 4852 672
rect 4818 638 4852 656
rect 4994 2669 5028 2703
rect 4906 2526 4940 2544
rect 4906 2510 4940 2526
rect 4906 2458 4940 2472
rect 4906 2438 4940 2458
rect 4906 2390 4940 2400
rect 4906 2366 4940 2390
rect 4906 2322 4940 2328
rect 4906 2294 4940 2322
rect 4906 2254 4940 2256
rect 4906 2222 4940 2254
rect 4906 2152 4940 2184
rect 4906 2150 4940 2152
rect 4906 2084 4940 2112
rect 4906 2078 4940 2084
rect 4906 2016 4940 2040
rect 4906 2006 4940 2016
rect 4906 1948 4940 1968
rect 4906 1934 4940 1948
rect 4906 1880 4940 1896
rect 4906 1862 4940 1880
rect 4906 1812 4940 1824
rect 4906 1790 4940 1812
rect 4906 1744 4940 1752
rect 4906 1718 4940 1744
rect 4906 1676 4940 1680
rect 4906 1646 4940 1676
rect 4906 1574 4940 1608
rect 4906 1506 4940 1536
rect 4906 1502 4940 1506
rect 4906 1438 4940 1464
rect 4906 1430 4940 1438
rect 4906 1370 4940 1392
rect 4906 1358 4940 1370
rect 4906 1302 4940 1320
rect 4906 1286 4940 1302
rect 4906 1234 4940 1248
rect 4906 1214 4940 1234
rect 4906 1166 4940 1176
rect 4906 1142 4940 1166
rect 4906 1098 4940 1104
rect 4906 1070 4940 1098
rect 4906 1030 4940 1032
rect 4906 998 4940 1030
rect 4906 928 4940 960
rect 4906 926 4940 928
rect 4906 860 4940 888
rect 4906 854 4940 860
rect 4906 792 4940 816
rect 4906 782 4940 792
rect 4906 724 4940 744
rect 4906 710 4940 724
rect 4906 656 4940 672
rect 4906 638 4940 656
rect 4994 2526 5028 2544
rect 4994 2510 5028 2526
rect 4994 2458 5028 2472
rect 4994 2438 5028 2458
rect 4994 2390 5028 2400
rect 4994 2366 5028 2390
rect 4994 2322 5028 2328
rect 4994 2294 5028 2322
rect 4994 2254 5028 2256
rect 4994 2222 5028 2254
rect 4994 2152 5028 2184
rect 4994 2150 5028 2152
rect 4994 2084 5028 2112
rect 4994 2078 5028 2084
rect 4994 2016 5028 2040
rect 4994 2006 5028 2016
rect 4994 1948 5028 1968
rect 4994 1934 5028 1948
rect 4994 1880 5028 1896
rect 4994 1862 5028 1880
rect 4994 1812 5028 1824
rect 4994 1790 5028 1812
rect 4994 1744 5028 1752
rect 4994 1718 5028 1744
rect 4994 1676 5028 1680
rect 4994 1646 5028 1676
rect 4994 1574 5028 1608
rect 4994 1506 5028 1536
rect 4994 1502 5028 1506
rect 4994 1438 5028 1464
rect 4994 1430 5028 1438
rect 4994 1370 5028 1392
rect 4994 1358 5028 1370
rect 4994 1302 5028 1320
rect 4994 1286 5028 1302
rect 4994 1234 5028 1248
rect 4994 1214 5028 1234
rect 4994 1166 5028 1176
rect 4994 1142 5028 1166
rect 4994 1098 5028 1104
rect 4994 1070 5028 1098
rect 4994 1030 5028 1032
rect 4994 998 5028 1030
rect 4994 928 5028 960
rect 4994 926 5028 928
rect 4994 860 5028 888
rect 4994 854 5028 860
rect 4994 792 5028 816
rect 4994 782 5028 792
rect 4994 724 5028 744
rect 4994 710 5028 724
rect 4994 656 5028 672
rect 4994 638 5028 656
rect 5170 2669 5204 2703
rect 5082 2526 5116 2544
rect 5082 2510 5116 2526
rect 5082 2458 5116 2472
rect 5082 2438 5116 2458
rect 5082 2390 5116 2400
rect 5082 2366 5116 2390
rect 5082 2322 5116 2328
rect 5082 2294 5116 2322
rect 5082 2254 5116 2256
rect 5082 2222 5116 2254
rect 5082 2152 5116 2184
rect 5082 2150 5116 2152
rect 5082 2084 5116 2112
rect 5082 2078 5116 2084
rect 5082 2016 5116 2040
rect 5082 2006 5116 2016
rect 5082 1948 5116 1968
rect 5082 1934 5116 1948
rect 5082 1880 5116 1896
rect 5082 1862 5116 1880
rect 5082 1812 5116 1824
rect 5082 1790 5116 1812
rect 5082 1744 5116 1752
rect 5082 1718 5116 1744
rect 5082 1676 5116 1680
rect 5082 1646 5116 1676
rect 5082 1574 5116 1608
rect 5082 1506 5116 1536
rect 5082 1502 5116 1506
rect 5082 1438 5116 1464
rect 5082 1430 5116 1438
rect 5082 1370 5116 1392
rect 5082 1358 5116 1370
rect 5082 1302 5116 1320
rect 5082 1286 5116 1302
rect 5082 1234 5116 1248
rect 5082 1214 5116 1234
rect 5082 1166 5116 1176
rect 5082 1142 5116 1166
rect 5082 1098 5116 1104
rect 5082 1070 5116 1098
rect 5082 1030 5116 1032
rect 5082 998 5116 1030
rect 5082 928 5116 960
rect 5082 926 5116 928
rect 5082 860 5116 888
rect 5082 854 5116 860
rect 5082 792 5116 816
rect 5082 782 5116 792
rect 5082 724 5116 744
rect 5082 710 5116 724
rect 5082 656 5116 672
rect 5082 638 5116 656
rect 5170 2526 5204 2544
rect 5170 2510 5204 2526
rect 5170 2458 5204 2472
rect 5170 2438 5204 2458
rect 5170 2390 5204 2400
rect 5170 2366 5204 2390
rect 5170 2322 5204 2328
rect 5170 2294 5204 2322
rect 5170 2254 5204 2256
rect 5170 2222 5204 2254
rect 5170 2152 5204 2184
rect 5170 2150 5204 2152
rect 5170 2084 5204 2112
rect 5170 2078 5204 2084
rect 5170 2016 5204 2040
rect 5170 2006 5204 2016
rect 5170 1948 5204 1968
rect 5170 1934 5204 1948
rect 5170 1880 5204 1896
rect 5170 1862 5204 1880
rect 5170 1812 5204 1824
rect 5170 1790 5204 1812
rect 5170 1744 5204 1752
rect 5170 1718 5204 1744
rect 5170 1676 5204 1680
rect 5170 1646 5204 1676
rect 5170 1574 5204 1608
rect 5170 1506 5204 1536
rect 5170 1502 5204 1506
rect 5170 1438 5204 1464
rect 5170 1430 5204 1438
rect 5170 1370 5204 1392
rect 5170 1358 5204 1370
rect 5170 1302 5204 1320
rect 5170 1286 5204 1302
rect 5170 1234 5204 1248
rect 5170 1214 5204 1234
rect 5170 1166 5204 1176
rect 5170 1142 5204 1166
rect 5170 1098 5204 1104
rect 5170 1070 5204 1098
rect 5170 1030 5204 1032
rect 5170 998 5204 1030
rect 5170 928 5204 960
rect 5170 926 5204 928
rect 5170 860 5204 888
rect 5170 854 5204 860
rect 5170 792 5204 816
rect 5170 782 5204 792
rect 5170 724 5204 744
rect 5170 710 5204 724
rect 5170 656 5204 672
rect 5170 638 5204 656
rect 5367 2669 5401 2703
rect 5258 2526 5292 2544
rect 5258 2510 5292 2526
rect 5258 2458 5292 2472
rect 5258 2438 5292 2458
rect 5258 2390 5292 2400
rect 5258 2366 5292 2390
rect 5258 2322 5292 2328
rect 5258 2294 5292 2322
rect 5258 2254 5292 2256
rect 5258 2222 5292 2254
rect 5258 2152 5292 2184
rect 5258 2150 5292 2152
rect 5258 2084 5292 2112
rect 5258 2078 5292 2084
rect 5258 2016 5292 2040
rect 5258 2006 5292 2016
rect 5258 1948 5292 1968
rect 5258 1934 5292 1948
rect 5258 1880 5292 1896
rect 5258 1862 5292 1880
rect 5258 1812 5292 1824
rect 5258 1790 5292 1812
rect 5258 1744 5292 1752
rect 5258 1718 5292 1744
rect 5258 1676 5292 1680
rect 5258 1646 5292 1676
rect 5258 1574 5292 1608
rect 5258 1506 5292 1536
rect 5258 1502 5292 1506
rect 5258 1438 5292 1464
rect 5258 1430 5292 1438
rect 5258 1370 5292 1392
rect 5258 1358 5292 1370
rect 5258 1302 5292 1320
rect 5258 1286 5292 1302
rect 5258 1234 5292 1248
rect 5258 1214 5292 1234
rect 5258 1166 5292 1176
rect 5258 1142 5292 1166
rect 5258 1098 5292 1104
rect 5258 1070 5292 1098
rect 5258 1030 5292 1032
rect 5258 998 5292 1030
rect 5258 928 5292 960
rect 5258 926 5292 928
rect 5258 860 5292 888
rect 5258 854 5292 860
rect 5258 792 5292 816
rect 5258 782 5292 792
rect 5258 724 5292 744
rect 5258 710 5292 724
rect 5258 656 5292 672
rect 5258 638 5292 656
rect 4378 490 4412 509
rect 4378 475 4412 490
rect 4554 490 4588 509
rect 4554 475 4588 490
rect 4730 490 4764 509
rect 4730 475 4764 490
rect 4906 490 4940 509
rect 4906 475 4940 490
rect 5082 490 5116 509
rect 5082 475 5116 490
<< metal1 >>
rect 279 3440 1104 3458
rect 279 3406 699 3440
rect 733 3406 875 3440
rect 909 3406 1051 3440
rect 1085 3406 1104 3440
rect 279 3388 1104 3406
rect 280 3010 350 3388
rect 680 3010 752 3388
rect 280 2992 752 3010
rect 280 2958 299 2992
rect 333 2958 752 2992
rect 280 2940 752 2958
rect 856 2940 928 3388
rect 1032 2940 1104 3388
rect 2792 3440 3740 3458
rect 2792 3406 2811 3440
rect 2845 3406 2987 3440
rect 3021 3406 3163 3440
rect 3197 3406 3740 3440
rect 2792 3388 3740 3406
rect 2044 3045 2069 3115
rect 2040 2940 2061 3010
rect 2792 2940 2864 3388
rect 2968 2940 3040 3388
rect 3144 3010 3216 3388
rect 3670 3010 3740 3388
rect 3144 2992 3740 3010
rect 3144 2958 3687 2992
rect 3721 2958 3740 2992
rect 3144 2940 3740 2958
rect 592 2877 5311 2906
rect 592 2843 4290 2877
rect 4324 2843 4466 2877
rect 4500 2843 4642 2877
rect 4676 2843 4818 2877
rect 4852 2843 4994 2877
rect 5028 2843 5170 2877
rect 5204 2843 5311 2877
rect 592 2807 5311 2843
rect 592 2775 4378 2807
rect 4269 2773 4378 2775
rect 4412 2773 4554 2807
rect 4588 2773 4730 2807
rect 4764 2773 4906 2807
rect 4940 2773 5082 2807
rect 5116 2773 5258 2807
rect 5292 2773 5311 2807
rect 4269 2755 5311 2773
rect 4130 2703 5531 2721
rect 4130 2702 4290 2703
rect 4130 2668 4149 2702
rect 4183 2669 4290 2702
rect 4324 2669 4466 2703
rect 4500 2669 4642 2703
rect 4676 2669 4818 2703
rect 4852 2669 4994 2703
rect 5028 2669 5170 2703
rect 5204 2669 5367 2703
rect 5401 2669 5531 2703
rect 4183 2668 5531 2669
rect 4130 2651 5531 2668
rect 4130 2650 4343 2651
rect 4284 2544 4330 2591
rect 4284 2510 4290 2544
rect 4324 2510 4330 2544
rect 4284 2472 4330 2510
rect 4284 2438 4290 2472
rect 4324 2438 4330 2472
rect 4284 2400 4330 2438
rect 4284 2366 4290 2400
rect 4324 2366 4330 2400
rect 4284 2328 4330 2366
rect 4284 2294 4290 2328
rect 4324 2294 4330 2328
rect 4284 2256 4330 2294
rect 4284 2222 4290 2256
rect 4324 2222 4330 2256
rect 4284 2184 4330 2222
rect 4284 2150 4290 2184
rect 4324 2150 4330 2184
rect 4284 2112 4330 2150
rect 4284 2078 4290 2112
rect 4324 2078 4330 2112
rect 4284 2040 4330 2078
rect 4284 2006 4290 2040
rect 4324 2006 4330 2040
rect 4284 1968 4330 2006
rect 4284 1934 4290 1968
rect 4324 1934 4330 1968
rect 4284 1896 4330 1934
rect 4284 1862 4290 1896
rect 4324 1862 4330 1896
rect 4284 1824 4330 1862
rect 4284 1790 4290 1824
rect 4324 1790 4330 1824
rect 4284 1752 4330 1790
rect 4284 1718 4290 1752
rect 4324 1718 4330 1752
rect 4284 1680 4330 1718
rect 4284 1646 4290 1680
rect 4324 1646 4330 1680
rect 4284 1608 4330 1646
rect 4284 1574 4290 1608
rect 4324 1574 4330 1608
rect 4284 1536 4330 1574
rect 4284 1502 4290 1536
rect 4324 1502 4330 1536
rect 4284 1464 4330 1502
rect 4284 1430 4290 1464
rect 4324 1430 4330 1464
rect 4284 1392 4330 1430
rect 4284 1358 4290 1392
rect 4324 1358 4330 1392
rect 4284 1320 4330 1358
rect 4284 1286 4290 1320
rect 4324 1286 4330 1320
rect 4284 1248 4330 1286
rect 4284 1214 4290 1248
rect 4324 1214 4330 1248
rect 4284 1176 4330 1214
rect 4284 1142 4290 1176
rect 4324 1142 4330 1176
rect 4284 1104 4330 1142
rect 4284 1070 4290 1104
rect 4324 1070 4330 1104
rect 4284 1032 4330 1070
rect 4284 998 4290 1032
rect 4324 998 4330 1032
rect 4284 960 4330 998
rect 4284 926 4290 960
rect 4324 926 4330 960
rect 4284 888 4330 926
rect 4284 854 4290 888
rect 4324 854 4330 888
rect 4284 816 4330 854
rect 4284 782 4290 816
rect 4324 782 4330 816
rect 4284 744 4330 782
rect 4284 710 4290 744
rect 4324 710 4330 744
rect 4284 672 4330 710
rect 4284 638 4290 672
rect 4324 638 4330 672
rect 4284 591 4330 638
rect 4372 2544 4418 2591
rect 4372 2510 4378 2544
rect 4412 2510 4418 2544
rect 4372 2472 4418 2510
rect 4372 2438 4378 2472
rect 4412 2438 4418 2472
rect 4372 2400 4418 2438
rect 4372 2366 4378 2400
rect 4412 2366 4418 2400
rect 4372 2328 4418 2366
rect 4372 2294 4378 2328
rect 4412 2294 4418 2328
rect 4372 2256 4418 2294
rect 4372 2222 4378 2256
rect 4412 2222 4418 2256
rect 4372 2184 4418 2222
rect 4372 2150 4378 2184
rect 4412 2150 4418 2184
rect 4372 2112 4418 2150
rect 4372 2078 4378 2112
rect 4412 2078 4418 2112
rect 4372 2040 4418 2078
rect 4372 2006 4378 2040
rect 4412 2006 4418 2040
rect 4372 1968 4418 2006
rect 4372 1934 4378 1968
rect 4412 1934 4418 1968
rect 4372 1896 4418 1934
rect 4372 1862 4378 1896
rect 4412 1862 4418 1896
rect 4372 1824 4418 1862
rect 4372 1790 4378 1824
rect 4412 1790 4418 1824
rect 4372 1752 4418 1790
rect 4372 1718 4378 1752
rect 4412 1718 4418 1752
rect 4372 1680 4418 1718
rect 4372 1646 4378 1680
rect 4412 1646 4418 1680
rect 4372 1608 4418 1646
rect 4372 1574 4378 1608
rect 4412 1574 4418 1608
rect 4372 1536 4418 1574
rect 4372 1502 4378 1536
rect 4412 1502 4418 1536
rect 4372 1464 4418 1502
rect 4372 1430 4378 1464
rect 4412 1430 4418 1464
rect 4372 1392 4418 1430
rect 4372 1358 4378 1392
rect 4412 1358 4418 1392
rect 4372 1320 4418 1358
rect 4372 1286 4378 1320
rect 4412 1286 4418 1320
rect 4372 1248 4418 1286
rect 4372 1214 4378 1248
rect 4412 1214 4418 1248
rect 4372 1176 4418 1214
rect 4372 1142 4378 1176
rect 4412 1142 4418 1176
rect 4372 1104 4418 1142
rect 4372 1070 4378 1104
rect 4412 1070 4418 1104
rect 4372 1032 4418 1070
rect 4372 998 4378 1032
rect 4412 998 4418 1032
rect 4372 960 4418 998
rect 4372 926 4378 960
rect 4412 926 4418 960
rect 4372 888 4418 926
rect 4372 854 4378 888
rect 4412 854 4418 888
rect 4372 816 4418 854
rect 4372 782 4378 816
rect 4412 782 4418 816
rect 4372 744 4418 782
rect 4372 710 4378 744
rect 4412 710 4418 744
rect 4372 672 4418 710
rect 4372 638 4378 672
rect 4412 638 4418 672
rect 4372 591 4418 638
rect 4460 2544 4506 2591
rect 4460 2510 4466 2544
rect 4500 2510 4506 2544
rect 4460 2472 4506 2510
rect 4460 2438 4466 2472
rect 4500 2438 4506 2472
rect 4460 2400 4506 2438
rect 4460 2366 4466 2400
rect 4500 2366 4506 2400
rect 4460 2328 4506 2366
rect 4460 2294 4466 2328
rect 4500 2294 4506 2328
rect 4460 2256 4506 2294
rect 4460 2222 4466 2256
rect 4500 2222 4506 2256
rect 4460 2184 4506 2222
rect 4460 2150 4466 2184
rect 4500 2150 4506 2184
rect 4460 2112 4506 2150
rect 4460 2078 4466 2112
rect 4500 2078 4506 2112
rect 4460 2040 4506 2078
rect 4460 2006 4466 2040
rect 4500 2006 4506 2040
rect 4460 1968 4506 2006
rect 4460 1934 4466 1968
rect 4500 1934 4506 1968
rect 4460 1896 4506 1934
rect 4460 1862 4466 1896
rect 4500 1862 4506 1896
rect 4460 1824 4506 1862
rect 4460 1790 4466 1824
rect 4500 1790 4506 1824
rect 4460 1752 4506 1790
rect 4460 1718 4466 1752
rect 4500 1718 4506 1752
rect 4460 1680 4506 1718
rect 4460 1646 4466 1680
rect 4500 1646 4506 1680
rect 4460 1608 4506 1646
rect 4460 1574 4466 1608
rect 4500 1574 4506 1608
rect 4460 1536 4506 1574
rect 4460 1502 4466 1536
rect 4500 1502 4506 1536
rect 4460 1464 4506 1502
rect 4460 1430 4466 1464
rect 4500 1430 4506 1464
rect 4460 1392 4506 1430
rect 4460 1358 4466 1392
rect 4500 1358 4506 1392
rect 4460 1320 4506 1358
rect 4460 1286 4466 1320
rect 4500 1286 4506 1320
rect 4460 1248 4506 1286
rect 4460 1214 4466 1248
rect 4500 1214 4506 1248
rect 4460 1176 4506 1214
rect 4460 1142 4466 1176
rect 4500 1142 4506 1176
rect 4460 1104 4506 1142
rect 4460 1070 4466 1104
rect 4500 1070 4506 1104
rect 4460 1032 4506 1070
rect 4460 998 4466 1032
rect 4500 998 4506 1032
rect 4460 960 4506 998
rect 4460 926 4466 960
rect 4500 926 4506 960
rect 4460 888 4506 926
rect 4460 854 4466 888
rect 4500 854 4506 888
rect 4460 816 4506 854
rect 4460 782 4466 816
rect 4500 782 4506 816
rect 4460 744 4506 782
rect 4460 710 4466 744
rect 4500 710 4506 744
rect 4460 672 4506 710
rect 4460 638 4466 672
rect 4500 638 4506 672
rect 4460 591 4506 638
rect 4548 2544 4594 2591
rect 4548 2510 4554 2544
rect 4588 2510 4594 2544
rect 4548 2472 4594 2510
rect 4548 2438 4554 2472
rect 4588 2438 4594 2472
rect 4548 2400 4594 2438
rect 4548 2366 4554 2400
rect 4588 2366 4594 2400
rect 4548 2328 4594 2366
rect 4548 2294 4554 2328
rect 4588 2294 4594 2328
rect 4548 2256 4594 2294
rect 4548 2222 4554 2256
rect 4588 2222 4594 2256
rect 4548 2184 4594 2222
rect 4548 2150 4554 2184
rect 4588 2150 4594 2184
rect 4548 2112 4594 2150
rect 4548 2078 4554 2112
rect 4588 2078 4594 2112
rect 4548 2040 4594 2078
rect 4548 2006 4554 2040
rect 4588 2006 4594 2040
rect 4548 1968 4594 2006
rect 4548 1934 4554 1968
rect 4588 1934 4594 1968
rect 4548 1896 4594 1934
rect 4548 1862 4554 1896
rect 4588 1862 4594 1896
rect 4548 1824 4594 1862
rect 4548 1790 4554 1824
rect 4588 1790 4594 1824
rect 4548 1752 4594 1790
rect 4548 1718 4554 1752
rect 4588 1718 4594 1752
rect 4548 1680 4594 1718
rect 4548 1646 4554 1680
rect 4588 1646 4594 1680
rect 4548 1608 4594 1646
rect 4548 1574 4554 1608
rect 4588 1574 4594 1608
rect 4548 1536 4594 1574
rect 4548 1502 4554 1536
rect 4588 1502 4594 1536
rect 4548 1464 4594 1502
rect 4548 1430 4554 1464
rect 4588 1430 4594 1464
rect 4548 1392 4594 1430
rect 4548 1358 4554 1392
rect 4588 1358 4594 1392
rect 4548 1320 4594 1358
rect 4548 1286 4554 1320
rect 4588 1286 4594 1320
rect 4548 1248 4594 1286
rect 4548 1214 4554 1248
rect 4588 1214 4594 1248
rect 4548 1176 4594 1214
rect 4548 1142 4554 1176
rect 4588 1142 4594 1176
rect 4548 1104 4594 1142
rect 4548 1070 4554 1104
rect 4588 1070 4594 1104
rect 4548 1032 4594 1070
rect 4548 998 4554 1032
rect 4588 998 4594 1032
rect 4548 960 4594 998
rect 4548 926 4554 960
rect 4588 926 4594 960
rect 4548 888 4594 926
rect 4548 854 4554 888
rect 4588 854 4594 888
rect 4548 816 4594 854
rect 4548 782 4554 816
rect 4588 782 4594 816
rect 4548 744 4594 782
rect 4548 710 4554 744
rect 4588 710 4594 744
rect 4548 672 4594 710
rect 4548 638 4554 672
rect 4588 638 4594 672
rect 4548 591 4594 638
rect 4636 2544 4682 2591
rect 4636 2510 4642 2544
rect 4676 2510 4682 2544
rect 4636 2472 4682 2510
rect 4636 2438 4642 2472
rect 4676 2438 4682 2472
rect 4636 2400 4682 2438
rect 4636 2366 4642 2400
rect 4676 2366 4682 2400
rect 4636 2328 4682 2366
rect 4636 2294 4642 2328
rect 4676 2294 4682 2328
rect 4636 2256 4682 2294
rect 4636 2222 4642 2256
rect 4676 2222 4682 2256
rect 4636 2184 4682 2222
rect 4636 2150 4642 2184
rect 4676 2150 4682 2184
rect 4636 2112 4682 2150
rect 4636 2078 4642 2112
rect 4676 2078 4682 2112
rect 4636 2040 4682 2078
rect 4636 2006 4642 2040
rect 4676 2006 4682 2040
rect 4636 1968 4682 2006
rect 4636 1934 4642 1968
rect 4676 1934 4682 1968
rect 4636 1896 4682 1934
rect 4636 1862 4642 1896
rect 4676 1862 4682 1896
rect 4636 1824 4682 1862
rect 4636 1790 4642 1824
rect 4676 1790 4682 1824
rect 4636 1752 4682 1790
rect 4636 1718 4642 1752
rect 4676 1718 4682 1752
rect 4636 1680 4682 1718
rect 4636 1646 4642 1680
rect 4676 1646 4682 1680
rect 4636 1608 4682 1646
rect 4636 1574 4642 1608
rect 4676 1574 4682 1608
rect 4636 1536 4682 1574
rect 4636 1502 4642 1536
rect 4676 1502 4682 1536
rect 4636 1464 4682 1502
rect 4636 1430 4642 1464
rect 4676 1430 4682 1464
rect 4636 1392 4682 1430
rect 4636 1358 4642 1392
rect 4676 1358 4682 1392
rect 4636 1320 4682 1358
rect 4636 1286 4642 1320
rect 4676 1286 4682 1320
rect 4636 1248 4682 1286
rect 4636 1214 4642 1248
rect 4676 1214 4682 1248
rect 4636 1176 4682 1214
rect 4636 1142 4642 1176
rect 4676 1142 4682 1176
rect 4636 1104 4682 1142
rect 4636 1070 4642 1104
rect 4676 1070 4682 1104
rect 4636 1032 4682 1070
rect 4636 998 4642 1032
rect 4676 998 4682 1032
rect 4636 960 4682 998
rect 4636 926 4642 960
rect 4676 926 4682 960
rect 4636 888 4682 926
rect 4636 854 4642 888
rect 4676 854 4682 888
rect 4636 816 4682 854
rect 4636 782 4642 816
rect 4676 782 4682 816
rect 4636 744 4682 782
rect 4636 710 4642 744
rect 4676 710 4682 744
rect 4636 672 4682 710
rect 4636 638 4642 672
rect 4676 638 4682 672
rect 4636 591 4682 638
rect 4724 2544 4770 2591
rect 4724 2510 4730 2544
rect 4764 2510 4770 2544
rect 4724 2472 4770 2510
rect 4724 2438 4730 2472
rect 4764 2438 4770 2472
rect 4724 2400 4770 2438
rect 4724 2366 4730 2400
rect 4764 2366 4770 2400
rect 4724 2328 4770 2366
rect 4724 2294 4730 2328
rect 4764 2294 4770 2328
rect 4724 2256 4770 2294
rect 4724 2222 4730 2256
rect 4764 2222 4770 2256
rect 4724 2184 4770 2222
rect 4724 2150 4730 2184
rect 4764 2150 4770 2184
rect 4724 2112 4770 2150
rect 4724 2078 4730 2112
rect 4764 2078 4770 2112
rect 4724 2040 4770 2078
rect 4724 2006 4730 2040
rect 4764 2006 4770 2040
rect 4724 1968 4770 2006
rect 4724 1934 4730 1968
rect 4764 1934 4770 1968
rect 4724 1896 4770 1934
rect 4724 1862 4730 1896
rect 4764 1862 4770 1896
rect 4724 1824 4770 1862
rect 4724 1790 4730 1824
rect 4764 1790 4770 1824
rect 4724 1752 4770 1790
rect 4724 1718 4730 1752
rect 4764 1718 4770 1752
rect 4724 1680 4770 1718
rect 4724 1646 4730 1680
rect 4764 1646 4770 1680
rect 4724 1608 4770 1646
rect 4724 1574 4730 1608
rect 4764 1574 4770 1608
rect 4724 1536 4770 1574
rect 4724 1502 4730 1536
rect 4764 1502 4770 1536
rect 4724 1464 4770 1502
rect 4724 1430 4730 1464
rect 4764 1430 4770 1464
rect 4724 1392 4770 1430
rect 4724 1358 4730 1392
rect 4764 1358 4770 1392
rect 4724 1320 4770 1358
rect 4724 1286 4730 1320
rect 4764 1286 4770 1320
rect 4724 1248 4770 1286
rect 4724 1214 4730 1248
rect 4764 1214 4770 1248
rect 4724 1176 4770 1214
rect 4724 1142 4730 1176
rect 4764 1142 4770 1176
rect 4724 1104 4770 1142
rect 4724 1070 4730 1104
rect 4764 1070 4770 1104
rect 4724 1032 4770 1070
rect 4724 998 4730 1032
rect 4764 998 4770 1032
rect 4724 960 4770 998
rect 4724 926 4730 960
rect 4764 926 4770 960
rect 4724 888 4770 926
rect 4724 854 4730 888
rect 4764 854 4770 888
rect 4724 816 4770 854
rect 4724 782 4730 816
rect 4764 782 4770 816
rect 4724 744 4770 782
rect 4724 710 4730 744
rect 4764 710 4770 744
rect 4724 672 4770 710
rect 4724 638 4730 672
rect 4764 638 4770 672
rect 4724 591 4770 638
rect 4812 2544 4858 2591
rect 4812 2510 4818 2544
rect 4852 2510 4858 2544
rect 4812 2472 4858 2510
rect 4812 2438 4818 2472
rect 4852 2438 4858 2472
rect 4812 2400 4858 2438
rect 4812 2366 4818 2400
rect 4852 2366 4858 2400
rect 4812 2328 4858 2366
rect 4812 2294 4818 2328
rect 4852 2294 4858 2328
rect 4812 2256 4858 2294
rect 4812 2222 4818 2256
rect 4852 2222 4858 2256
rect 4812 2184 4858 2222
rect 4812 2150 4818 2184
rect 4852 2150 4858 2184
rect 4812 2112 4858 2150
rect 4812 2078 4818 2112
rect 4852 2078 4858 2112
rect 4812 2040 4858 2078
rect 4812 2006 4818 2040
rect 4852 2006 4858 2040
rect 4812 1968 4858 2006
rect 4812 1934 4818 1968
rect 4852 1934 4858 1968
rect 4812 1896 4858 1934
rect 4812 1862 4818 1896
rect 4852 1862 4858 1896
rect 4812 1824 4858 1862
rect 4812 1790 4818 1824
rect 4852 1790 4858 1824
rect 4812 1752 4858 1790
rect 4812 1718 4818 1752
rect 4852 1718 4858 1752
rect 4812 1680 4858 1718
rect 4812 1646 4818 1680
rect 4852 1646 4858 1680
rect 4812 1608 4858 1646
rect 4812 1574 4818 1608
rect 4852 1574 4858 1608
rect 4812 1536 4858 1574
rect 4812 1502 4818 1536
rect 4852 1502 4858 1536
rect 4812 1464 4858 1502
rect 4812 1430 4818 1464
rect 4852 1430 4858 1464
rect 4812 1392 4858 1430
rect 4812 1358 4818 1392
rect 4852 1358 4858 1392
rect 4812 1320 4858 1358
rect 4812 1286 4818 1320
rect 4852 1286 4858 1320
rect 4812 1248 4858 1286
rect 4812 1214 4818 1248
rect 4852 1214 4858 1248
rect 4812 1176 4858 1214
rect 4812 1142 4818 1176
rect 4852 1142 4858 1176
rect 4812 1104 4858 1142
rect 4812 1070 4818 1104
rect 4852 1070 4858 1104
rect 4812 1032 4858 1070
rect 4812 998 4818 1032
rect 4852 998 4858 1032
rect 4812 960 4858 998
rect 4812 926 4818 960
rect 4852 926 4858 960
rect 4812 888 4858 926
rect 4812 854 4818 888
rect 4852 854 4858 888
rect 4812 816 4858 854
rect 4812 782 4818 816
rect 4852 782 4858 816
rect 4812 744 4858 782
rect 4812 710 4818 744
rect 4852 710 4858 744
rect 4812 672 4858 710
rect 4812 638 4818 672
rect 4852 638 4858 672
rect 4812 591 4858 638
rect 4900 2544 4946 2591
rect 4900 2510 4906 2544
rect 4940 2510 4946 2544
rect 4900 2472 4946 2510
rect 4900 2438 4906 2472
rect 4940 2438 4946 2472
rect 4900 2400 4946 2438
rect 4900 2366 4906 2400
rect 4940 2366 4946 2400
rect 4900 2328 4946 2366
rect 4900 2294 4906 2328
rect 4940 2294 4946 2328
rect 4900 2256 4946 2294
rect 4900 2222 4906 2256
rect 4940 2222 4946 2256
rect 4900 2184 4946 2222
rect 4900 2150 4906 2184
rect 4940 2150 4946 2184
rect 4900 2112 4946 2150
rect 4900 2078 4906 2112
rect 4940 2078 4946 2112
rect 4900 2040 4946 2078
rect 4900 2006 4906 2040
rect 4940 2006 4946 2040
rect 4900 1968 4946 2006
rect 4900 1934 4906 1968
rect 4940 1934 4946 1968
rect 4900 1896 4946 1934
rect 4900 1862 4906 1896
rect 4940 1862 4946 1896
rect 4900 1824 4946 1862
rect 4900 1790 4906 1824
rect 4940 1790 4946 1824
rect 4900 1752 4946 1790
rect 4900 1718 4906 1752
rect 4940 1718 4946 1752
rect 4900 1680 4946 1718
rect 4900 1646 4906 1680
rect 4940 1646 4946 1680
rect 4900 1608 4946 1646
rect 4900 1574 4906 1608
rect 4940 1574 4946 1608
rect 4900 1536 4946 1574
rect 4900 1502 4906 1536
rect 4940 1502 4946 1536
rect 4900 1464 4946 1502
rect 4900 1430 4906 1464
rect 4940 1430 4946 1464
rect 4900 1392 4946 1430
rect 4900 1358 4906 1392
rect 4940 1358 4946 1392
rect 4900 1320 4946 1358
rect 4900 1286 4906 1320
rect 4940 1286 4946 1320
rect 4900 1248 4946 1286
rect 4900 1214 4906 1248
rect 4940 1214 4946 1248
rect 4900 1176 4946 1214
rect 4900 1142 4906 1176
rect 4940 1142 4946 1176
rect 4900 1104 4946 1142
rect 4900 1070 4906 1104
rect 4940 1070 4946 1104
rect 4900 1032 4946 1070
rect 4900 998 4906 1032
rect 4940 998 4946 1032
rect 4900 960 4946 998
rect 4900 926 4906 960
rect 4940 926 4946 960
rect 4900 888 4946 926
rect 4900 854 4906 888
rect 4940 854 4946 888
rect 4900 816 4946 854
rect 4900 782 4906 816
rect 4940 782 4946 816
rect 4900 744 4946 782
rect 4900 710 4906 744
rect 4940 710 4946 744
rect 4900 672 4946 710
rect 4900 638 4906 672
rect 4940 638 4946 672
rect 4900 591 4946 638
rect 4988 2544 5034 2591
rect 4988 2510 4994 2544
rect 5028 2510 5034 2544
rect 4988 2472 5034 2510
rect 4988 2438 4994 2472
rect 5028 2438 5034 2472
rect 4988 2400 5034 2438
rect 4988 2366 4994 2400
rect 5028 2366 5034 2400
rect 4988 2328 5034 2366
rect 4988 2294 4994 2328
rect 5028 2294 5034 2328
rect 4988 2256 5034 2294
rect 4988 2222 4994 2256
rect 5028 2222 5034 2256
rect 4988 2184 5034 2222
rect 4988 2150 4994 2184
rect 5028 2150 5034 2184
rect 4988 2112 5034 2150
rect 4988 2078 4994 2112
rect 5028 2078 5034 2112
rect 4988 2040 5034 2078
rect 4988 2006 4994 2040
rect 5028 2006 5034 2040
rect 4988 1968 5034 2006
rect 4988 1934 4994 1968
rect 5028 1934 5034 1968
rect 4988 1896 5034 1934
rect 4988 1862 4994 1896
rect 5028 1862 5034 1896
rect 4988 1824 5034 1862
rect 4988 1790 4994 1824
rect 5028 1790 5034 1824
rect 4988 1752 5034 1790
rect 4988 1718 4994 1752
rect 5028 1718 5034 1752
rect 4988 1680 5034 1718
rect 4988 1646 4994 1680
rect 5028 1646 5034 1680
rect 4988 1608 5034 1646
rect 4988 1574 4994 1608
rect 5028 1574 5034 1608
rect 4988 1536 5034 1574
rect 4988 1502 4994 1536
rect 5028 1502 5034 1536
rect 4988 1464 5034 1502
rect 4988 1430 4994 1464
rect 5028 1430 5034 1464
rect 4988 1392 5034 1430
rect 4988 1358 4994 1392
rect 5028 1358 5034 1392
rect 4988 1320 5034 1358
rect 4988 1286 4994 1320
rect 5028 1286 5034 1320
rect 4988 1248 5034 1286
rect 4988 1214 4994 1248
rect 5028 1214 5034 1248
rect 4988 1176 5034 1214
rect 4988 1142 4994 1176
rect 5028 1142 5034 1176
rect 4988 1104 5034 1142
rect 4988 1070 4994 1104
rect 5028 1070 5034 1104
rect 4988 1032 5034 1070
rect 4988 998 4994 1032
rect 5028 998 5034 1032
rect 4988 960 5034 998
rect 4988 926 4994 960
rect 5028 926 5034 960
rect 4988 888 5034 926
rect 4988 854 4994 888
rect 5028 854 5034 888
rect 4988 816 5034 854
rect 4988 782 4994 816
rect 5028 782 5034 816
rect 4988 744 5034 782
rect 4988 710 4994 744
rect 5028 710 5034 744
rect 4988 672 5034 710
rect 4988 638 4994 672
rect 5028 638 5034 672
rect 4988 591 5034 638
rect 5076 2544 5122 2591
rect 5076 2510 5082 2544
rect 5116 2510 5122 2544
rect 5076 2472 5122 2510
rect 5076 2438 5082 2472
rect 5116 2438 5122 2472
rect 5076 2400 5122 2438
rect 5076 2366 5082 2400
rect 5116 2366 5122 2400
rect 5076 2328 5122 2366
rect 5076 2294 5082 2328
rect 5116 2294 5122 2328
rect 5076 2256 5122 2294
rect 5076 2222 5082 2256
rect 5116 2222 5122 2256
rect 5076 2184 5122 2222
rect 5076 2150 5082 2184
rect 5116 2150 5122 2184
rect 5076 2112 5122 2150
rect 5076 2078 5082 2112
rect 5116 2078 5122 2112
rect 5076 2040 5122 2078
rect 5076 2006 5082 2040
rect 5116 2006 5122 2040
rect 5076 1968 5122 2006
rect 5076 1934 5082 1968
rect 5116 1934 5122 1968
rect 5076 1896 5122 1934
rect 5076 1862 5082 1896
rect 5116 1862 5122 1896
rect 5076 1824 5122 1862
rect 5076 1790 5082 1824
rect 5116 1790 5122 1824
rect 5076 1752 5122 1790
rect 5076 1718 5082 1752
rect 5116 1718 5122 1752
rect 5076 1680 5122 1718
rect 5076 1646 5082 1680
rect 5116 1646 5122 1680
rect 5076 1608 5122 1646
rect 5076 1574 5082 1608
rect 5116 1574 5122 1608
rect 5076 1536 5122 1574
rect 5076 1502 5082 1536
rect 5116 1502 5122 1536
rect 5076 1464 5122 1502
rect 5076 1430 5082 1464
rect 5116 1430 5122 1464
rect 5076 1392 5122 1430
rect 5076 1358 5082 1392
rect 5116 1358 5122 1392
rect 5076 1320 5122 1358
rect 5076 1286 5082 1320
rect 5116 1286 5122 1320
rect 5076 1248 5122 1286
rect 5076 1214 5082 1248
rect 5116 1214 5122 1248
rect 5076 1176 5122 1214
rect 5076 1142 5082 1176
rect 5116 1142 5122 1176
rect 5076 1104 5122 1142
rect 5076 1070 5082 1104
rect 5116 1070 5122 1104
rect 5076 1032 5122 1070
rect 5076 998 5082 1032
rect 5116 998 5122 1032
rect 5076 960 5122 998
rect 5076 926 5082 960
rect 5116 926 5122 960
rect 5076 888 5122 926
rect 5076 854 5082 888
rect 5116 854 5122 888
rect 5076 816 5122 854
rect 5076 782 5082 816
rect 5116 782 5122 816
rect 5076 744 5122 782
rect 5076 710 5082 744
rect 5116 710 5122 744
rect 5076 672 5122 710
rect 5076 638 5082 672
rect 5116 638 5122 672
rect 5076 591 5122 638
rect 5164 2544 5210 2591
rect 5164 2510 5170 2544
rect 5204 2510 5210 2544
rect 5164 2472 5210 2510
rect 5164 2438 5170 2472
rect 5204 2438 5210 2472
rect 5164 2400 5210 2438
rect 5164 2366 5170 2400
rect 5204 2366 5210 2400
rect 5164 2328 5210 2366
rect 5164 2294 5170 2328
rect 5204 2294 5210 2328
rect 5164 2256 5210 2294
rect 5164 2222 5170 2256
rect 5204 2222 5210 2256
rect 5164 2184 5210 2222
rect 5164 2150 5170 2184
rect 5204 2150 5210 2184
rect 5164 2112 5210 2150
rect 5164 2078 5170 2112
rect 5204 2078 5210 2112
rect 5164 2040 5210 2078
rect 5164 2006 5170 2040
rect 5204 2006 5210 2040
rect 5164 1968 5210 2006
rect 5164 1934 5170 1968
rect 5204 1934 5210 1968
rect 5164 1896 5210 1934
rect 5164 1862 5170 1896
rect 5204 1862 5210 1896
rect 5164 1824 5210 1862
rect 5164 1790 5170 1824
rect 5204 1790 5210 1824
rect 5164 1752 5210 1790
rect 5164 1718 5170 1752
rect 5204 1718 5210 1752
rect 5164 1680 5210 1718
rect 5164 1646 5170 1680
rect 5204 1646 5210 1680
rect 5164 1608 5210 1646
rect 5164 1574 5170 1608
rect 5204 1574 5210 1608
rect 5164 1536 5210 1574
rect 5164 1502 5170 1536
rect 5204 1502 5210 1536
rect 5164 1464 5210 1502
rect 5164 1430 5170 1464
rect 5204 1430 5210 1464
rect 5164 1392 5210 1430
rect 5164 1358 5170 1392
rect 5204 1358 5210 1392
rect 5164 1320 5210 1358
rect 5164 1286 5170 1320
rect 5204 1286 5210 1320
rect 5164 1248 5210 1286
rect 5164 1214 5170 1248
rect 5204 1214 5210 1248
rect 5164 1176 5210 1214
rect 5164 1142 5170 1176
rect 5204 1142 5210 1176
rect 5164 1104 5210 1142
rect 5164 1070 5170 1104
rect 5204 1070 5210 1104
rect 5164 1032 5210 1070
rect 5164 998 5170 1032
rect 5204 998 5210 1032
rect 5164 960 5210 998
rect 5164 926 5170 960
rect 5204 926 5210 960
rect 5164 888 5210 926
rect 5164 854 5170 888
rect 5204 854 5210 888
rect 5164 816 5210 854
rect 5164 782 5170 816
rect 5204 782 5210 816
rect 5164 744 5210 782
rect 5164 710 5170 744
rect 5204 710 5210 744
rect 5164 672 5210 710
rect 5164 638 5170 672
rect 5204 638 5210 672
rect 5164 591 5210 638
rect 5252 2544 5298 2591
rect 5252 2510 5258 2544
rect 5292 2510 5298 2544
rect 5252 2472 5298 2510
rect 5252 2438 5258 2472
rect 5292 2438 5298 2472
rect 5252 2400 5298 2438
rect 5252 2366 5258 2400
rect 5292 2366 5298 2400
rect 5252 2328 5298 2366
rect 5252 2294 5258 2328
rect 5292 2294 5298 2328
rect 5252 2256 5298 2294
rect 5252 2222 5258 2256
rect 5292 2222 5298 2256
rect 5252 2184 5298 2222
rect 5252 2150 5258 2184
rect 5292 2150 5298 2184
rect 5252 2112 5298 2150
rect 5252 2078 5258 2112
rect 5292 2078 5298 2112
rect 5252 2040 5298 2078
rect 5252 2006 5258 2040
rect 5292 2006 5298 2040
rect 5252 1968 5298 2006
rect 5252 1934 5258 1968
rect 5292 1934 5298 1968
rect 5252 1896 5298 1934
rect 5252 1862 5258 1896
rect 5292 1862 5298 1896
rect 5252 1824 5298 1862
rect 5252 1790 5258 1824
rect 5292 1790 5298 1824
rect 5252 1752 5298 1790
rect 5252 1718 5258 1752
rect 5292 1718 5298 1752
rect 5252 1680 5298 1718
rect 5252 1646 5258 1680
rect 5292 1646 5298 1680
rect 5252 1608 5298 1646
rect 5252 1574 5258 1608
rect 5292 1574 5298 1608
rect 5252 1536 5298 1574
rect 5252 1502 5258 1536
rect 5292 1502 5298 1536
rect 5252 1464 5298 1502
rect 5252 1430 5258 1464
rect 5292 1430 5298 1464
rect 5252 1392 5298 1430
rect 5252 1358 5258 1392
rect 5292 1358 5298 1392
rect 5252 1320 5298 1358
rect 5252 1286 5258 1320
rect 5292 1286 5298 1320
rect 5252 1248 5298 1286
rect 5252 1214 5258 1248
rect 5292 1214 5298 1248
rect 5252 1176 5298 1214
rect 5252 1142 5258 1176
rect 5292 1142 5298 1176
rect 5252 1104 5298 1142
rect 5252 1070 5258 1104
rect 5292 1070 5298 1104
rect 5252 1032 5298 1070
rect 5252 998 5258 1032
rect 5292 998 5298 1032
rect 5252 960 5298 998
rect 5252 926 5258 960
rect 5292 926 5298 960
rect 5252 888 5298 926
rect 5252 854 5258 888
rect 5292 854 5298 888
rect 5252 816 5298 854
rect 5252 782 5258 816
rect 5292 782 5298 816
rect 5252 744 5298 782
rect 5252 710 5258 744
rect 5292 710 5298 744
rect 5252 672 5298 710
rect 5252 638 5258 672
rect 5292 638 5298 672
rect 5252 591 5298 638
rect 1943 418 1966 555
rect 2911 553 4802 555
rect 2911 509 5159 553
rect 2911 475 4378 509
rect 4412 475 4554 509
rect 4588 475 4730 509
rect 4764 475 4906 509
rect 4940 475 5082 509
rect 5116 475 5159 509
rect 2911 418 5159 475
use cascode  cascode_0
timestamp 1636132012
transform 1 0 599 0 1 719
box -773 -653 3221 2834
<< labels >>
rlabel metal1 s 2055 3115 2055 3115 4 D2
port 1 nsew
rlabel metal1 s 2049 3010 2049 3010 4 S1
port 2 nsew
rlabel metal1 s 1955 418 1955 418 4 G1
port 3 nsew
rlabel metal1 s 5531 2671 5531 2671 4 VDD
port 4 nsew
<< end >>
