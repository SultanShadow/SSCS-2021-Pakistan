magic
tech sky130A
magscale 1 2
timestamp 1635855079
<< metal4 >>
rect -3351 2518 3351 2600
rect -3351 2282 3095 2518
rect 3331 2282 3351 2518
rect -3351 2198 3351 2282
rect -3351 1962 3095 2198
rect 3331 1962 3351 2198
rect -3351 1878 3351 1962
rect -3351 1642 3095 1878
rect 3331 1642 3351 1878
rect -3351 1558 3351 1642
rect -3351 1322 3095 1558
rect 3331 1322 3351 1558
rect -3351 1238 3351 1322
rect -3351 1002 3095 1238
rect 3331 1002 3351 1238
rect -3351 918 3351 1002
rect -3351 682 3095 918
rect 3331 682 3351 918
rect -3351 598 3351 682
rect -3351 362 3095 598
rect 3331 362 3351 598
rect -3351 278 3351 362
rect -3351 42 3095 278
rect 3331 42 3351 278
rect -3351 -42 3351 42
rect -3351 -278 3095 -42
rect 3331 -278 3351 -42
rect -3351 -362 3351 -278
rect -3351 -598 3095 -362
rect 3331 -598 3351 -362
rect -3351 -682 3351 -598
rect -3351 -918 3095 -682
rect 3331 -918 3351 -682
rect -3351 -1002 3351 -918
rect -3351 -1238 3095 -1002
rect 3331 -1238 3351 -1002
rect -3351 -1322 3351 -1238
rect -3351 -1558 3095 -1322
rect 3331 -1558 3351 -1322
rect -3351 -1642 3351 -1558
rect -3351 -1878 3095 -1642
rect 3331 -1878 3351 -1642
rect -3351 -1962 3351 -1878
rect -3351 -2198 3095 -1962
rect 3331 -2198 3351 -1962
rect -3351 -2282 3351 -2198
rect -3351 -2518 3095 -2282
rect 3331 -2518 3351 -2282
rect -3351 -2600 3351 -2518
<< via4 >>
rect 3095 2282 3331 2518
rect 3095 1962 3331 2198
rect 3095 1642 3331 1878
rect 3095 1322 3331 1558
rect 3095 1002 3331 1238
rect 3095 682 3331 918
rect 3095 362 3331 598
rect 3095 42 3331 278
rect 3095 -278 3331 -42
rect 3095 -598 3331 -362
rect 3095 -918 3331 -682
rect 3095 -1238 3331 -1002
rect 3095 -1558 3331 -1322
rect 3095 -1878 3331 -1642
rect 3095 -2198 3331 -1962
rect 3095 -2518 3331 -2282
<< mimcap2 >>
rect -3251 2358 2749 2500
rect -3251 -2358 -3089 2358
rect 2587 -2358 2749 2358
rect -3251 -2500 2749 -2358
<< mimcap2contact >>
rect -3089 -2358 2587 2358
<< metal5 >>
rect 3053 2518 3373 2601
rect -3235 2358 2733 2484
rect -3235 -2358 -3089 2358
rect 2587 -2358 2733 2358
rect -3235 -2484 2733 -2358
rect 3053 2282 3095 2518
rect 3331 2282 3373 2518
rect 3053 2198 3373 2282
rect 3053 1962 3095 2198
rect 3331 1962 3373 2198
rect 3053 1878 3373 1962
rect 3053 1642 3095 1878
rect 3331 1642 3373 1878
rect 3053 1558 3373 1642
rect 3053 1322 3095 1558
rect 3331 1322 3373 1558
rect 3053 1238 3373 1322
rect 3053 1002 3095 1238
rect 3331 1002 3373 1238
rect 3053 918 3373 1002
rect 3053 682 3095 918
rect 3331 682 3373 918
rect 3053 598 3373 682
rect 3053 362 3095 598
rect 3331 362 3373 598
rect 3053 278 3373 362
rect 3053 42 3095 278
rect 3331 42 3373 278
rect 3053 -42 3373 42
rect 3053 -278 3095 -42
rect 3331 -278 3373 -42
rect 3053 -362 3373 -278
rect 3053 -598 3095 -362
rect 3331 -598 3373 -362
rect 3053 -682 3373 -598
rect 3053 -918 3095 -682
rect 3331 -918 3373 -682
rect 3053 -1002 3373 -918
rect 3053 -1238 3095 -1002
rect 3331 -1238 3373 -1002
rect 3053 -1322 3373 -1238
rect 3053 -1558 3095 -1322
rect 3331 -1558 3373 -1322
rect 3053 -1642 3373 -1558
rect 3053 -1878 3095 -1642
rect 3331 -1878 3373 -1642
rect 3053 -1962 3373 -1878
rect 3053 -2198 3095 -1962
rect 3331 -2198 3373 -1962
rect 3053 -2282 3373 -2198
rect 3053 -2518 3095 -2282
rect 3331 -2518 3373 -2282
rect 3053 -2601 3373 -2518
<< properties >>
string FIXED_BBOX -3351 -2600 2849 2600
<< end >>
