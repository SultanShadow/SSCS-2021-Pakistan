magic
tech sky130A
magscale 1 2
timestamp 1637060811
<< metal4 >>
rect -1851 1558 1851 1600
rect -1851 1322 1595 1558
rect 1831 1322 1851 1558
rect -1851 1238 1851 1322
rect -1851 1002 1595 1238
rect 1831 1002 1851 1238
rect -1851 918 1851 1002
rect -1851 682 1595 918
rect 1831 682 1851 918
rect -1851 598 1851 682
rect -1851 362 1595 598
rect 1831 362 1851 598
rect -1851 278 1851 362
rect -1851 42 1595 278
rect 1831 42 1851 278
rect -1851 -42 1851 42
rect -1851 -278 1595 -42
rect 1831 -278 1851 -42
rect -1851 -362 1851 -278
rect -1851 -598 1595 -362
rect 1831 -598 1851 -362
rect -1851 -682 1851 -598
rect -1851 -918 1595 -682
rect 1831 -918 1851 -682
rect -1851 -1002 1851 -918
rect -1851 -1238 1595 -1002
rect 1831 -1238 1851 -1002
rect -1851 -1322 1851 -1238
rect -1851 -1558 1595 -1322
rect 1831 -1558 1851 -1322
rect -1851 -1600 1851 -1558
<< via4 >>
rect 1595 1322 1831 1558
rect 1595 1002 1831 1238
rect 1595 682 1831 918
rect 1595 362 1831 598
rect 1595 42 1831 278
rect 1595 -278 1831 -42
rect 1595 -598 1831 -362
rect 1595 -918 1831 -682
rect 1595 -1238 1831 -1002
rect 1595 -1558 1831 -1322
<< mimcap2 >>
rect -1751 1398 1249 1500
rect -1751 -1398 -1649 1398
rect 1147 -1398 1249 1398
rect -1751 -1500 1249 -1398
<< mimcap2contact >>
rect -1649 -1398 1147 1398
<< metal5 >>
rect 1553 1558 1873 1601
rect -1735 1398 1233 1484
rect -1735 -1398 -1649 1398
rect 1147 -1398 1233 1398
rect -1735 -1484 1233 -1398
rect 1553 1322 1595 1558
rect 1831 1322 1873 1558
rect 1553 1238 1873 1322
rect 1553 1002 1595 1238
rect 1831 1002 1873 1238
rect 1553 918 1873 1002
rect 1553 682 1595 918
rect 1831 682 1873 918
rect 1553 598 1873 682
rect 1553 362 1595 598
rect 1831 362 1873 598
rect 1553 278 1873 362
rect 1553 42 1595 278
rect 1831 42 1873 278
rect 1553 -42 1873 42
rect 1553 -278 1595 -42
rect 1831 -278 1873 -42
rect 1553 -362 1873 -278
rect 1553 -598 1595 -362
rect 1831 -598 1873 -362
rect 1553 -682 1873 -598
rect 1553 -918 1595 -682
rect 1831 -918 1873 -682
rect 1553 -1002 1873 -918
rect 1553 -1238 1595 -1002
rect 1831 -1238 1873 -1002
rect 1553 -1322 1873 -1238
rect 1553 -1558 1595 -1322
rect 1831 -1558 1873 -1322
rect 1553 -1601 1873 -1558
<< properties >>
string FIXED_BBOX -1851 -1600 1349 1600
<< end >>
