magic
tech sky130A
magscale 1 2
timestamp 1637060811
<< error_p >>
rect -73 -600 -15 600
rect 15 -600 73 600
<< pwell >>
rect -99 -626 99 626
<< nmoslvt >>
rect -15 -600 15 600
<< ndiff >>
rect -73 561 -15 600
rect -73 527 -61 561
rect -27 527 -15 561
rect -73 493 -15 527
rect -73 459 -61 493
rect -27 459 -15 493
rect -73 425 -15 459
rect -73 391 -61 425
rect -27 391 -15 425
rect -73 357 -15 391
rect -73 323 -61 357
rect -27 323 -15 357
rect -73 289 -15 323
rect -73 255 -61 289
rect -27 255 -15 289
rect -73 221 -15 255
rect -73 187 -61 221
rect -27 187 -15 221
rect -73 153 -15 187
rect -73 119 -61 153
rect -27 119 -15 153
rect -73 85 -15 119
rect -73 51 -61 85
rect -27 51 -15 85
rect -73 17 -15 51
rect -73 -17 -61 17
rect -27 -17 -15 17
rect -73 -51 -15 -17
rect -73 -85 -61 -51
rect -27 -85 -15 -51
rect -73 -119 -15 -85
rect -73 -153 -61 -119
rect -27 -153 -15 -119
rect -73 -187 -15 -153
rect -73 -221 -61 -187
rect -27 -221 -15 -187
rect -73 -255 -15 -221
rect -73 -289 -61 -255
rect -27 -289 -15 -255
rect -73 -323 -15 -289
rect -73 -357 -61 -323
rect -27 -357 -15 -323
rect -73 -391 -15 -357
rect -73 -425 -61 -391
rect -27 -425 -15 -391
rect -73 -459 -15 -425
rect -73 -493 -61 -459
rect -27 -493 -15 -459
rect -73 -527 -15 -493
rect -73 -561 -61 -527
rect -27 -561 -15 -527
rect -73 -600 -15 -561
rect 15 561 73 600
rect 15 527 27 561
rect 61 527 73 561
rect 15 493 73 527
rect 15 459 27 493
rect 61 459 73 493
rect 15 425 73 459
rect 15 391 27 425
rect 61 391 73 425
rect 15 357 73 391
rect 15 323 27 357
rect 61 323 73 357
rect 15 289 73 323
rect 15 255 27 289
rect 61 255 73 289
rect 15 221 73 255
rect 15 187 27 221
rect 61 187 73 221
rect 15 153 73 187
rect 15 119 27 153
rect 61 119 73 153
rect 15 85 73 119
rect 15 51 27 85
rect 61 51 73 85
rect 15 17 73 51
rect 15 -17 27 17
rect 61 -17 73 17
rect 15 -51 73 -17
rect 15 -85 27 -51
rect 61 -85 73 -51
rect 15 -119 73 -85
rect 15 -153 27 -119
rect 61 -153 73 -119
rect 15 -187 73 -153
rect 15 -221 27 -187
rect 61 -221 73 -187
rect 15 -255 73 -221
rect 15 -289 27 -255
rect 61 -289 73 -255
rect 15 -323 73 -289
rect 15 -357 27 -323
rect 61 -357 73 -323
rect 15 -391 73 -357
rect 15 -425 27 -391
rect 61 -425 73 -391
rect 15 -459 73 -425
rect 15 -493 27 -459
rect 61 -493 73 -459
rect 15 -527 73 -493
rect 15 -561 27 -527
rect 61 -561 73 -527
rect 15 -600 73 -561
<< ndiffc >>
rect -61 527 -27 561
rect -61 459 -27 493
rect -61 391 -27 425
rect -61 323 -27 357
rect -61 255 -27 289
rect -61 187 -27 221
rect -61 119 -27 153
rect -61 51 -27 85
rect -61 -17 -27 17
rect -61 -85 -27 -51
rect -61 -153 -27 -119
rect -61 -221 -27 -187
rect -61 -289 -27 -255
rect -61 -357 -27 -323
rect -61 -425 -27 -391
rect -61 -493 -27 -459
rect -61 -561 -27 -527
rect 27 527 61 561
rect 27 459 61 493
rect 27 391 61 425
rect 27 323 61 357
rect 27 255 61 289
rect 27 187 61 221
rect 27 119 61 153
rect 27 51 61 85
rect 27 -17 61 17
rect 27 -85 61 -51
rect 27 -153 61 -119
rect 27 -221 61 -187
rect 27 -289 61 -255
rect 27 -357 61 -323
rect 27 -425 61 -391
rect 27 -493 61 -459
rect 27 -561 61 -527
<< poly >>
rect -15 600 15 626
rect -15 -626 15 -600
<< locali >>
rect -61 561 -27 604
rect -61 493 -27 523
rect -61 425 -27 451
rect -61 357 -27 379
rect -61 289 -27 307
rect -61 221 -27 235
rect -61 153 -27 163
rect -61 85 -27 91
rect -61 17 -27 19
rect -61 -19 -27 -17
rect -61 -91 -27 -85
rect -61 -163 -27 -153
rect -61 -235 -27 -221
rect -61 -307 -27 -289
rect -61 -379 -27 -357
rect -61 -451 -27 -425
rect -61 -523 -27 -493
rect -61 -604 -27 -561
rect 27 561 61 604
rect 27 493 61 523
rect 27 425 61 451
rect 27 357 61 379
rect 27 289 61 307
rect 27 221 61 235
rect 27 153 61 163
rect 27 85 61 91
rect 27 17 61 19
rect 27 -19 61 -17
rect 27 -91 61 -85
rect 27 -163 61 -153
rect 27 -235 61 -221
rect 27 -307 61 -289
rect 27 -379 61 -357
rect 27 -451 61 -425
rect 27 -523 61 -493
rect 27 -604 61 -561
<< viali >>
rect -61 527 -27 557
rect -61 523 -27 527
rect -61 459 -27 485
rect -61 451 -27 459
rect -61 391 -27 413
rect -61 379 -27 391
rect -61 323 -27 341
rect -61 307 -27 323
rect -61 255 -27 269
rect -61 235 -27 255
rect -61 187 -27 197
rect -61 163 -27 187
rect -61 119 -27 125
rect -61 91 -27 119
rect -61 51 -27 53
rect -61 19 -27 51
rect -61 -51 -27 -19
rect -61 -53 -27 -51
rect -61 -119 -27 -91
rect -61 -125 -27 -119
rect -61 -187 -27 -163
rect -61 -197 -27 -187
rect -61 -255 -27 -235
rect -61 -269 -27 -255
rect -61 -323 -27 -307
rect -61 -341 -27 -323
rect -61 -391 -27 -379
rect -61 -413 -27 -391
rect -61 -459 -27 -451
rect -61 -485 -27 -459
rect -61 -527 -27 -523
rect -61 -557 -27 -527
rect 27 527 61 557
rect 27 523 61 527
rect 27 459 61 485
rect 27 451 61 459
rect 27 391 61 413
rect 27 379 61 391
rect 27 323 61 341
rect 27 307 61 323
rect 27 255 61 269
rect 27 235 61 255
rect 27 187 61 197
rect 27 163 61 187
rect 27 119 61 125
rect 27 91 61 119
rect 27 51 61 53
rect 27 19 61 51
rect 27 -51 61 -19
rect 27 -53 61 -51
rect 27 -119 61 -91
rect 27 -125 61 -119
rect 27 -187 61 -163
rect 27 -197 61 -187
rect 27 -255 61 -235
rect 27 -269 61 -255
rect 27 -323 61 -307
rect 27 -341 61 -323
rect 27 -391 61 -379
rect 27 -413 61 -391
rect 27 -459 61 -451
rect 27 -485 61 -459
rect 27 -527 61 -523
rect 27 -557 61 -527
<< metal1 >>
rect -67 557 -21 600
rect -67 523 -61 557
rect -27 523 -21 557
rect -67 485 -21 523
rect -67 451 -61 485
rect -27 451 -21 485
rect -67 413 -21 451
rect -67 379 -61 413
rect -27 379 -21 413
rect -67 341 -21 379
rect -67 307 -61 341
rect -27 307 -21 341
rect -67 269 -21 307
rect -67 235 -61 269
rect -27 235 -21 269
rect -67 197 -21 235
rect -67 163 -61 197
rect -27 163 -21 197
rect -67 125 -21 163
rect -67 91 -61 125
rect -27 91 -21 125
rect -67 53 -21 91
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -91 -21 -53
rect -67 -125 -61 -91
rect -27 -125 -21 -91
rect -67 -163 -21 -125
rect -67 -197 -61 -163
rect -27 -197 -21 -163
rect -67 -235 -21 -197
rect -67 -269 -61 -235
rect -27 -269 -21 -235
rect -67 -307 -21 -269
rect -67 -341 -61 -307
rect -27 -341 -21 -307
rect -67 -379 -21 -341
rect -67 -413 -61 -379
rect -27 -413 -21 -379
rect -67 -451 -21 -413
rect -67 -485 -61 -451
rect -27 -485 -21 -451
rect -67 -523 -21 -485
rect -67 -557 -61 -523
rect -27 -557 -21 -523
rect -67 -600 -21 -557
rect 21 557 67 600
rect 21 523 27 557
rect 61 523 67 557
rect 21 485 67 523
rect 21 451 27 485
rect 61 451 67 485
rect 21 413 67 451
rect 21 379 27 413
rect 61 379 67 413
rect 21 341 67 379
rect 21 307 27 341
rect 61 307 67 341
rect 21 269 67 307
rect 21 235 27 269
rect 61 235 67 269
rect 21 197 67 235
rect 21 163 27 197
rect 61 163 67 197
rect 21 125 67 163
rect 21 91 27 125
rect 61 91 67 125
rect 21 53 67 91
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -91 67 -53
rect 21 -125 27 -91
rect 61 -125 67 -91
rect 21 -163 67 -125
rect 21 -197 27 -163
rect 61 -197 67 -163
rect 21 -235 67 -197
rect 21 -269 27 -235
rect 61 -269 67 -235
rect 21 -307 67 -269
rect 21 -341 27 -307
rect 61 -341 67 -307
rect 21 -379 67 -341
rect 21 -413 27 -379
rect 61 -413 67 -379
rect 21 -451 67 -413
rect 21 -485 27 -451
rect 61 -485 67 -451
rect 21 -523 67 -485
rect 21 -557 27 -523
rect 61 -557 67 -523
rect 21 -600 67 -557
<< end >>
