magic
tech sky130A
magscale 1 2
timestamp 1635855079
<< metal3 >>
rect -90032 -88468 7414 6314
rect -90032 -88800 7438 -88468
rect -83242 -89592 7438 -88800
<< metal4 >>
rect -85808 7468 4410 8920
rect -85790 -85968 -84576 7468
rect -79572 -85738 -78358 7468
rect -73126 -86058 -71912 7468
rect -66720 -85938 -65506 7468
rect -60354 -86138 -59140 7468
rect -54270 -86258 -53056 7468
rect -47904 -86098 -46690 7468
rect -41378 -85978 -40164 7468
rect -35174 -85818 -33960 7468
rect -28768 -85698 -27554 7468
rect -22762 -85538 -21548 7468
rect -16518 -85578 -15304 7468
rect -10112 -85338 -8898 7468
rect -3466 -85218 -2252 7468
rect 2660 -85218 3874 7468
rect -82316 -88468 -82128 -88080
rect -76018 -88468 -75830 -88170
rect -69672 -88468 -69484 -88164
rect -63366 -88468 -63178 -88160
rect -57032 -88468 -56844 -88092
rect -50696 -88468 -50508 -88118
rect -44378 -88468 -44190 -88108
rect -38092 -88468 -37904 -88046
rect -31770 -88468 -31582 -88186
rect -25416 -88468 -25228 -88068
rect -19096 -88468 -18908 -88056
rect -12792 -88468 -12604 -87990
rect -6488 -88468 -6300 -87980
rect -148 -88468 40 -87976
rect 6162 -88468 6350 -88048
rect -83242 -89592 7438 -88468
use sky130_fd_pr__cap_mim_m3_1_ZP6U3S  sky130_fd_pr__cap_mim_m3_1_ZP6U3S_0
timestamp 1635855079
transform 1 0 -41083 0 1 -41000
box -47383 -47250 47382 47250
<< labels >>
rlabel metal4 s -44568 7904 -44568 7904 4 VIN
port 1 nsew
rlabel metal4 s -41466 -89242 -41466 -89242 4 VOUT
port 2 nsew
<< end >>
