magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< error_p >>
rect -31 8072 31 8078
rect -31 8038 -17 8072
rect -31 8032 31 8038
rect -31 -8038 31 -8032
rect -31 -8072 -17 -8038
rect -31 -8078 31 -8072
<< pwell >>
rect -221 -8200 221 8200
<< nmoslvt >>
rect -35 -8000 35 8000
<< ndiff >>
rect -93 7973 -35 8000
rect -93 7939 -81 7973
rect -47 7939 -35 7973
rect -93 7905 -35 7939
rect -93 7871 -81 7905
rect -47 7871 -35 7905
rect -93 7837 -35 7871
rect -93 7803 -81 7837
rect -47 7803 -35 7837
rect -93 7769 -35 7803
rect -93 7735 -81 7769
rect -47 7735 -35 7769
rect -93 7701 -35 7735
rect -93 7667 -81 7701
rect -47 7667 -35 7701
rect -93 7633 -35 7667
rect -93 7599 -81 7633
rect -47 7599 -35 7633
rect -93 7565 -35 7599
rect -93 7531 -81 7565
rect -47 7531 -35 7565
rect -93 7497 -35 7531
rect -93 7463 -81 7497
rect -47 7463 -35 7497
rect -93 7429 -35 7463
rect -93 7395 -81 7429
rect -47 7395 -35 7429
rect -93 7361 -35 7395
rect -93 7327 -81 7361
rect -47 7327 -35 7361
rect -93 7293 -35 7327
rect -93 7259 -81 7293
rect -47 7259 -35 7293
rect -93 7225 -35 7259
rect -93 7191 -81 7225
rect -47 7191 -35 7225
rect -93 7157 -35 7191
rect -93 7123 -81 7157
rect -47 7123 -35 7157
rect -93 7089 -35 7123
rect -93 7055 -81 7089
rect -47 7055 -35 7089
rect -93 7021 -35 7055
rect -93 6987 -81 7021
rect -47 6987 -35 7021
rect -93 6953 -35 6987
rect -93 6919 -81 6953
rect -47 6919 -35 6953
rect -93 6885 -35 6919
rect -93 6851 -81 6885
rect -47 6851 -35 6885
rect -93 6817 -35 6851
rect -93 6783 -81 6817
rect -47 6783 -35 6817
rect -93 6749 -35 6783
rect -93 6715 -81 6749
rect -47 6715 -35 6749
rect -93 6681 -35 6715
rect -93 6647 -81 6681
rect -47 6647 -35 6681
rect -93 6613 -35 6647
rect -93 6579 -81 6613
rect -47 6579 -35 6613
rect -93 6545 -35 6579
rect -93 6511 -81 6545
rect -47 6511 -35 6545
rect -93 6477 -35 6511
rect -93 6443 -81 6477
rect -47 6443 -35 6477
rect -93 6409 -35 6443
rect -93 6375 -81 6409
rect -47 6375 -35 6409
rect -93 6341 -35 6375
rect -93 6307 -81 6341
rect -47 6307 -35 6341
rect -93 6273 -35 6307
rect -93 6239 -81 6273
rect -47 6239 -35 6273
rect -93 6205 -35 6239
rect -93 6171 -81 6205
rect -47 6171 -35 6205
rect -93 6137 -35 6171
rect -93 6103 -81 6137
rect -47 6103 -35 6137
rect -93 6069 -35 6103
rect -93 6035 -81 6069
rect -47 6035 -35 6069
rect -93 6001 -35 6035
rect -93 5967 -81 6001
rect -47 5967 -35 6001
rect -93 5933 -35 5967
rect -93 5899 -81 5933
rect -47 5899 -35 5933
rect -93 5865 -35 5899
rect -93 5831 -81 5865
rect -47 5831 -35 5865
rect -93 5797 -35 5831
rect -93 5763 -81 5797
rect -47 5763 -35 5797
rect -93 5729 -35 5763
rect -93 5695 -81 5729
rect -47 5695 -35 5729
rect -93 5661 -35 5695
rect -93 5627 -81 5661
rect -47 5627 -35 5661
rect -93 5593 -35 5627
rect -93 5559 -81 5593
rect -47 5559 -35 5593
rect -93 5525 -35 5559
rect -93 5491 -81 5525
rect -47 5491 -35 5525
rect -93 5457 -35 5491
rect -93 5423 -81 5457
rect -47 5423 -35 5457
rect -93 5389 -35 5423
rect -93 5355 -81 5389
rect -47 5355 -35 5389
rect -93 5321 -35 5355
rect -93 5287 -81 5321
rect -47 5287 -35 5321
rect -93 5253 -35 5287
rect -93 5219 -81 5253
rect -47 5219 -35 5253
rect -93 5185 -35 5219
rect -93 5151 -81 5185
rect -47 5151 -35 5185
rect -93 5117 -35 5151
rect -93 5083 -81 5117
rect -47 5083 -35 5117
rect -93 5049 -35 5083
rect -93 5015 -81 5049
rect -47 5015 -35 5049
rect -93 4981 -35 5015
rect -93 4947 -81 4981
rect -47 4947 -35 4981
rect -93 4913 -35 4947
rect -93 4879 -81 4913
rect -47 4879 -35 4913
rect -93 4845 -35 4879
rect -93 4811 -81 4845
rect -47 4811 -35 4845
rect -93 4777 -35 4811
rect -93 4743 -81 4777
rect -47 4743 -35 4777
rect -93 4709 -35 4743
rect -93 4675 -81 4709
rect -47 4675 -35 4709
rect -93 4641 -35 4675
rect -93 4607 -81 4641
rect -47 4607 -35 4641
rect -93 4573 -35 4607
rect -93 4539 -81 4573
rect -47 4539 -35 4573
rect -93 4505 -35 4539
rect -93 4471 -81 4505
rect -47 4471 -35 4505
rect -93 4437 -35 4471
rect -93 4403 -81 4437
rect -47 4403 -35 4437
rect -93 4369 -35 4403
rect -93 4335 -81 4369
rect -47 4335 -35 4369
rect -93 4301 -35 4335
rect -93 4267 -81 4301
rect -47 4267 -35 4301
rect -93 4233 -35 4267
rect -93 4199 -81 4233
rect -47 4199 -35 4233
rect -93 4165 -35 4199
rect -93 4131 -81 4165
rect -47 4131 -35 4165
rect -93 4097 -35 4131
rect -93 4063 -81 4097
rect -47 4063 -35 4097
rect -93 4029 -35 4063
rect -93 3995 -81 4029
rect -47 3995 -35 4029
rect -93 3961 -35 3995
rect -93 3927 -81 3961
rect -47 3927 -35 3961
rect -93 3893 -35 3927
rect -93 3859 -81 3893
rect -47 3859 -35 3893
rect -93 3825 -35 3859
rect -93 3791 -81 3825
rect -47 3791 -35 3825
rect -93 3757 -35 3791
rect -93 3723 -81 3757
rect -47 3723 -35 3757
rect -93 3689 -35 3723
rect -93 3655 -81 3689
rect -47 3655 -35 3689
rect -93 3621 -35 3655
rect -93 3587 -81 3621
rect -47 3587 -35 3621
rect -93 3553 -35 3587
rect -93 3519 -81 3553
rect -47 3519 -35 3553
rect -93 3485 -35 3519
rect -93 3451 -81 3485
rect -47 3451 -35 3485
rect -93 3417 -35 3451
rect -93 3383 -81 3417
rect -47 3383 -35 3417
rect -93 3349 -35 3383
rect -93 3315 -81 3349
rect -47 3315 -35 3349
rect -93 3281 -35 3315
rect -93 3247 -81 3281
rect -47 3247 -35 3281
rect -93 3213 -35 3247
rect -93 3179 -81 3213
rect -47 3179 -35 3213
rect -93 3145 -35 3179
rect -93 3111 -81 3145
rect -47 3111 -35 3145
rect -93 3077 -35 3111
rect -93 3043 -81 3077
rect -47 3043 -35 3077
rect -93 3009 -35 3043
rect -93 2975 -81 3009
rect -47 2975 -35 3009
rect -93 2941 -35 2975
rect -93 2907 -81 2941
rect -47 2907 -35 2941
rect -93 2873 -35 2907
rect -93 2839 -81 2873
rect -47 2839 -35 2873
rect -93 2805 -35 2839
rect -93 2771 -81 2805
rect -47 2771 -35 2805
rect -93 2737 -35 2771
rect -93 2703 -81 2737
rect -47 2703 -35 2737
rect -93 2669 -35 2703
rect -93 2635 -81 2669
rect -47 2635 -35 2669
rect -93 2601 -35 2635
rect -93 2567 -81 2601
rect -47 2567 -35 2601
rect -93 2533 -35 2567
rect -93 2499 -81 2533
rect -47 2499 -35 2533
rect -93 2465 -35 2499
rect -93 2431 -81 2465
rect -47 2431 -35 2465
rect -93 2397 -35 2431
rect -93 2363 -81 2397
rect -47 2363 -35 2397
rect -93 2329 -35 2363
rect -93 2295 -81 2329
rect -47 2295 -35 2329
rect -93 2261 -35 2295
rect -93 2227 -81 2261
rect -47 2227 -35 2261
rect -93 2193 -35 2227
rect -93 2159 -81 2193
rect -47 2159 -35 2193
rect -93 2125 -35 2159
rect -93 2091 -81 2125
rect -47 2091 -35 2125
rect -93 2057 -35 2091
rect -93 2023 -81 2057
rect -47 2023 -35 2057
rect -93 1989 -35 2023
rect -93 1955 -81 1989
rect -47 1955 -35 1989
rect -93 1921 -35 1955
rect -93 1887 -81 1921
rect -47 1887 -35 1921
rect -93 1853 -35 1887
rect -93 1819 -81 1853
rect -47 1819 -35 1853
rect -93 1785 -35 1819
rect -93 1751 -81 1785
rect -47 1751 -35 1785
rect -93 1717 -35 1751
rect -93 1683 -81 1717
rect -47 1683 -35 1717
rect -93 1649 -35 1683
rect -93 1615 -81 1649
rect -47 1615 -35 1649
rect -93 1581 -35 1615
rect -93 1547 -81 1581
rect -47 1547 -35 1581
rect -93 1513 -35 1547
rect -93 1479 -81 1513
rect -47 1479 -35 1513
rect -93 1445 -35 1479
rect -93 1411 -81 1445
rect -47 1411 -35 1445
rect -93 1377 -35 1411
rect -93 1343 -81 1377
rect -47 1343 -35 1377
rect -93 1309 -35 1343
rect -93 1275 -81 1309
rect -47 1275 -35 1309
rect -93 1241 -35 1275
rect -93 1207 -81 1241
rect -47 1207 -35 1241
rect -93 1173 -35 1207
rect -93 1139 -81 1173
rect -47 1139 -35 1173
rect -93 1105 -35 1139
rect -93 1071 -81 1105
rect -47 1071 -35 1105
rect -93 1037 -35 1071
rect -93 1003 -81 1037
rect -47 1003 -35 1037
rect -93 969 -35 1003
rect -93 935 -81 969
rect -47 935 -35 969
rect -93 901 -35 935
rect -93 867 -81 901
rect -47 867 -35 901
rect -93 833 -35 867
rect -93 799 -81 833
rect -47 799 -35 833
rect -93 765 -35 799
rect -93 731 -81 765
rect -47 731 -35 765
rect -93 697 -35 731
rect -93 663 -81 697
rect -47 663 -35 697
rect -93 629 -35 663
rect -93 595 -81 629
rect -47 595 -35 629
rect -93 561 -35 595
rect -93 527 -81 561
rect -47 527 -35 561
rect -93 493 -35 527
rect -93 459 -81 493
rect -47 459 -35 493
rect -93 425 -35 459
rect -93 391 -81 425
rect -47 391 -35 425
rect -93 357 -35 391
rect -93 323 -81 357
rect -47 323 -35 357
rect -93 289 -35 323
rect -93 255 -81 289
rect -47 255 -35 289
rect -93 221 -35 255
rect -93 187 -81 221
rect -47 187 -35 221
rect -93 153 -35 187
rect -93 119 -81 153
rect -47 119 -35 153
rect -93 85 -35 119
rect -93 51 -81 85
rect -47 51 -35 85
rect -93 17 -35 51
rect -93 -17 -81 17
rect -47 -17 -35 17
rect -93 -51 -35 -17
rect -93 -85 -81 -51
rect -47 -85 -35 -51
rect -93 -119 -35 -85
rect -93 -153 -81 -119
rect -47 -153 -35 -119
rect -93 -187 -35 -153
rect -93 -221 -81 -187
rect -47 -221 -35 -187
rect -93 -255 -35 -221
rect -93 -289 -81 -255
rect -47 -289 -35 -255
rect -93 -323 -35 -289
rect -93 -357 -81 -323
rect -47 -357 -35 -323
rect -93 -391 -35 -357
rect -93 -425 -81 -391
rect -47 -425 -35 -391
rect -93 -459 -35 -425
rect -93 -493 -81 -459
rect -47 -493 -35 -459
rect -93 -527 -35 -493
rect -93 -561 -81 -527
rect -47 -561 -35 -527
rect -93 -595 -35 -561
rect -93 -629 -81 -595
rect -47 -629 -35 -595
rect -93 -663 -35 -629
rect -93 -697 -81 -663
rect -47 -697 -35 -663
rect -93 -731 -35 -697
rect -93 -765 -81 -731
rect -47 -765 -35 -731
rect -93 -799 -35 -765
rect -93 -833 -81 -799
rect -47 -833 -35 -799
rect -93 -867 -35 -833
rect -93 -901 -81 -867
rect -47 -901 -35 -867
rect -93 -935 -35 -901
rect -93 -969 -81 -935
rect -47 -969 -35 -935
rect -93 -1003 -35 -969
rect -93 -1037 -81 -1003
rect -47 -1037 -35 -1003
rect -93 -1071 -35 -1037
rect -93 -1105 -81 -1071
rect -47 -1105 -35 -1071
rect -93 -1139 -35 -1105
rect -93 -1173 -81 -1139
rect -47 -1173 -35 -1139
rect -93 -1207 -35 -1173
rect -93 -1241 -81 -1207
rect -47 -1241 -35 -1207
rect -93 -1275 -35 -1241
rect -93 -1309 -81 -1275
rect -47 -1309 -35 -1275
rect -93 -1343 -35 -1309
rect -93 -1377 -81 -1343
rect -47 -1377 -35 -1343
rect -93 -1411 -35 -1377
rect -93 -1445 -81 -1411
rect -47 -1445 -35 -1411
rect -93 -1479 -35 -1445
rect -93 -1513 -81 -1479
rect -47 -1513 -35 -1479
rect -93 -1547 -35 -1513
rect -93 -1581 -81 -1547
rect -47 -1581 -35 -1547
rect -93 -1615 -35 -1581
rect -93 -1649 -81 -1615
rect -47 -1649 -35 -1615
rect -93 -1683 -35 -1649
rect -93 -1717 -81 -1683
rect -47 -1717 -35 -1683
rect -93 -1751 -35 -1717
rect -93 -1785 -81 -1751
rect -47 -1785 -35 -1751
rect -93 -1819 -35 -1785
rect -93 -1853 -81 -1819
rect -47 -1853 -35 -1819
rect -93 -1887 -35 -1853
rect -93 -1921 -81 -1887
rect -47 -1921 -35 -1887
rect -93 -1955 -35 -1921
rect -93 -1989 -81 -1955
rect -47 -1989 -35 -1955
rect -93 -2023 -35 -1989
rect -93 -2057 -81 -2023
rect -47 -2057 -35 -2023
rect -93 -2091 -35 -2057
rect -93 -2125 -81 -2091
rect -47 -2125 -35 -2091
rect -93 -2159 -35 -2125
rect -93 -2193 -81 -2159
rect -47 -2193 -35 -2159
rect -93 -2227 -35 -2193
rect -93 -2261 -81 -2227
rect -47 -2261 -35 -2227
rect -93 -2295 -35 -2261
rect -93 -2329 -81 -2295
rect -47 -2329 -35 -2295
rect -93 -2363 -35 -2329
rect -93 -2397 -81 -2363
rect -47 -2397 -35 -2363
rect -93 -2431 -35 -2397
rect -93 -2465 -81 -2431
rect -47 -2465 -35 -2431
rect -93 -2499 -35 -2465
rect -93 -2533 -81 -2499
rect -47 -2533 -35 -2499
rect -93 -2567 -35 -2533
rect -93 -2601 -81 -2567
rect -47 -2601 -35 -2567
rect -93 -2635 -35 -2601
rect -93 -2669 -81 -2635
rect -47 -2669 -35 -2635
rect -93 -2703 -35 -2669
rect -93 -2737 -81 -2703
rect -47 -2737 -35 -2703
rect -93 -2771 -35 -2737
rect -93 -2805 -81 -2771
rect -47 -2805 -35 -2771
rect -93 -2839 -35 -2805
rect -93 -2873 -81 -2839
rect -47 -2873 -35 -2839
rect -93 -2907 -35 -2873
rect -93 -2941 -81 -2907
rect -47 -2941 -35 -2907
rect -93 -2975 -35 -2941
rect -93 -3009 -81 -2975
rect -47 -3009 -35 -2975
rect -93 -3043 -35 -3009
rect -93 -3077 -81 -3043
rect -47 -3077 -35 -3043
rect -93 -3111 -35 -3077
rect -93 -3145 -81 -3111
rect -47 -3145 -35 -3111
rect -93 -3179 -35 -3145
rect -93 -3213 -81 -3179
rect -47 -3213 -35 -3179
rect -93 -3247 -35 -3213
rect -93 -3281 -81 -3247
rect -47 -3281 -35 -3247
rect -93 -3315 -35 -3281
rect -93 -3349 -81 -3315
rect -47 -3349 -35 -3315
rect -93 -3383 -35 -3349
rect -93 -3417 -81 -3383
rect -47 -3417 -35 -3383
rect -93 -3451 -35 -3417
rect -93 -3485 -81 -3451
rect -47 -3485 -35 -3451
rect -93 -3519 -35 -3485
rect -93 -3553 -81 -3519
rect -47 -3553 -35 -3519
rect -93 -3587 -35 -3553
rect -93 -3621 -81 -3587
rect -47 -3621 -35 -3587
rect -93 -3655 -35 -3621
rect -93 -3689 -81 -3655
rect -47 -3689 -35 -3655
rect -93 -3723 -35 -3689
rect -93 -3757 -81 -3723
rect -47 -3757 -35 -3723
rect -93 -3791 -35 -3757
rect -93 -3825 -81 -3791
rect -47 -3825 -35 -3791
rect -93 -3859 -35 -3825
rect -93 -3893 -81 -3859
rect -47 -3893 -35 -3859
rect -93 -3927 -35 -3893
rect -93 -3961 -81 -3927
rect -47 -3961 -35 -3927
rect -93 -3995 -35 -3961
rect -93 -4029 -81 -3995
rect -47 -4029 -35 -3995
rect -93 -4063 -35 -4029
rect -93 -4097 -81 -4063
rect -47 -4097 -35 -4063
rect -93 -4131 -35 -4097
rect -93 -4165 -81 -4131
rect -47 -4165 -35 -4131
rect -93 -4199 -35 -4165
rect -93 -4233 -81 -4199
rect -47 -4233 -35 -4199
rect -93 -4267 -35 -4233
rect -93 -4301 -81 -4267
rect -47 -4301 -35 -4267
rect -93 -4335 -35 -4301
rect -93 -4369 -81 -4335
rect -47 -4369 -35 -4335
rect -93 -4403 -35 -4369
rect -93 -4437 -81 -4403
rect -47 -4437 -35 -4403
rect -93 -4471 -35 -4437
rect -93 -4505 -81 -4471
rect -47 -4505 -35 -4471
rect -93 -4539 -35 -4505
rect -93 -4573 -81 -4539
rect -47 -4573 -35 -4539
rect -93 -4607 -35 -4573
rect -93 -4641 -81 -4607
rect -47 -4641 -35 -4607
rect -93 -4675 -35 -4641
rect -93 -4709 -81 -4675
rect -47 -4709 -35 -4675
rect -93 -4743 -35 -4709
rect -93 -4777 -81 -4743
rect -47 -4777 -35 -4743
rect -93 -4811 -35 -4777
rect -93 -4845 -81 -4811
rect -47 -4845 -35 -4811
rect -93 -4879 -35 -4845
rect -93 -4913 -81 -4879
rect -47 -4913 -35 -4879
rect -93 -4947 -35 -4913
rect -93 -4981 -81 -4947
rect -47 -4981 -35 -4947
rect -93 -5015 -35 -4981
rect -93 -5049 -81 -5015
rect -47 -5049 -35 -5015
rect -93 -5083 -35 -5049
rect -93 -5117 -81 -5083
rect -47 -5117 -35 -5083
rect -93 -5151 -35 -5117
rect -93 -5185 -81 -5151
rect -47 -5185 -35 -5151
rect -93 -5219 -35 -5185
rect -93 -5253 -81 -5219
rect -47 -5253 -35 -5219
rect -93 -5287 -35 -5253
rect -93 -5321 -81 -5287
rect -47 -5321 -35 -5287
rect -93 -5355 -35 -5321
rect -93 -5389 -81 -5355
rect -47 -5389 -35 -5355
rect -93 -5423 -35 -5389
rect -93 -5457 -81 -5423
rect -47 -5457 -35 -5423
rect -93 -5491 -35 -5457
rect -93 -5525 -81 -5491
rect -47 -5525 -35 -5491
rect -93 -5559 -35 -5525
rect -93 -5593 -81 -5559
rect -47 -5593 -35 -5559
rect -93 -5627 -35 -5593
rect -93 -5661 -81 -5627
rect -47 -5661 -35 -5627
rect -93 -5695 -35 -5661
rect -93 -5729 -81 -5695
rect -47 -5729 -35 -5695
rect -93 -5763 -35 -5729
rect -93 -5797 -81 -5763
rect -47 -5797 -35 -5763
rect -93 -5831 -35 -5797
rect -93 -5865 -81 -5831
rect -47 -5865 -35 -5831
rect -93 -5899 -35 -5865
rect -93 -5933 -81 -5899
rect -47 -5933 -35 -5899
rect -93 -5967 -35 -5933
rect -93 -6001 -81 -5967
rect -47 -6001 -35 -5967
rect -93 -6035 -35 -6001
rect -93 -6069 -81 -6035
rect -47 -6069 -35 -6035
rect -93 -6103 -35 -6069
rect -93 -6137 -81 -6103
rect -47 -6137 -35 -6103
rect -93 -6171 -35 -6137
rect -93 -6205 -81 -6171
rect -47 -6205 -35 -6171
rect -93 -6239 -35 -6205
rect -93 -6273 -81 -6239
rect -47 -6273 -35 -6239
rect -93 -6307 -35 -6273
rect -93 -6341 -81 -6307
rect -47 -6341 -35 -6307
rect -93 -6375 -35 -6341
rect -93 -6409 -81 -6375
rect -47 -6409 -35 -6375
rect -93 -6443 -35 -6409
rect -93 -6477 -81 -6443
rect -47 -6477 -35 -6443
rect -93 -6511 -35 -6477
rect -93 -6545 -81 -6511
rect -47 -6545 -35 -6511
rect -93 -6579 -35 -6545
rect -93 -6613 -81 -6579
rect -47 -6613 -35 -6579
rect -93 -6647 -35 -6613
rect -93 -6681 -81 -6647
rect -47 -6681 -35 -6647
rect -93 -6715 -35 -6681
rect -93 -6749 -81 -6715
rect -47 -6749 -35 -6715
rect -93 -6783 -35 -6749
rect -93 -6817 -81 -6783
rect -47 -6817 -35 -6783
rect -93 -6851 -35 -6817
rect -93 -6885 -81 -6851
rect -47 -6885 -35 -6851
rect -93 -6919 -35 -6885
rect -93 -6953 -81 -6919
rect -47 -6953 -35 -6919
rect -93 -6987 -35 -6953
rect -93 -7021 -81 -6987
rect -47 -7021 -35 -6987
rect -93 -7055 -35 -7021
rect -93 -7089 -81 -7055
rect -47 -7089 -35 -7055
rect -93 -7123 -35 -7089
rect -93 -7157 -81 -7123
rect -47 -7157 -35 -7123
rect -93 -7191 -35 -7157
rect -93 -7225 -81 -7191
rect -47 -7225 -35 -7191
rect -93 -7259 -35 -7225
rect -93 -7293 -81 -7259
rect -47 -7293 -35 -7259
rect -93 -7327 -35 -7293
rect -93 -7361 -81 -7327
rect -47 -7361 -35 -7327
rect -93 -7395 -35 -7361
rect -93 -7429 -81 -7395
rect -47 -7429 -35 -7395
rect -93 -7463 -35 -7429
rect -93 -7497 -81 -7463
rect -47 -7497 -35 -7463
rect -93 -7531 -35 -7497
rect -93 -7565 -81 -7531
rect -47 -7565 -35 -7531
rect -93 -7599 -35 -7565
rect -93 -7633 -81 -7599
rect -47 -7633 -35 -7599
rect -93 -7667 -35 -7633
rect -93 -7701 -81 -7667
rect -47 -7701 -35 -7667
rect -93 -7735 -35 -7701
rect -93 -7769 -81 -7735
rect -47 -7769 -35 -7735
rect -93 -7803 -35 -7769
rect -93 -7837 -81 -7803
rect -47 -7837 -35 -7803
rect -93 -7871 -35 -7837
rect -93 -7905 -81 -7871
rect -47 -7905 -35 -7871
rect -93 -7939 -35 -7905
rect -93 -7973 -81 -7939
rect -47 -7973 -35 -7939
rect -93 -8000 -35 -7973
rect 35 7973 93 8000
rect 35 7939 47 7973
rect 81 7939 93 7973
rect 35 7905 93 7939
rect 35 7871 47 7905
rect 81 7871 93 7905
rect 35 7837 93 7871
rect 35 7803 47 7837
rect 81 7803 93 7837
rect 35 7769 93 7803
rect 35 7735 47 7769
rect 81 7735 93 7769
rect 35 7701 93 7735
rect 35 7667 47 7701
rect 81 7667 93 7701
rect 35 7633 93 7667
rect 35 7599 47 7633
rect 81 7599 93 7633
rect 35 7565 93 7599
rect 35 7531 47 7565
rect 81 7531 93 7565
rect 35 7497 93 7531
rect 35 7463 47 7497
rect 81 7463 93 7497
rect 35 7429 93 7463
rect 35 7395 47 7429
rect 81 7395 93 7429
rect 35 7361 93 7395
rect 35 7327 47 7361
rect 81 7327 93 7361
rect 35 7293 93 7327
rect 35 7259 47 7293
rect 81 7259 93 7293
rect 35 7225 93 7259
rect 35 7191 47 7225
rect 81 7191 93 7225
rect 35 7157 93 7191
rect 35 7123 47 7157
rect 81 7123 93 7157
rect 35 7089 93 7123
rect 35 7055 47 7089
rect 81 7055 93 7089
rect 35 7021 93 7055
rect 35 6987 47 7021
rect 81 6987 93 7021
rect 35 6953 93 6987
rect 35 6919 47 6953
rect 81 6919 93 6953
rect 35 6885 93 6919
rect 35 6851 47 6885
rect 81 6851 93 6885
rect 35 6817 93 6851
rect 35 6783 47 6817
rect 81 6783 93 6817
rect 35 6749 93 6783
rect 35 6715 47 6749
rect 81 6715 93 6749
rect 35 6681 93 6715
rect 35 6647 47 6681
rect 81 6647 93 6681
rect 35 6613 93 6647
rect 35 6579 47 6613
rect 81 6579 93 6613
rect 35 6545 93 6579
rect 35 6511 47 6545
rect 81 6511 93 6545
rect 35 6477 93 6511
rect 35 6443 47 6477
rect 81 6443 93 6477
rect 35 6409 93 6443
rect 35 6375 47 6409
rect 81 6375 93 6409
rect 35 6341 93 6375
rect 35 6307 47 6341
rect 81 6307 93 6341
rect 35 6273 93 6307
rect 35 6239 47 6273
rect 81 6239 93 6273
rect 35 6205 93 6239
rect 35 6171 47 6205
rect 81 6171 93 6205
rect 35 6137 93 6171
rect 35 6103 47 6137
rect 81 6103 93 6137
rect 35 6069 93 6103
rect 35 6035 47 6069
rect 81 6035 93 6069
rect 35 6001 93 6035
rect 35 5967 47 6001
rect 81 5967 93 6001
rect 35 5933 93 5967
rect 35 5899 47 5933
rect 81 5899 93 5933
rect 35 5865 93 5899
rect 35 5831 47 5865
rect 81 5831 93 5865
rect 35 5797 93 5831
rect 35 5763 47 5797
rect 81 5763 93 5797
rect 35 5729 93 5763
rect 35 5695 47 5729
rect 81 5695 93 5729
rect 35 5661 93 5695
rect 35 5627 47 5661
rect 81 5627 93 5661
rect 35 5593 93 5627
rect 35 5559 47 5593
rect 81 5559 93 5593
rect 35 5525 93 5559
rect 35 5491 47 5525
rect 81 5491 93 5525
rect 35 5457 93 5491
rect 35 5423 47 5457
rect 81 5423 93 5457
rect 35 5389 93 5423
rect 35 5355 47 5389
rect 81 5355 93 5389
rect 35 5321 93 5355
rect 35 5287 47 5321
rect 81 5287 93 5321
rect 35 5253 93 5287
rect 35 5219 47 5253
rect 81 5219 93 5253
rect 35 5185 93 5219
rect 35 5151 47 5185
rect 81 5151 93 5185
rect 35 5117 93 5151
rect 35 5083 47 5117
rect 81 5083 93 5117
rect 35 5049 93 5083
rect 35 5015 47 5049
rect 81 5015 93 5049
rect 35 4981 93 5015
rect 35 4947 47 4981
rect 81 4947 93 4981
rect 35 4913 93 4947
rect 35 4879 47 4913
rect 81 4879 93 4913
rect 35 4845 93 4879
rect 35 4811 47 4845
rect 81 4811 93 4845
rect 35 4777 93 4811
rect 35 4743 47 4777
rect 81 4743 93 4777
rect 35 4709 93 4743
rect 35 4675 47 4709
rect 81 4675 93 4709
rect 35 4641 93 4675
rect 35 4607 47 4641
rect 81 4607 93 4641
rect 35 4573 93 4607
rect 35 4539 47 4573
rect 81 4539 93 4573
rect 35 4505 93 4539
rect 35 4471 47 4505
rect 81 4471 93 4505
rect 35 4437 93 4471
rect 35 4403 47 4437
rect 81 4403 93 4437
rect 35 4369 93 4403
rect 35 4335 47 4369
rect 81 4335 93 4369
rect 35 4301 93 4335
rect 35 4267 47 4301
rect 81 4267 93 4301
rect 35 4233 93 4267
rect 35 4199 47 4233
rect 81 4199 93 4233
rect 35 4165 93 4199
rect 35 4131 47 4165
rect 81 4131 93 4165
rect 35 4097 93 4131
rect 35 4063 47 4097
rect 81 4063 93 4097
rect 35 4029 93 4063
rect 35 3995 47 4029
rect 81 3995 93 4029
rect 35 3961 93 3995
rect 35 3927 47 3961
rect 81 3927 93 3961
rect 35 3893 93 3927
rect 35 3859 47 3893
rect 81 3859 93 3893
rect 35 3825 93 3859
rect 35 3791 47 3825
rect 81 3791 93 3825
rect 35 3757 93 3791
rect 35 3723 47 3757
rect 81 3723 93 3757
rect 35 3689 93 3723
rect 35 3655 47 3689
rect 81 3655 93 3689
rect 35 3621 93 3655
rect 35 3587 47 3621
rect 81 3587 93 3621
rect 35 3553 93 3587
rect 35 3519 47 3553
rect 81 3519 93 3553
rect 35 3485 93 3519
rect 35 3451 47 3485
rect 81 3451 93 3485
rect 35 3417 93 3451
rect 35 3383 47 3417
rect 81 3383 93 3417
rect 35 3349 93 3383
rect 35 3315 47 3349
rect 81 3315 93 3349
rect 35 3281 93 3315
rect 35 3247 47 3281
rect 81 3247 93 3281
rect 35 3213 93 3247
rect 35 3179 47 3213
rect 81 3179 93 3213
rect 35 3145 93 3179
rect 35 3111 47 3145
rect 81 3111 93 3145
rect 35 3077 93 3111
rect 35 3043 47 3077
rect 81 3043 93 3077
rect 35 3009 93 3043
rect 35 2975 47 3009
rect 81 2975 93 3009
rect 35 2941 93 2975
rect 35 2907 47 2941
rect 81 2907 93 2941
rect 35 2873 93 2907
rect 35 2839 47 2873
rect 81 2839 93 2873
rect 35 2805 93 2839
rect 35 2771 47 2805
rect 81 2771 93 2805
rect 35 2737 93 2771
rect 35 2703 47 2737
rect 81 2703 93 2737
rect 35 2669 93 2703
rect 35 2635 47 2669
rect 81 2635 93 2669
rect 35 2601 93 2635
rect 35 2567 47 2601
rect 81 2567 93 2601
rect 35 2533 93 2567
rect 35 2499 47 2533
rect 81 2499 93 2533
rect 35 2465 93 2499
rect 35 2431 47 2465
rect 81 2431 93 2465
rect 35 2397 93 2431
rect 35 2363 47 2397
rect 81 2363 93 2397
rect 35 2329 93 2363
rect 35 2295 47 2329
rect 81 2295 93 2329
rect 35 2261 93 2295
rect 35 2227 47 2261
rect 81 2227 93 2261
rect 35 2193 93 2227
rect 35 2159 47 2193
rect 81 2159 93 2193
rect 35 2125 93 2159
rect 35 2091 47 2125
rect 81 2091 93 2125
rect 35 2057 93 2091
rect 35 2023 47 2057
rect 81 2023 93 2057
rect 35 1989 93 2023
rect 35 1955 47 1989
rect 81 1955 93 1989
rect 35 1921 93 1955
rect 35 1887 47 1921
rect 81 1887 93 1921
rect 35 1853 93 1887
rect 35 1819 47 1853
rect 81 1819 93 1853
rect 35 1785 93 1819
rect 35 1751 47 1785
rect 81 1751 93 1785
rect 35 1717 93 1751
rect 35 1683 47 1717
rect 81 1683 93 1717
rect 35 1649 93 1683
rect 35 1615 47 1649
rect 81 1615 93 1649
rect 35 1581 93 1615
rect 35 1547 47 1581
rect 81 1547 93 1581
rect 35 1513 93 1547
rect 35 1479 47 1513
rect 81 1479 93 1513
rect 35 1445 93 1479
rect 35 1411 47 1445
rect 81 1411 93 1445
rect 35 1377 93 1411
rect 35 1343 47 1377
rect 81 1343 93 1377
rect 35 1309 93 1343
rect 35 1275 47 1309
rect 81 1275 93 1309
rect 35 1241 93 1275
rect 35 1207 47 1241
rect 81 1207 93 1241
rect 35 1173 93 1207
rect 35 1139 47 1173
rect 81 1139 93 1173
rect 35 1105 93 1139
rect 35 1071 47 1105
rect 81 1071 93 1105
rect 35 1037 93 1071
rect 35 1003 47 1037
rect 81 1003 93 1037
rect 35 969 93 1003
rect 35 935 47 969
rect 81 935 93 969
rect 35 901 93 935
rect 35 867 47 901
rect 81 867 93 901
rect 35 833 93 867
rect 35 799 47 833
rect 81 799 93 833
rect 35 765 93 799
rect 35 731 47 765
rect 81 731 93 765
rect 35 697 93 731
rect 35 663 47 697
rect 81 663 93 697
rect 35 629 93 663
rect 35 595 47 629
rect 81 595 93 629
rect 35 561 93 595
rect 35 527 47 561
rect 81 527 93 561
rect 35 493 93 527
rect 35 459 47 493
rect 81 459 93 493
rect 35 425 93 459
rect 35 391 47 425
rect 81 391 93 425
rect 35 357 93 391
rect 35 323 47 357
rect 81 323 93 357
rect 35 289 93 323
rect 35 255 47 289
rect 81 255 93 289
rect 35 221 93 255
rect 35 187 47 221
rect 81 187 93 221
rect 35 153 93 187
rect 35 119 47 153
rect 81 119 93 153
rect 35 85 93 119
rect 35 51 47 85
rect 81 51 93 85
rect 35 17 93 51
rect 35 -17 47 17
rect 81 -17 93 17
rect 35 -51 93 -17
rect 35 -85 47 -51
rect 81 -85 93 -51
rect 35 -119 93 -85
rect 35 -153 47 -119
rect 81 -153 93 -119
rect 35 -187 93 -153
rect 35 -221 47 -187
rect 81 -221 93 -187
rect 35 -255 93 -221
rect 35 -289 47 -255
rect 81 -289 93 -255
rect 35 -323 93 -289
rect 35 -357 47 -323
rect 81 -357 93 -323
rect 35 -391 93 -357
rect 35 -425 47 -391
rect 81 -425 93 -391
rect 35 -459 93 -425
rect 35 -493 47 -459
rect 81 -493 93 -459
rect 35 -527 93 -493
rect 35 -561 47 -527
rect 81 -561 93 -527
rect 35 -595 93 -561
rect 35 -629 47 -595
rect 81 -629 93 -595
rect 35 -663 93 -629
rect 35 -697 47 -663
rect 81 -697 93 -663
rect 35 -731 93 -697
rect 35 -765 47 -731
rect 81 -765 93 -731
rect 35 -799 93 -765
rect 35 -833 47 -799
rect 81 -833 93 -799
rect 35 -867 93 -833
rect 35 -901 47 -867
rect 81 -901 93 -867
rect 35 -935 93 -901
rect 35 -969 47 -935
rect 81 -969 93 -935
rect 35 -1003 93 -969
rect 35 -1037 47 -1003
rect 81 -1037 93 -1003
rect 35 -1071 93 -1037
rect 35 -1105 47 -1071
rect 81 -1105 93 -1071
rect 35 -1139 93 -1105
rect 35 -1173 47 -1139
rect 81 -1173 93 -1139
rect 35 -1207 93 -1173
rect 35 -1241 47 -1207
rect 81 -1241 93 -1207
rect 35 -1275 93 -1241
rect 35 -1309 47 -1275
rect 81 -1309 93 -1275
rect 35 -1343 93 -1309
rect 35 -1377 47 -1343
rect 81 -1377 93 -1343
rect 35 -1411 93 -1377
rect 35 -1445 47 -1411
rect 81 -1445 93 -1411
rect 35 -1479 93 -1445
rect 35 -1513 47 -1479
rect 81 -1513 93 -1479
rect 35 -1547 93 -1513
rect 35 -1581 47 -1547
rect 81 -1581 93 -1547
rect 35 -1615 93 -1581
rect 35 -1649 47 -1615
rect 81 -1649 93 -1615
rect 35 -1683 93 -1649
rect 35 -1717 47 -1683
rect 81 -1717 93 -1683
rect 35 -1751 93 -1717
rect 35 -1785 47 -1751
rect 81 -1785 93 -1751
rect 35 -1819 93 -1785
rect 35 -1853 47 -1819
rect 81 -1853 93 -1819
rect 35 -1887 93 -1853
rect 35 -1921 47 -1887
rect 81 -1921 93 -1887
rect 35 -1955 93 -1921
rect 35 -1989 47 -1955
rect 81 -1989 93 -1955
rect 35 -2023 93 -1989
rect 35 -2057 47 -2023
rect 81 -2057 93 -2023
rect 35 -2091 93 -2057
rect 35 -2125 47 -2091
rect 81 -2125 93 -2091
rect 35 -2159 93 -2125
rect 35 -2193 47 -2159
rect 81 -2193 93 -2159
rect 35 -2227 93 -2193
rect 35 -2261 47 -2227
rect 81 -2261 93 -2227
rect 35 -2295 93 -2261
rect 35 -2329 47 -2295
rect 81 -2329 93 -2295
rect 35 -2363 93 -2329
rect 35 -2397 47 -2363
rect 81 -2397 93 -2363
rect 35 -2431 93 -2397
rect 35 -2465 47 -2431
rect 81 -2465 93 -2431
rect 35 -2499 93 -2465
rect 35 -2533 47 -2499
rect 81 -2533 93 -2499
rect 35 -2567 93 -2533
rect 35 -2601 47 -2567
rect 81 -2601 93 -2567
rect 35 -2635 93 -2601
rect 35 -2669 47 -2635
rect 81 -2669 93 -2635
rect 35 -2703 93 -2669
rect 35 -2737 47 -2703
rect 81 -2737 93 -2703
rect 35 -2771 93 -2737
rect 35 -2805 47 -2771
rect 81 -2805 93 -2771
rect 35 -2839 93 -2805
rect 35 -2873 47 -2839
rect 81 -2873 93 -2839
rect 35 -2907 93 -2873
rect 35 -2941 47 -2907
rect 81 -2941 93 -2907
rect 35 -2975 93 -2941
rect 35 -3009 47 -2975
rect 81 -3009 93 -2975
rect 35 -3043 93 -3009
rect 35 -3077 47 -3043
rect 81 -3077 93 -3043
rect 35 -3111 93 -3077
rect 35 -3145 47 -3111
rect 81 -3145 93 -3111
rect 35 -3179 93 -3145
rect 35 -3213 47 -3179
rect 81 -3213 93 -3179
rect 35 -3247 93 -3213
rect 35 -3281 47 -3247
rect 81 -3281 93 -3247
rect 35 -3315 93 -3281
rect 35 -3349 47 -3315
rect 81 -3349 93 -3315
rect 35 -3383 93 -3349
rect 35 -3417 47 -3383
rect 81 -3417 93 -3383
rect 35 -3451 93 -3417
rect 35 -3485 47 -3451
rect 81 -3485 93 -3451
rect 35 -3519 93 -3485
rect 35 -3553 47 -3519
rect 81 -3553 93 -3519
rect 35 -3587 93 -3553
rect 35 -3621 47 -3587
rect 81 -3621 93 -3587
rect 35 -3655 93 -3621
rect 35 -3689 47 -3655
rect 81 -3689 93 -3655
rect 35 -3723 93 -3689
rect 35 -3757 47 -3723
rect 81 -3757 93 -3723
rect 35 -3791 93 -3757
rect 35 -3825 47 -3791
rect 81 -3825 93 -3791
rect 35 -3859 93 -3825
rect 35 -3893 47 -3859
rect 81 -3893 93 -3859
rect 35 -3927 93 -3893
rect 35 -3961 47 -3927
rect 81 -3961 93 -3927
rect 35 -3995 93 -3961
rect 35 -4029 47 -3995
rect 81 -4029 93 -3995
rect 35 -4063 93 -4029
rect 35 -4097 47 -4063
rect 81 -4097 93 -4063
rect 35 -4131 93 -4097
rect 35 -4165 47 -4131
rect 81 -4165 93 -4131
rect 35 -4199 93 -4165
rect 35 -4233 47 -4199
rect 81 -4233 93 -4199
rect 35 -4267 93 -4233
rect 35 -4301 47 -4267
rect 81 -4301 93 -4267
rect 35 -4335 93 -4301
rect 35 -4369 47 -4335
rect 81 -4369 93 -4335
rect 35 -4403 93 -4369
rect 35 -4437 47 -4403
rect 81 -4437 93 -4403
rect 35 -4471 93 -4437
rect 35 -4505 47 -4471
rect 81 -4505 93 -4471
rect 35 -4539 93 -4505
rect 35 -4573 47 -4539
rect 81 -4573 93 -4539
rect 35 -4607 93 -4573
rect 35 -4641 47 -4607
rect 81 -4641 93 -4607
rect 35 -4675 93 -4641
rect 35 -4709 47 -4675
rect 81 -4709 93 -4675
rect 35 -4743 93 -4709
rect 35 -4777 47 -4743
rect 81 -4777 93 -4743
rect 35 -4811 93 -4777
rect 35 -4845 47 -4811
rect 81 -4845 93 -4811
rect 35 -4879 93 -4845
rect 35 -4913 47 -4879
rect 81 -4913 93 -4879
rect 35 -4947 93 -4913
rect 35 -4981 47 -4947
rect 81 -4981 93 -4947
rect 35 -5015 93 -4981
rect 35 -5049 47 -5015
rect 81 -5049 93 -5015
rect 35 -5083 93 -5049
rect 35 -5117 47 -5083
rect 81 -5117 93 -5083
rect 35 -5151 93 -5117
rect 35 -5185 47 -5151
rect 81 -5185 93 -5151
rect 35 -5219 93 -5185
rect 35 -5253 47 -5219
rect 81 -5253 93 -5219
rect 35 -5287 93 -5253
rect 35 -5321 47 -5287
rect 81 -5321 93 -5287
rect 35 -5355 93 -5321
rect 35 -5389 47 -5355
rect 81 -5389 93 -5355
rect 35 -5423 93 -5389
rect 35 -5457 47 -5423
rect 81 -5457 93 -5423
rect 35 -5491 93 -5457
rect 35 -5525 47 -5491
rect 81 -5525 93 -5491
rect 35 -5559 93 -5525
rect 35 -5593 47 -5559
rect 81 -5593 93 -5559
rect 35 -5627 93 -5593
rect 35 -5661 47 -5627
rect 81 -5661 93 -5627
rect 35 -5695 93 -5661
rect 35 -5729 47 -5695
rect 81 -5729 93 -5695
rect 35 -5763 93 -5729
rect 35 -5797 47 -5763
rect 81 -5797 93 -5763
rect 35 -5831 93 -5797
rect 35 -5865 47 -5831
rect 81 -5865 93 -5831
rect 35 -5899 93 -5865
rect 35 -5933 47 -5899
rect 81 -5933 93 -5899
rect 35 -5967 93 -5933
rect 35 -6001 47 -5967
rect 81 -6001 93 -5967
rect 35 -6035 93 -6001
rect 35 -6069 47 -6035
rect 81 -6069 93 -6035
rect 35 -6103 93 -6069
rect 35 -6137 47 -6103
rect 81 -6137 93 -6103
rect 35 -6171 93 -6137
rect 35 -6205 47 -6171
rect 81 -6205 93 -6171
rect 35 -6239 93 -6205
rect 35 -6273 47 -6239
rect 81 -6273 93 -6239
rect 35 -6307 93 -6273
rect 35 -6341 47 -6307
rect 81 -6341 93 -6307
rect 35 -6375 93 -6341
rect 35 -6409 47 -6375
rect 81 -6409 93 -6375
rect 35 -6443 93 -6409
rect 35 -6477 47 -6443
rect 81 -6477 93 -6443
rect 35 -6511 93 -6477
rect 35 -6545 47 -6511
rect 81 -6545 93 -6511
rect 35 -6579 93 -6545
rect 35 -6613 47 -6579
rect 81 -6613 93 -6579
rect 35 -6647 93 -6613
rect 35 -6681 47 -6647
rect 81 -6681 93 -6647
rect 35 -6715 93 -6681
rect 35 -6749 47 -6715
rect 81 -6749 93 -6715
rect 35 -6783 93 -6749
rect 35 -6817 47 -6783
rect 81 -6817 93 -6783
rect 35 -6851 93 -6817
rect 35 -6885 47 -6851
rect 81 -6885 93 -6851
rect 35 -6919 93 -6885
rect 35 -6953 47 -6919
rect 81 -6953 93 -6919
rect 35 -6987 93 -6953
rect 35 -7021 47 -6987
rect 81 -7021 93 -6987
rect 35 -7055 93 -7021
rect 35 -7089 47 -7055
rect 81 -7089 93 -7055
rect 35 -7123 93 -7089
rect 35 -7157 47 -7123
rect 81 -7157 93 -7123
rect 35 -7191 93 -7157
rect 35 -7225 47 -7191
rect 81 -7225 93 -7191
rect 35 -7259 93 -7225
rect 35 -7293 47 -7259
rect 81 -7293 93 -7259
rect 35 -7327 93 -7293
rect 35 -7361 47 -7327
rect 81 -7361 93 -7327
rect 35 -7395 93 -7361
rect 35 -7429 47 -7395
rect 81 -7429 93 -7395
rect 35 -7463 93 -7429
rect 35 -7497 47 -7463
rect 81 -7497 93 -7463
rect 35 -7531 93 -7497
rect 35 -7565 47 -7531
rect 81 -7565 93 -7531
rect 35 -7599 93 -7565
rect 35 -7633 47 -7599
rect 81 -7633 93 -7599
rect 35 -7667 93 -7633
rect 35 -7701 47 -7667
rect 81 -7701 93 -7667
rect 35 -7735 93 -7701
rect 35 -7769 47 -7735
rect 81 -7769 93 -7735
rect 35 -7803 93 -7769
rect 35 -7837 47 -7803
rect 81 -7837 93 -7803
rect 35 -7871 93 -7837
rect 35 -7905 47 -7871
rect 81 -7905 93 -7871
rect 35 -7939 93 -7905
rect 35 -7973 47 -7939
rect 81 -7973 93 -7939
rect 35 -8000 93 -7973
<< ndiffc >>
rect -81 7939 -47 7973
rect -81 7871 -47 7905
rect -81 7803 -47 7837
rect -81 7735 -47 7769
rect -81 7667 -47 7701
rect -81 7599 -47 7633
rect -81 7531 -47 7565
rect -81 7463 -47 7497
rect -81 7395 -47 7429
rect -81 7327 -47 7361
rect -81 7259 -47 7293
rect -81 7191 -47 7225
rect -81 7123 -47 7157
rect -81 7055 -47 7089
rect -81 6987 -47 7021
rect -81 6919 -47 6953
rect -81 6851 -47 6885
rect -81 6783 -47 6817
rect -81 6715 -47 6749
rect -81 6647 -47 6681
rect -81 6579 -47 6613
rect -81 6511 -47 6545
rect -81 6443 -47 6477
rect -81 6375 -47 6409
rect -81 6307 -47 6341
rect -81 6239 -47 6273
rect -81 6171 -47 6205
rect -81 6103 -47 6137
rect -81 6035 -47 6069
rect -81 5967 -47 6001
rect -81 5899 -47 5933
rect -81 5831 -47 5865
rect -81 5763 -47 5797
rect -81 5695 -47 5729
rect -81 5627 -47 5661
rect -81 5559 -47 5593
rect -81 5491 -47 5525
rect -81 5423 -47 5457
rect -81 5355 -47 5389
rect -81 5287 -47 5321
rect -81 5219 -47 5253
rect -81 5151 -47 5185
rect -81 5083 -47 5117
rect -81 5015 -47 5049
rect -81 4947 -47 4981
rect -81 4879 -47 4913
rect -81 4811 -47 4845
rect -81 4743 -47 4777
rect -81 4675 -47 4709
rect -81 4607 -47 4641
rect -81 4539 -47 4573
rect -81 4471 -47 4505
rect -81 4403 -47 4437
rect -81 4335 -47 4369
rect -81 4267 -47 4301
rect -81 4199 -47 4233
rect -81 4131 -47 4165
rect -81 4063 -47 4097
rect -81 3995 -47 4029
rect -81 3927 -47 3961
rect -81 3859 -47 3893
rect -81 3791 -47 3825
rect -81 3723 -47 3757
rect -81 3655 -47 3689
rect -81 3587 -47 3621
rect -81 3519 -47 3553
rect -81 3451 -47 3485
rect -81 3383 -47 3417
rect -81 3315 -47 3349
rect -81 3247 -47 3281
rect -81 3179 -47 3213
rect -81 3111 -47 3145
rect -81 3043 -47 3077
rect -81 2975 -47 3009
rect -81 2907 -47 2941
rect -81 2839 -47 2873
rect -81 2771 -47 2805
rect -81 2703 -47 2737
rect -81 2635 -47 2669
rect -81 2567 -47 2601
rect -81 2499 -47 2533
rect -81 2431 -47 2465
rect -81 2363 -47 2397
rect -81 2295 -47 2329
rect -81 2227 -47 2261
rect -81 2159 -47 2193
rect -81 2091 -47 2125
rect -81 2023 -47 2057
rect -81 1955 -47 1989
rect -81 1887 -47 1921
rect -81 1819 -47 1853
rect -81 1751 -47 1785
rect -81 1683 -47 1717
rect -81 1615 -47 1649
rect -81 1547 -47 1581
rect -81 1479 -47 1513
rect -81 1411 -47 1445
rect -81 1343 -47 1377
rect -81 1275 -47 1309
rect -81 1207 -47 1241
rect -81 1139 -47 1173
rect -81 1071 -47 1105
rect -81 1003 -47 1037
rect -81 935 -47 969
rect -81 867 -47 901
rect -81 799 -47 833
rect -81 731 -47 765
rect -81 663 -47 697
rect -81 595 -47 629
rect -81 527 -47 561
rect -81 459 -47 493
rect -81 391 -47 425
rect -81 323 -47 357
rect -81 255 -47 289
rect -81 187 -47 221
rect -81 119 -47 153
rect -81 51 -47 85
rect -81 -17 -47 17
rect -81 -85 -47 -51
rect -81 -153 -47 -119
rect -81 -221 -47 -187
rect -81 -289 -47 -255
rect -81 -357 -47 -323
rect -81 -425 -47 -391
rect -81 -493 -47 -459
rect -81 -561 -47 -527
rect -81 -629 -47 -595
rect -81 -697 -47 -663
rect -81 -765 -47 -731
rect -81 -833 -47 -799
rect -81 -901 -47 -867
rect -81 -969 -47 -935
rect -81 -1037 -47 -1003
rect -81 -1105 -47 -1071
rect -81 -1173 -47 -1139
rect -81 -1241 -47 -1207
rect -81 -1309 -47 -1275
rect -81 -1377 -47 -1343
rect -81 -1445 -47 -1411
rect -81 -1513 -47 -1479
rect -81 -1581 -47 -1547
rect -81 -1649 -47 -1615
rect -81 -1717 -47 -1683
rect -81 -1785 -47 -1751
rect -81 -1853 -47 -1819
rect -81 -1921 -47 -1887
rect -81 -1989 -47 -1955
rect -81 -2057 -47 -2023
rect -81 -2125 -47 -2091
rect -81 -2193 -47 -2159
rect -81 -2261 -47 -2227
rect -81 -2329 -47 -2295
rect -81 -2397 -47 -2363
rect -81 -2465 -47 -2431
rect -81 -2533 -47 -2499
rect -81 -2601 -47 -2567
rect -81 -2669 -47 -2635
rect -81 -2737 -47 -2703
rect -81 -2805 -47 -2771
rect -81 -2873 -47 -2839
rect -81 -2941 -47 -2907
rect -81 -3009 -47 -2975
rect -81 -3077 -47 -3043
rect -81 -3145 -47 -3111
rect -81 -3213 -47 -3179
rect -81 -3281 -47 -3247
rect -81 -3349 -47 -3315
rect -81 -3417 -47 -3383
rect -81 -3485 -47 -3451
rect -81 -3553 -47 -3519
rect -81 -3621 -47 -3587
rect -81 -3689 -47 -3655
rect -81 -3757 -47 -3723
rect -81 -3825 -47 -3791
rect -81 -3893 -47 -3859
rect -81 -3961 -47 -3927
rect -81 -4029 -47 -3995
rect -81 -4097 -47 -4063
rect -81 -4165 -47 -4131
rect -81 -4233 -47 -4199
rect -81 -4301 -47 -4267
rect -81 -4369 -47 -4335
rect -81 -4437 -47 -4403
rect -81 -4505 -47 -4471
rect -81 -4573 -47 -4539
rect -81 -4641 -47 -4607
rect -81 -4709 -47 -4675
rect -81 -4777 -47 -4743
rect -81 -4845 -47 -4811
rect -81 -4913 -47 -4879
rect -81 -4981 -47 -4947
rect -81 -5049 -47 -5015
rect -81 -5117 -47 -5083
rect -81 -5185 -47 -5151
rect -81 -5253 -47 -5219
rect -81 -5321 -47 -5287
rect -81 -5389 -47 -5355
rect -81 -5457 -47 -5423
rect -81 -5525 -47 -5491
rect -81 -5593 -47 -5559
rect -81 -5661 -47 -5627
rect -81 -5729 -47 -5695
rect -81 -5797 -47 -5763
rect -81 -5865 -47 -5831
rect -81 -5933 -47 -5899
rect -81 -6001 -47 -5967
rect -81 -6069 -47 -6035
rect -81 -6137 -47 -6103
rect -81 -6205 -47 -6171
rect -81 -6273 -47 -6239
rect -81 -6341 -47 -6307
rect -81 -6409 -47 -6375
rect -81 -6477 -47 -6443
rect -81 -6545 -47 -6511
rect -81 -6613 -47 -6579
rect -81 -6681 -47 -6647
rect -81 -6749 -47 -6715
rect -81 -6817 -47 -6783
rect -81 -6885 -47 -6851
rect -81 -6953 -47 -6919
rect -81 -7021 -47 -6987
rect -81 -7089 -47 -7055
rect -81 -7157 -47 -7123
rect -81 -7225 -47 -7191
rect -81 -7293 -47 -7259
rect -81 -7361 -47 -7327
rect -81 -7429 -47 -7395
rect -81 -7497 -47 -7463
rect -81 -7565 -47 -7531
rect -81 -7633 -47 -7599
rect -81 -7701 -47 -7667
rect -81 -7769 -47 -7735
rect -81 -7837 -47 -7803
rect -81 -7905 -47 -7871
rect -81 -7973 -47 -7939
rect 47 7939 81 7973
rect 47 7871 81 7905
rect 47 7803 81 7837
rect 47 7735 81 7769
rect 47 7667 81 7701
rect 47 7599 81 7633
rect 47 7531 81 7565
rect 47 7463 81 7497
rect 47 7395 81 7429
rect 47 7327 81 7361
rect 47 7259 81 7293
rect 47 7191 81 7225
rect 47 7123 81 7157
rect 47 7055 81 7089
rect 47 6987 81 7021
rect 47 6919 81 6953
rect 47 6851 81 6885
rect 47 6783 81 6817
rect 47 6715 81 6749
rect 47 6647 81 6681
rect 47 6579 81 6613
rect 47 6511 81 6545
rect 47 6443 81 6477
rect 47 6375 81 6409
rect 47 6307 81 6341
rect 47 6239 81 6273
rect 47 6171 81 6205
rect 47 6103 81 6137
rect 47 6035 81 6069
rect 47 5967 81 6001
rect 47 5899 81 5933
rect 47 5831 81 5865
rect 47 5763 81 5797
rect 47 5695 81 5729
rect 47 5627 81 5661
rect 47 5559 81 5593
rect 47 5491 81 5525
rect 47 5423 81 5457
rect 47 5355 81 5389
rect 47 5287 81 5321
rect 47 5219 81 5253
rect 47 5151 81 5185
rect 47 5083 81 5117
rect 47 5015 81 5049
rect 47 4947 81 4981
rect 47 4879 81 4913
rect 47 4811 81 4845
rect 47 4743 81 4777
rect 47 4675 81 4709
rect 47 4607 81 4641
rect 47 4539 81 4573
rect 47 4471 81 4505
rect 47 4403 81 4437
rect 47 4335 81 4369
rect 47 4267 81 4301
rect 47 4199 81 4233
rect 47 4131 81 4165
rect 47 4063 81 4097
rect 47 3995 81 4029
rect 47 3927 81 3961
rect 47 3859 81 3893
rect 47 3791 81 3825
rect 47 3723 81 3757
rect 47 3655 81 3689
rect 47 3587 81 3621
rect 47 3519 81 3553
rect 47 3451 81 3485
rect 47 3383 81 3417
rect 47 3315 81 3349
rect 47 3247 81 3281
rect 47 3179 81 3213
rect 47 3111 81 3145
rect 47 3043 81 3077
rect 47 2975 81 3009
rect 47 2907 81 2941
rect 47 2839 81 2873
rect 47 2771 81 2805
rect 47 2703 81 2737
rect 47 2635 81 2669
rect 47 2567 81 2601
rect 47 2499 81 2533
rect 47 2431 81 2465
rect 47 2363 81 2397
rect 47 2295 81 2329
rect 47 2227 81 2261
rect 47 2159 81 2193
rect 47 2091 81 2125
rect 47 2023 81 2057
rect 47 1955 81 1989
rect 47 1887 81 1921
rect 47 1819 81 1853
rect 47 1751 81 1785
rect 47 1683 81 1717
rect 47 1615 81 1649
rect 47 1547 81 1581
rect 47 1479 81 1513
rect 47 1411 81 1445
rect 47 1343 81 1377
rect 47 1275 81 1309
rect 47 1207 81 1241
rect 47 1139 81 1173
rect 47 1071 81 1105
rect 47 1003 81 1037
rect 47 935 81 969
rect 47 867 81 901
rect 47 799 81 833
rect 47 731 81 765
rect 47 663 81 697
rect 47 595 81 629
rect 47 527 81 561
rect 47 459 81 493
rect 47 391 81 425
rect 47 323 81 357
rect 47 255 81 289
rect 47 187 81 221
rect 47 119 81 153
rect 47 51 81 85
rect 47 -17 81 17
rect 47 -85 81 -51
rect 47 -153 81 -119
rect 47 -221 81 -187
rect 47 -289 81 -255
rect 47 -357 81 -323
rect 47 -425 81 -391
rect 47 -493 81 -459
rect 47 -561 81 -527
rect 47 -629 81 -595
rect 47 -697 81 -663
rect 47 -765 81 -731
rect 47 -833 81 -799
rect 47 -901 81 -867
rect 47 -969 81 -935
rect 47 -1037 81 -1003
rect 47 -1105 81 -1071
rect 47 -1173 81 -1139
rect 47 -1241 81 -1207
rect 47 -1309 81 -1275
rect 47 -1377 81 -1343
rect 47 -1445 81 -1411
rect 47 -1513 81 -1479
rect 47 -1581 81 -1547
rect 47 -1649 81 -1615
rect 47 -1717 81 -1683
rect 47 -1785 81 -1751
rect 47 -1853 81 -1819
rect 47 -1921 81 -1887
rect 47 -1989 81 -1955
rect 47 -2057 81 -2023
rect 47 -2125 81 -2091
rect 47 -2193 81 -2159
rect 47 -2261 81 -2227
rect 47 -2329 81 -2295
rect 47 -2397 81 -2363
rect 47 -2465 81 -2431
rect 47 -2533 81 -2499
rect 47 -2601 81 -2567
rect 47 -2669 81 -2635
rect 47 -2737 81 -2703
rect 47 -2805 81 -2771
rect 47 -2873 81 -2839
rect 47 -2941 81 -2907
rect 47 -3009 81 -2975
rect 47 -3077 81 -3043
rect 47 -3145 81 -3111
rect 47 -3213 81 -3179
rect 47 -3281 81 -3247
rect 47 -3349 81 -3315
rect 47 -3417 81 -3383
rect 47 -3485 81 -3451
rect 47 -3553 81 -3519
rect 47 -3621 81 -3587
rect 47 -3689 81 -3655
rect 47 -3757 81 -3723
rect 47 -3825 81 -3791
rect 47 -3893 81 -3859
rect 47 -3961 81 -3927
rect 47 -4029 81 -3995
rect 47 -4097 81 -4063
rect 47 -4165 81 -4131
rect 47 -4233 81 -4199
rect 47 -4301 81 -4267
rect 47 -4369 81 -4335
rect 47 -4437 81 -4403
rect 47 -4505 81 -4471
rect 47 -4573 81 -4539
rect 47 -4641 81 -4607
rect 47 -4709 81 -4675
rect 47 -4777 81 -4743
rect 47 -4845 81 -4811
rect 47 -4913 81 -4879
rect 47 -4981 81 -4947
rect 47 -5049 81 -5015
rect 47 -5117 81 -5083
rect 47 -5185 81 -5151
rect 47 -5253 81 -5219
rect 47 -5321 81 -5287
rect 47 -5389 81 -5355
rect 47 -5457 81 -5423
rect 47 -5525 81 -5491
rect 47 -5593 81 -5559
rect 47 -5661 81 -5627
rect 47 -5729 81 -5695
rect 47 -5797 81 -5763
rect 47 -5865 81 -5831
rect 47 -5933 81 -5899
rect 47 -6001 81 -5967
rect 47 -6069 81 -6035
rect 47 -6137 81 -6103
rect 47 -6205 81 -6171
rect 47 -6273 81 -6239
rect 47 -6341 81 -6307
rect 47 -6409 81 -6375
rect 47 -6477 81 -6443
rect 47 -6545 81 -6511
rect 47 -6613 81 -6579
rect 47 -6681 81 -6647
rect 47 -6749 81 -6715
rect 47 -6817 81 -6783
rect 47 -6885 81 -6851
rect 47 -6953 81 -6919
rect 47 -7021 81 -6987
rect 47 -7089 81 -7055
rect 47 -7157 81 -7123
rect 47 -7225 81 -7191
rect 47 -7293 81 -7259
rect 47 -7361 81 -7327
rect 47 -7429 81 -7395
rect 47 -7497 81 -7463
rect 47 -7565 81 -7531
rect 47 -7633 81 -7599
rect 47 -7701 81 -7667
rect 47 -7769 81 -7735
rect 47 -7837 81 -7803
rect 47 -7905 81 -7871
rect 47 -7973 81 -7939
<< psubdiff >>
rect -195 8140 -85 8174
rect -51 8140 -17 8174
rect 17 8140 51 8174
rect 85 8140 195 8174
rect -195 8075 -161 8140
rect -195 8007 -161 8041
rect 161 8075 195 8140
rect 161 8007 195 8041
rect -195 7939 -161 7973
rect -195 7871 -161 7905
rect -195 7803 -161 7837
rect -195 7735 -161 7769
rect -195 7667 -161 7701
rect -195 7599 -161 7633
rect -195 7531 -161 7565
rect -195 7463 -161 7497
rect -195 7395 -161 7429
rect -195 7327 -161 7361
rect -195 7259 -161 7293
rect -195 7191 -161 7225
rect -195 7123 -161 7157
rect -195 7055 -161 7089
rect -195 6987 -161 7021
rect -195 6919 -161 6953
rect -195 6851 -161 6885
rect -195 6783 -161 6817
rect -195 6715 -161 6749
rect -195 6647 -161 6681
rect -195 6579 -161 6613
rect -195 6511 -161 6545
rect -195 6443 -161 6477
rect -195 6375 -161 6409
rect -195 6307 -161 6341
rect -195 6239 -161 6273
rect -195 6171 -161 6205
rect -195 6103 -161 6137
rect -195 6035 -161 6069
rect -195 5967 -161 6001
rect -195 5899 -161 5933
rect -195 5831 -161 5865
rect -195 5763 -161 5797
rect -195 5695 -161 5729
rect -195 5627 -161 5661
rect -195 5559 -161 5593
rect -195 5491 -161 5525
rect -195 5423 -161 5457
rect -195 5355 -161 5389
rect -195 5287 -161 5321
rect -195 5219 -161 5253
rect -195 5151 -161 5185
rect -195 5083 -161 5117
rect -195 5015 -161 5049
rect -195 4947 -161 4981
rect -195 4879 -161 4913
rect -195 4811 -161 4845
rect -195 4743 -161 4777
rect -195 4675 -161 4709
rect -195 4607 -161 4641
rect -195 4539 -161 4573
rect -195 4471 -161 4505
rect -195 4403 -161 4437
rect -195 4335 -161 4369
rect -195 4267 -161 4301
rect -195 4199 -161 4233
rect -195 4131 -161 4165
rect -195 4063 -161 4097
rect -195 3995 -161 4029
rect -195 3927 -161 3961
rect -195 3859 -161 3893
rect -195 3791 -161 3825
rect -195 3723 -161 3757
rect -195 3655 -161 3689
rect -195 3587 -161 3621
rect -195 3519 -161 3553
rect -195 3451 -161 3485
rect -195 3383 -161 3417
rect -195 3315 -161 3349
rect -195 3247 -161 3281
rect -195 3179 -161 3213
rect -195 3111 -161 3145
rect -195 3043 -161 3077
rect -195 2975 -161 3009
rect -195 2907 -161 2941
rect -195 2839 -161 2873
rect -195 2771 -161 2805
rect -195 2703 -161 2737
rect -195 2635 -161 2669
rect -195 2567 -161 2601
rect -195 2499 -161 2533
rect -195 2431 -161 2465
rect -195 2363 -161 2397
rect -195 2295 -161 2329
rect -195 2227 -161 2261
rect -195 2159 -161 2193
rect -195 2091 -161 2125
rect -195 2023 -161 2057
rect -195 1955 -161 1989
rect -195 1887 -161 1921
rect -195 1819 -161 1853
rect -195 1751 -161 1785
rect -195 1683 -161 1717
rect -195 1615 -161 1649
rect -195 1547 -161 1581
rect -195 1479 -161 1513
rect -195 1411 -161 1445
rect -195 1343 -161 1377
rect -195 1275 -161 1309
rect -195 1207 -161 1241
rect -195 1139 -161 1173
rect -195 1071 -161 1105
rect -195 1003 -161 1037
rect -195 935 -161 969
rect -195 867 -161 901
rect -195 799 -161 833
rect -195 731 -161 765
rect -195 663 -161 697
rect -195 595 -161 629
rect -195 527 -161 561
rect -195 459 -161 493
rect -195 391 -161 425
rect -195 323 -161 357
rect -195 255 -161 289
rect -195 187 -161 221
rect -195 119 -161 153
rect -195 51 -161 85
rect -195 -17 -161 17
rect -195 -85 -161 -51
rect -195 -153 -161 -119
rect -195 -221 -161 -187
rect -195 -289 -161 -255
rect -195 -357 -161 -323
rect -195 -425 -161 -391
rect -195 -493 -161 -459
rect -195 -561 -161 -527
rect -195 -629 -161 -595
rect -195 -697 -161 -663
rect -195 -765 -161 -731
rect -195 -833 -161 -799
rect -195 -901 -161 -867
rect -195 -969 -161 -935
rect -195 -1037 -161 -1003
rect -195 -1105 -161 -1071
rect -195 -1173 -161 -1139
rect -195 -1241 -161 -1207
rect -195 -1309 -161 -1275
rect -195 -1377 -161 -1343
rect -195 -1445 -161 -1411
rect -195 -1513 -161 -1479
rect -195 -1581 -161 -1547
rect -195 -1649 -161 -1615
rect -195 -1717 -161 -1683
rect -195 -1785 -161 -1751
rect -195 -1853 -161 -1819
rect -195 -1921 -161 -1887
rect -195 -1989 -161 -1955
rect -195 -2057 -161 -2023
rect -195 -2125 -161 -2091
rect -195 -2193 -161 -2159
rect -195 -2261 -161 -2227
rect -195 -2329 -161 -2295
rect -195 -2397 -161 -2363
rect -195 -2465 -161 -2431
rect -195 -2533 -161 -2499
rect -195 -2601 -161 -2567
rect -195 -2669 -161 -2635
rect -195 -2737 -161 -2703
rect -195 -2805 -161 -2771
rect -195 -2873 -161 -2839
rect -195 -2941 -161 -2907
rect -195 -3009 -161 -2975
rect -195 -3077 -161 -3043
rect -195 -3145 -161 -3111
rect -195 -3213 -161 -3179
rect -195 -3281 -161 -3247
rect -195 -3349 -161 -3315
rect -195 -3417 -161 -3383
rect -195 -3485 -161 -3451
rect -195 -3553 -161 -3519
rect -195 -3621 -161 -3587
rect -195 -3689 -161 -3655
rect -195 -3757 -161 -3723
rect -195 -3825 -161 -3791
rect -195 -3893 -161 -3859
rect -195 -3961 -161 -3927
rect -195 -4029 -161 -3995
rect -195 -4097 -161 -4063
rect -195 -4165 -161 -4131
rect -195 -4233 -161 -4199
rect -195 -4301 -161 -4267
rect -195 -4369 -161 -4335
rect -195 -4437 -161 -4403
rect -195 -4505 -161 -4471
rect -195 -4573 -161 -4539
rect -195 -4641 -161 -4607
rect -195 -4709 -161 -4675
rect -195 -4777 -161 -4743
rect -195 -4845 -161 -4811
rect -195 -4913 -161 -4879
rect -195 -4981 -161 -4947
rect -195 -5049 -161 -5015
rect -195 -5117 -161 -5083
rect -195 -5185 -161 -5151
rect -195 -5253 -161 -5219
rect -195 -5321 -161 -5287
rect -195 -5389 -161 -5355
rect -195 -5457 -161 -5423
rect -195 -5525 -161 -5491
rect -195 -5593 -161 -5559
rect -195 -5661 -161 -5627
rect -195 -5729 -161 -5695
rect -195 -5797 -161 -5763
rect -195 -5865 -161 -5831
rect -195 -5933 -161 -5899
rect -195 -6001 -161 -5967
rect -195 -6069 -161 -6035
rect -195 -6137 -161 -6103
rect -195 -6205 -161 -6171
rect -195 -6273 -161 -6239
rect -195 -6341 -161 -6307
rect -195 -6409 -161 -6375
rect -195 -6477 -161 -6443
rect -195 -6545 -161 -6511
rect -195 -6613 -161 -6579
rect -195 -6681 -161 -6647
rect -195 -6749 -161 -6715
rect -195 -6817 -161 -6783
rect -195 -6885 -161 -6851
rect -195 -6953 -161 -6919
rect -195 -7021 -161 -6987
rect -195 -7089 -161 -7055
rect -195 -7157 -161 -7123
rect -195 -7225 -161 -7191
rect -195 -7293 -161 -7259
rect -195 -7361 -161 -7327
rect -195 -7429 -161 -7395
rect -195 -7497 -161 -7463
rect -195 -7565 -161 -7531
rect -195 -7633 -161 -7599
rect -195 -7701 -161 -7667
rect -195 -7769 -161 -7735
rect -195 -7837 -161 -7803
rect -195 -7905 -161 -7871
rect -195 -7973 -161 -7939
rect 161 7939 195 7973
rect 161 7871 195 7905
rect 161 7803 195 7837
rect 161 7735 195 7769
rect 161 7667 195 7701
rect 161 7599 195 7633
rect 161 7531 195 7565
rect 161 7463 195 7497
rect 161 7395 195 7429
rect 161 7327 195 7361
rect 161 7259 195 7293
rect 161 7191 195 7225
rect 161 7123 195 7157
rect 161 7055 195 7089
rect 161 6987 195 7021
rect 161 6919 195 6953
rect 161 6851 195 6885
rect 161 6783 195 6817
rect 161 6715 195 6749
rect 161 6647 195 6681
rect 161 6579 195 6613
rect 161 6511 195 6545
rect 161 6443 195 6477
rect 161 6375 195 6409
rect 161 6307 195 6341
rect 161 6239 195 6273
rect 161 6171 195 6205
rect 161 6103 195 6137
rect 161 6035 195 6069
rect 161 5967 195 6001
rect 161 5899 195 5933
rect 161 5831 195 5865
rect 161 5763 195 5797
rect 161 5695 195 5729
rect 161 5627 195 5661
rect 161 5559 195 5593
rect 161 5491 195 5525
rect 161 5423 195 5457
rect 161 5355 195 5389
rect 161 5287 195 5321
rect 161 5219 195 5253
rect 161 5151 195 5185
rect 161 5083 195 5117
rect 161 5015 195 5049
rect 161 4947 195 4981
rect 161 4879 195 4913
rect 161 4811 195 4845
rect 161 4743 195 4777
rect 161 4675 195 4709
rect 161 4607 195 4641
rect 161 4539 195 4573
rect 161 4471 195 4505
rect 161 4403 195 4437
rect 161 4335 195 4369
rect 161 4267 195 4301
rect 161 4199 195 4233
rect 161 4131 195 4165
rect 161 4063 195 4097
rect 161 3995 195 4029
rect 161 3927 195 3961
rect 161 3859 195 3893
rect 161 3791 195 3825
rect 161 3723 195 3757
rect 161 3655 195 3689
rect 161 3587 195 3621
rect 161 3519 195 3553
rect 161 3451 195 3485
rect 161 3383 195 3417
rect 161 3315 195 3349
rect 161 3247 195 3281
rect 161 3179 195 3213
rect 161 3111 195 3145
rect 161 3043 195 3077
rect 161 2975 195 3009
rect 161 2907 195 2941
rect 161 2839 195 2873
rect 161 2771 195 2805
rect 161 2703 195 2737
rect 161 2635 195 2669
rect 161 2567 195 2601
rect 161 2499 195 2533
rect 161 2431 195 2465
rect 161 2363 195 2397
rect 161 2295 195 2329
rect 161 2227 195 2261
rect 161 2159 195 2193
rect 161 2091 195 2125
rect 161 2023 195 2057
rect 161 1955 195 1989
rect 161 1887 195 1921
rect 161 1819 195 1853
rect 161 1751 195 1785
rect 161 1683 195 1717
rect 161 1615 195 1649
rect 161 1547 195 1581
rect 161 1479 195 1513
rect 161 1411 195 1445
rect 161 1343 195 1377
rect 161 1275 195 1309
rect 161 1207 195 1241
rect 161 1139 195 1173
rect 161 1071 195 1105
rect 161 1003 195 1037
rect 161 935 195 969
rect 161 867 195 901
rect 161 799 195 833
rect 161 731 195 765
rect 161 663 195 697
rect 161 595 195 629
rect 161 527 195 561
rect 161 459 195 493
rect 161 391 195 425
rect 161 323 195 357
rect 161 255 195 289
rect 161 187 195 221
rect 161 119 195 153
rect 161 51 195 85
rect 161 -17 195 17
rect 161 -85 195 -51
rect 161 -153 195 -119
rect 161 -221 195 -187
rect 161 -289 195 -255
rect 161 -357 195 -323
rect 161 -425 195 -391
rect 161 -493 195 -459
rect 161 -561 195 -527
rect 161 -629 195 -595
rect 161 -697 195 -663
rect 161 -765 195 -731
rect 161 -833 195 -799
rect 161 -901 195 -867
rect 161 -969 195 -935
rect 161 -1037 195 -1003
rect 161 -1105 195 -1071
rect 161 -1173 195 -1139
rect 161 -1241 195 -1207
rect 161 -1309 195 -1275
rect 161 -1377 195 -1343
rect 161 -1445 195 -1411
rect 161 -1513 195 -1479
rect 161 -1581 195 -1547
rect 161 -1649 195 -1615
rect 161 -1717 195 -1683
rect 161 -1785 195 -1751
rect 161 -1853 195 -1819
rect 161 -1921 195 -1887
rect 161 -1989 195 -1955
rect 161 -2057 195 -2023
rect 161 -2125 195 -2091
rect 161 -2193 195 -2159
rect 161 -2261 195 -2227
rect 161 -2329 195 -2295
rect 161 -2397 195 -2363
rect 161 -2465 195 -2431
rect 161 -2533 195 -2499
rect 161 -2601 195 -2567
rect 161 -2669 195 -2635
rect 161 -2737 195 -2703
rect 161 -2805 195 -2771
rect 161 -2873 195 -2839
rect 161 -2941 195 -2907
rect 161 -3009 195 -2975
rect 161 -3077 195 -3043
rect 161 -3145 195 -3111
rect 161 -3213 195 -3179
rect 161 -3281 195 -3247
rect 161 -3349 195 -3315
rect 161 -3417 195 -3383
rect 161 -3485 195 -3451
rect 161 -3553 195 -3519
rect 161 -3621 195 -3587
rect 161 -3689 195 -3655
rect 161 -3757 195 -3723
rect 161 -3825 195 -3791
rect 161 -3893 195 -3859
rect 161 -3961 195 -3927
rect 161 -4029 195 -3995
rect 161 -4097 195 -4063
rect 161 -4165 195 -4131
rect 161 -4233 195 -4199
rect 161 -4301 195 -4267
rect 161 -4369 195 -4335
rect 161 -4437 195 -4403
rect 161 -4505 195 -4471
rect 161 -4573 195 -4539
rect 161 -4641 195 -4607
rect 161 -4709 195 -4675
rect 161 -4777 195 -4743
rect 161 -4845 195 -4811
rect 161 -4913 195 -4879
rect 161 -4981 195 -4947
rect 161 -5049 195 -5015
rect 161 -5117 195 -5083
rect 161 -5185 195 -5151
rect 161 -5253 195 -5219
rect 161 -5321 195 -5287
rect 161 -5389 195 -5355
rect 161 -5457 195 -5423
rect 161 -5525 195 -5491
rect 161 -5593 195 -5559
rect 161 -5661 195 -5627
rect 161 -5729 195 -5695
rect 161 -5797 195 -5763
rect 161 -5865 195 -5831
rect 161 -5933 195 -5899
rect 161 -6001 195 -5967
rect 161 -6069 195 -6035
rect 161 -6137 195 -6103
rect 161 -6205 195 -6171
rect 161 -6273 195 -6239
rect 161 -6341 195 -6307
rect 161 -6409 195 -6375
rect 161 -6477 195 -6443
rect 161 -6545 195 -6511
rect 161 -6613 195 -6579
rect 161 -6681 195 -6647
rect 161 -6749 195 -6715
rect 161 -6817 195 -6783
rect 161 -6885 195 -6851
rect 161 -6953 195 -6919
rect 161 -7021 195 -6987
rect 161 -7089 195 -7055
rect 161 -7157 195 -7123
rect 161 -7225 195 -7191
rect 161 -7293 195 -7259
rect 161 -7361 195 -7327
rect 161 -7429 195 -7395
rect 161 -7497 195 -7463
rect 161 -7565 195 -7531
rect 161 -7633 195 -7599
rect 161 -7701 195 -7667
rect 161 -7769 195 -7735
rect 161 -7837 195 -7803
rect 161 -7905 195 -7871
rect 161 -7973 195 -7939
rect -195 -8041 -161 -8007
rect -195 -8140 -161 -8075
rect 161 -8041 195 -8007
rect 161 -8140 195 -8075
rect -195 -8174 -85 -8140
rect -51 -8174 -17 -8140
rect 17 -8174 51 -8140
rect 85 -8174 195 -8140
<< psubdiffcont >>
rect -85 8140 -51 8174
rect -17 8140 17 8174
rect 51 8140 85 8174
rect -195 8041 -161 8075
rect -195 7973 -161 8007
rect 161 8041 195 8075
rect -195 7905 -161 7939
rect -195 7837 -161 7871
rect -195 7769 -161 7803
rect -195 7701 -161 7735
rect -195 7633 -161 7667
rect -195 7565 -161 7599
rect -195 7497 -161 7531
rect -195 7429 -161 7463
rect -195 7361 -161 7395
rect -195 7293 -161 7327
rect -195 7225 -161 7259
rect -195 7157 -161 7191
rect -195 7089 -161 7123
rect -195 7021 -161 7055
rect -195 6953 -161 6987
rect -195 6885 -161 6919
rect -195 6817 -161 6851
rect -195 6749 -161 6783
rect -195 6681 -161 6715
rect -195 6613 -161 6647
rect -195 6545 -161 6579
rect -195 6477 -161 6511
rect -195 6409 -161 6443
rect -195 6341 -161 6375
rect -195 6273 -161 6307
rect -195 6205 -161 6239
rect -195 6137 -161 6171
rect -195 6069 -161 6103
rect -195 6001 -161 6035
rect -195 5933 -161 5967
rect -195 5865 -161 5899
rect -195 5797 -161 5831
rect -195 5729 -161 5763
rect -195 5661 -161 5695
rect -195 5593 -161 5627
rect -195 5525 -161 5559
rect -195 5457 -161 5491
rect -195 5389 -161 5423
rect -195 5321 -161 5355
rect -195 5253 -161 5287
rect -195 5185 -161 5219
rect -195 5117 -161 5151
rect -195 5049 -161 5083
rect -195 4981 -161 5015
rect -195 4913 -161 4947
rect -195 4845 -161 4879
rect -195 4777 -161 4811
rect -195 4709 -161 4743
rect -195 4641 -161 4675
rect -195 4573 -161 4607
rect -195 4505 -161 4539
rect -195 4437 -161 4471
rect -195 4369 -161 4403
rect -195 4301 -161 4335
rect -195 4233 -161 4267
rect -195 4165 -161 4199
rect -195 4097 -161 4131
rect -195 4029 -161 4063
rect -195 3961 -161 3995
rect -195 3893 -161 3927
rect -195 3825 -161 3859
rect -195 3757 -161 3791
rect -195 3689 -161 3723
rect -195 3621 -161 3655
rect -195 3553 -161 3587
rect -195 3485 -161 3519
rect -195 3417 -161 3451
rect -195 3349 -161 3383
rect -195 3281 -161 3315
rect -195 3213 -161 3247
rect -195 3145 -161 3179
rect -195 3077 -161 3111
rect -195 3009 -161 3043
rect -195 2941 -161 2975
rect -195 2873 -161 2907
rect -195 2805 -161 2839
rect -195 2737 -161 2771
rect -195 2669 -161 2703
rect -195 2601 -161 2635
rect -195 2533 -161 2567
rect -195 2465 -161 2499
rect -195 2397 -161 2431
rect -195 2329 -161 2363
rect -195 2261 -161 2295
rect -195 2193 -161 2227
rect -195 2125 -161 2159
rect -195 2057 -161 2091
rect -195 1989 -161 2023
rect -195 1921 -161 1955
rect -195 1853 -161 1887
rect -195 1785 -161 1819
rect -195 1717 -161 1751
rect -195 1649 -161 1683
rect -195 1581 -161 1615
rect -195 1513 -161 1547
rect -195 1445 -161 1479
rect -195 1377 -161 1411
rect -195 1309 -161 1343
rect -195 1241 -161 1275
rect -195 1173 -161 1207
rect -195 1105 -161 1139
rect -195 1037 -161 1071
rect -195 969 -161 1003
rect -195 901 -161 935
rect -195 833 -161 867
rect -195 765 -161 799
rect -195 697 -161 731
rect -195 629 -161 663
rect -195 561 -161 595
rect -195 493 -161 527
rect -195 425 -161 459
rect -195 357 -161 391
rect -195 289 -161 323
rect -195 221 -161 255
rect -195 153 -161 187
rect -195 85 -161 119
rect -195 17 -161 51
rect -195 -51 -161 -17
rect -195 -119 -161 -85
rect -195 -187 -161 -153
rect -195 -255 -161 -221
rect -195 -323 -161 -289
rect -195 -391 -161 -357
rect -195 -459 -161 -425
rect -195 -527 -161 -493
rect -195 -595 -161 -561
rect -195 -663 -161 -629
rect -195 -731 -161 -697
rect -195 -799 -161 -765
rect -195 -867 -161 -833
rect -195 -935 -161 -901
rect -195 -1003 -161 -969
rect -195 -1071 -161 -1037
rect -195 -1139 -161 -1105
rect -195 -1207 -161 -1173
rect -195 -1275 -161 -1241
rect -195 -1343 -161 -1309
rect -195 -1411 -161 -1377
rect -195 -1479 -161 -1445
rect -195 -1547 -161 -1513
rect -195 -1615 -161 -1581
rect -195 -1683 -161 -1649
rect -195 -1751 -161 -1717
rect -195 -1819 -161 -1785
rect -195 -1887 -161 -1853
rect -195 -1955 -161 -1921
rect -195 -2023 -161 -1989
rect -195 -2091 -161 -2057
rect -195 -2159 -161 -2125
rect -195 -2227 -161 -2193
rect -195 -2295 -161 -2261
rect -195 -2363 -161 -2329
rect -195 -2431 -161 -2397
rect -195 -2499 -161 -2465
rect -195 -2567 -161 -2533
rect -195 -2635 -161 -2601
rect -195 -2703 -161 -2669
rect -195 -2771 -161 -2737
rect -195 -2839 -161 -2805
rect -195 -2907 -161 -2873
rect -195 -2975 -161 -2941
rect -195 -3043 -161 -3009
rect -195 -3111 -161 -3077
rect -195 -3179 -161 -3145
rect -195 -3247 -161 -3213
rect -195 -3315 -161 -3281
rect -195 -3383 -161 -3349
rect -195 -3451 -161 -3417
rect -195 -3519 -161 -3485
rect -195 -3587 -161 -3553
rect -195 -3655 -161 -3621
rect -195 -3723 -161 -3689
rect -195 -3791 -161 -3757
rect -195 -3859 -161 -3825
rect -195 -3927 -161 -3893
rect -195 -3995 -161 -3961
rect -195 -4063 -161 -4029
rect -195 -4131 -161 -4097
rect -195 -4199 -161 -4165
rect -195 -4267 -161 -4233
rect -195 -4335 -161 -4301
rect -195 -4403 -161 -4369
rect -195 -4471 -161 -4437
rect -195 -4539 -161 -4505
rect -195 -4607 -161 -4573
rect -195 -4675 -161 -4641
rect -195 -4743 -161 -4709
rect -195 -4811 -161 -4777
rect -195 -4879 -161 -4845
rect -195 -4947 -161 -4913
rect -195 -5015 -161 -4981
rect -195 -5083 -161 -5049
rect -195 -5151 -161 -5117
rect -195 -5219 -161 -5185
rect -195 -5287 -161 -5253
rect -195 -5355 -161 -5321
rect -195 -5423 -161 -5389
rect -195 -5491 -161 -5457
rect -195 -5559 -161 -5525
rect -195 -5627 -161 -5593
rect -195 -5695 -161 -5661
rect -195 -5763 -161 -5729
rect -195 -5831 -161 -5797
rect -195 -5899 -161 -5865
rect -195 -5967 -161 -5933
rect -195 -6035 -161 -6001
rect -195 -6103 -161 -6069
rect -195 -6171 -161 -6137
rect -195 -6239 -161 -6205
rect -195 -6307 -161 -6273
rect -195 -6375 -161 -6341
rect -195 -6443 -161 -6409
rect -195 -6511 -161 -6477
rect -195 -6579 -161 -6545
rect -195 -6647 -161 -6613
rect -195 -6715 -161 -6681
rect -195 -6783 -161 -6749
rect -195 -6851 -161 -6817
rect -195 -6919 -161 -6885
rect -195 -6987 -161 -6953
rect -195 -7055 -161 -7021
rect -195 -7123 -161 -7089
rect -195 -7191 -161 -7157
rect -195 -7259 -161 -7225
rect -195 -7327 -161 -7293
rect -195 -7395 -161 -7361
rect -195 -7463 -161 -7429
rect -195 -7531 -161 -7497
rect -195 -7599 -161 -7565
rect -195 -7667 -161 -7633
rect -195 -7735 -161 -7701
rect -195 -7803 -161 -7769
rect -195 -7871 -161 -7837
rect -195 -7939 -161 -7905
rect -195 -8007 -161 -7973
rect 161 7973 195 8007
rect 161 7905 195 7939
rect 161 7837 195 7871
rect 161 7769 195 7803
rect 161 7701 195 7735
rect 161 7633 195 7667
rect 161 7565 195 7599
rect 161 7497 195 7531
rect 161 7429 195 7463
rect 161 7361 195 7395
rect 161 7293 195 7327
rect 161 7225 195 7259
rect 161 7157 195 7191
rect 161 7089 195 7123
rect 161 7021 195 7055
rect 161 6953 195 6987
rect 161 6885 195 6919
rect 161 6817 195 6851
rect 161 6749 195 6783
rect 161 6681 195 6715
rect 161 6613 195 6647
rect 161 6545 195 6579
rect 161 6477 195 6511
rect 161 6409 195 6443
rect 161 6341 195 6375
rect 161 6273 195 6307
rect 161 6205 195 6239
rect 161 6137 195 6171
rect 161 6069 195 6103
rect 161 6001 195 6035
rect 161 5933 195 5967
rect 161 5865 195 5899
rect 161 5797 195 5831
rect 161 5729 195 5763
rect 161 5661 195 5695
rect 161 5593 195 5627
rect 161 5525 195 5559
rect 161 5457 195 5491
rect 161 5389 195 5423
rect 161 5321 195 5355
rect 161 5253 195 5287
rect 161 5185 195 5219
rect 161 5117 195 5151
rect 161 5049 195 5083
rect 161 4981 195 5015
rect 161 4913 195 4947
rect 161 4845 195 4879
rect 161 4777 195 4811
rect 161 4709 195 4743
rect 161 4641 195 4675
rect 161 4573 195 4607
rect 161 4505 195 4539
rect 161 4437 195 4471
rect 161 4369 195 4403
rect 161 4301 195 4335
rect 161 4233 195 4267
rect 161 4165 195 4199
rect 161 4097 195 4131
rect 161 4029 195 4063
rect 161 3961 195 3995
rect 161 3893 195 3927
rect 161 3825 195 3859
rect 161 3757 195 3791
rect 161 3689 195 3723
rect 161 3621 195 3655
rect 161 3553 195 3587
rect 161 3485 195 3519
rect 161 3417 195 3451
rect 161 3349 195 3383
rect 161 3281 195 3315
rect 161 3213 195 3247
rect 161 3145 195 3179
rect 161 3077 195 3111
rect 161 3009 195 3043
rect 161 2941 195 2975
rect 161 2873 195 2907
rect 161 2805 195 2839
rect 161 2737 195 2771
rect 161 2669 195 2703
rect 161 2601 195 2635
rect 161 2533 195 2567
rect 161 2465 195 2499
rect 161 2397 195 2431
rect 161 2329 195 2363
rect 161 2261 195 2295
rect 161 2193 195 2227
rect 161 2125 195 2159
rect 161 2057 195 2091
rect 161 1989 195 2023
rect 161 1921 195 1955
rect 161 1853 195 1887
rect 161 1785 195 1819
rect 161 1717 195 1751
rect 161 1649 195 1683
rect 161 1581 195 1615
rect 161 1513 195 1547
rect 161 1445 195 1479
rect 161 1377 195 1411
rect 161 1309 195 1343
rect 161 1241 195 1275
rect 161 1173 195 1207
rect 161 1105 195 1139
rect 161 1037 195 1071
rect 161 969 195 1003
rect 161 901 195 935
rect 161 833 195 867
rect 161 765 195 799
rect 161 697 195 731
rect 161 629 195 663
rect 161 561 195 595
rect 161 493 195 527
rect 161 425 195 459
rect 161 357 195 391
rect 161 289 195 323
rect 161 221 195 255
rect 161 153 195 187
rect 161 85 195 119
rect 161 17 195 51
rect 161 -51 195 -17
rect 161 -119 195 -85
rect 161 -187 195 -153
rect 161 -255 195 -221
rect 161 -323 195 -289
rect 161 -391 195 -357
rect 161 -459 195 -425
rect 161 -527 195 -493
rect 161 -595 195 -561
rect 161 -663 195 -629
rect 161 -731 195 -697
rect 161 -799 195 -765
rect 161 -867 195 -833
rect 161 -935 195 -901
rect 161 -1003 195 -969
rect 161 -1071 195 -1037
rect 161 -1139 195 -1105
rect 161 -1207 195 -1173
rect 161 -1275 195 -1241
rect 161 -1343 195 -1309
rect 161 -1411 195 -1377
rect 161 -1479 195 -1445
rect 161 -1547 195 -1513
rect 161 -1615 195 -1581
rect 161 -1683 195 -1649
rect 161 -1751 195 -1717
rect 161 -1819 195 -1785
rect 161 -1887 195 -1853
rect 161 -1955 195 -1921
rect 161 -2023 195 -1989
rect 161 -2091 195 -2057
rect 161 -2159 195 -2125
rect 161 -2227 195 -2193
rect 161 -2295 195 -2261
rect 161 -2363 195 -2329
rect 161 -2431 195 -2397
rect 161 -2499 195 -2465
rect 161 -2567 195 -2533
rect 161 -2635 195 -2601
rect 161 -2703 195 -2669
rect 161 -2771 195 -2737
rect 161 -2839 195 -2805
rect 161 -2907 195 -2873
rect 161 -2975 195 -2941
rect 161 -3043 195 -3009
rect 161 -3111 195 -3077
rect 161 -3179 195 -3145
rect 161 -3247 195 -3213
rect 161 -3315 195 -3281
rect 161 -3383 195 -3349
rect 161 -3451 195 -3417
rect 161 -3519 195 -3485
rect 161 -3587 195 -3553
rect 161 -3655 195 -3621
rect 161 -3723 195 -3689
rect 161 -3791 195 -3757
rect 161 -3859 195 -3825
rect 161 -3927 195 -3893
rect 161 -3995 195 -3961
rect 161 -4063 195 -4029
rect 161 -4131 195 -4097
rect 161 -4199 195 -4165
rect 161 -4267 195 -4233
rect 161 -4335 195 -4301
rect 161 -4403 195 -4369
rect 161 -4471 195 -4437
rect 161 -4539 195 -4505
rect 161 -4607 195 -4573
rect 161 -4675 195 -4641
rect 161 -4743 195 -4709
rect 161 -4811 195 -4777
rect 161 -4879 195 -4845
rect 161 -4947 195 -4913
rect 161 -5015 195 -4981
rect 161 -5083 195 -5049
rect 161 -5151 195 -5117
rect 161 -5219 195 -5185
rect 161 -5287 195 -5253
rect 161 -5355 195 -5321
rect 161 -5423 195 -5389
rect 161 -5491 195 -5457
rect 161 -5559 195 -5525
rect 161 -5627 195 -5593
rect 161 -5695 195 -5661
rect 161 -5763 195 -5729
rect 161 -5831 195 -5797
rect 161 -5899 195 -5865
rect 161 -5967 195 -5933
rect 161 -6035 195 -6001
rect 161 -6103 195 -6069
rect 161 -6171 195 -6137
rect 161 -6239 195 -6205
rect 161 -6307 195 -6273
rect 161 -6375 195 -6341
rect 161 -6443 195 -6409
rect 161 -6511 195 -6477
rect 161 -6579 195 -6545
rect 161 -6647 195 -6613
rect 161 -6715 195 -6681
rect 161 -6783 195 -6749
rect 161 -6851 195 -6817
rect 161 -6919 195 -6885
rect 161 -6987 195 -6953
rect 161 -7055 195 -7021
rect 161 -7123 195 -7089
rect 161 -7191 195 -7157
rect 161 -7259 195 -7225
rect 161 -7327 195 -7293
rect 161 -7395 195 -7361
rect 161 -7463 195 -7429
rect 161 -7531 195 -7497
rect 161 -7599 195 -7565
rect 161 -7667 195 -7633
rect 161 -7735 195 -7701
rect 161 -7803 195 -7769
rect 161 -7871 195 -7837
rect 161 -7939 195 -7905
rect -195 -8075 -161 -8041
rect 161 -8007 195 -7973
rect 161 -8075 195 -8041
rect -85 -8174 -51 -8140
rect -17 -8174 17 -8140
rect 51 -8174 85 -8140
<< poly >>
rect -35 8072 35 8088
rect -35 8038 -17 8072
rect 17 8038 35 8072
rect -35 8000 35 8038
rect -35 -8038 35 -8000
rect -35 -8072 -17 -8038
rect 17 -8072 35 -8038
rect -35 -8088 35 -8072
<< polycont >>
rect -17 8038 17 8072
rect -17 -8072 17 -8038
<< locali >>
rect -195 8140 -85 8174
rect -51 8140 -17 8174
rect 17 8140 51 8174
rect 85 8140 195 8174
rect -195 8075 -161 8140
rect 161 8075 195 8140
rect -195 8007 -161 8041
rect -35 8038 -17 8072
rect 17 8038 35 8072
rect 161 8007 195 8041
rect -195 7939 -161 7973
rect -195 7871 -161 7905
rect -195 7803 -161 7837
rect -195 7735 -161 7769
rect -195 7667 -161 7701
rect -195 7599 -161 7633
rect -195 7531 -161 7565
rect -195 7463 -161 7497
rect -195 7395 -161 7429
rect -195 7327 -161 7361
rect -195 7259 -161 7293
rect -195 7191 -161 7225
rect -195 7123 -161 7157
rect -195 7055 -161 7089
rect -195 6987 -161 7021
rect -195 6919 -161 6953
rect -195 6851 -161 6885
rect -195 6783 -161 6817
rect -195 6715 -161 6749
rect -195 6647 -161 6681
rect -195 6579 -161 6613
rect -195 6511 -161 6545
rect -195 6443 -161 6477
rect -195 6375 -161 6409
rect -195 6307 -161 6341
rect -195 6239 -161 6273
rect -195 6171 -161 6205
rect -195 6103 -161 6137
rect -195 6035 -161 6069
rect -195 5967 -161 6001
rect -195 5899 -161 5933
rect -195 5831 -161 5865
rect -195 5763 -161 5797
rect -195 5695 -161 5729
rect -195 5627 -161 5661
rect -195 5559 -161 5593
rect -195 5491 -161 5525
rect -195 5423 -161 5457
rect -195 5355 -161 5389
rect -195 5287 -161 5321
rect -195 5219 -161 5253
rect -195 5151 -161 5185
rect -195 5083 -161 5117
rect -195 5015 -161 5049
rect -195 4947 -161 4981
rect -195 4879 -161 4913
rect -195 4811 -161 4845
rect -195 4743 -161 4777
rect -195 4675 -161 4709
rect -195 4607 -161 4641
rect -195 4539 -161 4573
rect -195 4471 -161 4505
rect -195 4403 -161 4437
rect -195 4335 -161 4369
rect -195 4267 -161 4301
rect -195 4199 -161 4233
rect -195 4131 -161 4165
rect -195 4063 -161 4097
rect -195 3995 -161 4029
rect -195 3927 -161 3961
rect -195 3859 -161 3893
rect -195 3791 -161 3825
rect -195 3723 -161 3757
rect -195 3655 -161 3689
rect -195 3587 -161 3621
rect -195 3519 -161 3553
rect -195 3451 -161 3485
rect -195 3383 -161 3417
rect -195 3315 -161 3349
rect -195 3247 -161 3281
rect -195 3179 -161 3213
rect -195 3111 -161 3145
rect -195 3043 -161 3077
rect -195 2975 -161 3009
rect -195 2907 -161 2941
rect -195 2839 -161 2873
rect -195 2771 -161 2805
rect -195 2703 -161 2737
rect -195 2635 -161 2669
rect -195 2567 -161 2601
rect -195 2499 -161 2533
rect -195 2431 -161 2465
rect -195 2363 -161 2397
rect -195 2295 -161 2329
rect -195 2227 -161 2261
rect -195 2159 -161 2193
rect -195 2091 -161 2125
rect -195 2023 -161 2057
rect -195 1955 -161 1989
rect -195 1887 -161 1921
rect -195 1819 -161 1853
rect -195 1751 -161 1785
rect -195 1683 -161 1717
rect -195 1615 -161 1649
rect -195 1547 -161 1581
rect -195 1479 -161 1513
rect -195 1411 -161 1445
rect -195 1343 -161 1377
rect -195 1275 -161 1309
rect -195 1207 -161 1241
rect -195 1139 -161 1173
rect -195 1071 -161 1105
rect -195 1003 -161 1037
rect -195 935 -161 969
rect -195 867 -161 901
rect -195 799 -161 833
rect -195 731 -161 765
rect -195 663 -161 697
rect -195 595 -161 629
rect -195 527 -161 561
rect -195 459 -161 493
rect -195 391 -161 425
rect -195 323 -161 357
rect -195 255 -161 289
rect -195 187 -161 221
rect -195 119 -161 153
rect -195 51 -161 85
rect -195 -17 -161 17
rect -195 -85 -161 -51
rect -195 -153 -161 -119
rect -195 -221 -161 -187
rect -195 -289 -161 -255
rect -195 -357 -161 -323
rect -195 -425 -161 -391
rect -195 -493 -161 -459
rect -195 -561 -161 -527
rect -195 -629 -161 -595
rect -195 -697 -161 -663
rect -195 -765 -161 -731
rect -195 -833 -161 -799
rect -195 -901 -161 -867
rect -195 -969 -161 -935
rect -195 -1037 -161 -1003
rect -195 -1105 -161 -1071
rect -195 -1173 -161 -1139
rect -195 -1241 -161 -1207
rect -195 -1309 -161 -1275
rect -195 -1377 -161 -1343
rect -195 -1445 -161 -1411
rect -195 -1513 -161 -1479
rect -195 -1581 -161 -1547
rect -195 -1649 -161 -1615
rect -195 -1717 -161 -1683
rect -195 -1785 -161 -1751
rect -195 -1853 -161 -1819
rect -195 -1921 -161 -1887
rect -195 -1989 -161 -1955
rect -195 -2057 -161 -2023
rect -195 -2125 -161 -2091
rect -195 -2193 -161 -2159
rect -195 -2261 -161 -2227
rect -195 -2329 -161 -2295
rect -195 -2397 -161 -2363
rect -195 -2465 -161 -2431
rect -195 -2533 -161 -2499
rect -195 -2601 -161 -2567
rect -195 -2669 -161 -2635
rect -195 -2737 -161 -2703
rect -195 -2805 -161 -2771
rect -195 -2873 -161 -2839
rect -195 -2941 -161 -2907
rect -195 -3009 -161 -2975
rect -195 -3077 -161 -3043
rect -195 -3145 -161 -3111
rect -195 -3213 -161 -3179
rect -195 -3281 -161 -3247
rect -195 -3349 -161 -3315
rect -195 -3417 -161 -3383
rect -195 -3485 -161 -3451
rect -195 -3553 -161 -3519
rect -195 -3621 -161 -3587
rect -195 -3689 -161 -3655
rect -195 -3757 -161 -3723
rect -195 -3825 -161 -3791
rect -195 -3893 -161 -3859
rect -195 -3961 -161 -3927
rect -195 -4029 -161 -3995
rect -195 -4097 -161 -4063
rect -195 -4165 -161 -4131
rect -195 -4233 -161 -4199
rect -195 -4301 -161 -4267
rect -195 -4369 -161 -4335
rect -195 -4437 -161 -4403
rect -195 -4505 -161 -4471
rect -195 -4573 -161 -4539
rect -195 -4641 -161 -4607
rect -195 -4709 -161 -4675
rect -195 -4777 -161 -4743
rect -195 -4845 -161 -4811
rect -195 -4913 -161 -4879
rect -195 -4981 -161 -4947
rect -195 -5049 -161 -5015
rect -195 -5117 -161 -5083
rect -195 -5185 -161 -5151
rect -195 -5253 -161 -5219
rect -195 -5321 -161 -5287
rect -195 -5389 -161 -5355
rect -195 -5457 -161 -5423
rect -195 -5525 -161 -5491
rect -195 -5593 -161 -5559
rect -195 -5661 -161 -5627
rect -195 -5729 -161 -5695
rect -195 -5797 -161 -5763
rect -195 -5865 -161 -5831
rect -195 -5933 -161 -5899
rect -195 -6001 -161 -5967
rect -195 -6069 -161 -6035
rect -195 -6137 -161 -6103
rect -195 -6205 -161 -6171
rect -195 -6273 -161 -6239
rect -195 -6341 -161 -6307
rect -195 -6409 -161 -6375
rect -195 -6477 -161 -6443
rect -195 -6545 -161 -6511
rect -195 -6613 -161 -6579
rect -195 -6681 -161 -6647
rect -195 -6749 -161 -6715
rect -195 -6817 -161 -6783
rect -195 -6885 -161 -6851
rect -195 -6953 -161 -6919
rect -195 -7021 -161 -6987
rect -195 -7089 -161 -7055
rect -195 -7157 -161 -7123
rect -195 -7225 -161 -7191
rect -195 -7293 -161 -7259
rect -195 -7361 -161 -7327
rect -195 -7429 -161 -7395
rect -195 -7497 -161 -7463
rect -195 -7565 -161 -7531
rect -195 -7633 -161 -7599
rect -195 -7701 -161 -7667
rect -195 -7769 -161 -7735
rect -195 -7837 -161 -7803
rect -195 -7905 -161 -7871
rect -195 -7973 -161 -7939
rect -81 7973 -47 8004
rect -81 7905 -47 7939
rect -81 7837 -47 7867
rect -81 7769 -47 7795
rect -81 7701 -47 7723
rect -81 7633 -47 7651
rect -81 7565 -47 7579
rect -81 7497 -47 7507
rect -81 7429 -47 7435
rect -81 7361 -47 7363
rect -81 7325 -47 7327
rect -81 7253 -47 7259
rect -81 7181 -47 7191
rect -81 7109 -47 7123
rect -81 7037 -47 7055
rect -81 6965 -47 6987
rect -81 6893 -47 6919
rect -81 6821 -47 6851
rect -81 6749 -47 6783
rect -81 6681 -47 6715
rect -81 6613 -47 6643
rect -81 6545 -47 6571
rect -81 6477 -47 6499
rect -81 6409 -47 6427
rect -81 6341 -47 6355
rect -81 6273 -47 6283
rect -81 6205 -47 6211
rect -81 6137 -47 6139
rect -81 6101 -47 6103
rect -81 6029 -47 6035
rect -81 5957 -47 5967
rect -81 5885 -47 5899
rect -81 5813 -47 5831
rect -81 5741 -47 5763
rect -81 5669 -47 5695
rect -81 5597 -47 5627
rect -81 5525 -47 5559
rect -81 5457 -47 5491
rect -81 5389 -47 5419
rect -81 5321 -47 5347
rect -81 5253 -47 5275
rect -81 5185 -47 5203
rect -81 5117 -47 5131
rect -81 5049 -47 5059
rect -81 4981 -47 4987
rect -81 4913 -47 4915
rect -81 4877 -47 4879
rect -81 4805 -47 4811
rect -81 4733 -47 4743
rect -81 4661 -47 4675
rect -81 4589 -47 4607
rect -81 4517 -47 4539
rect -81 4445 -47 4471
rect -81 4373 -47 4403
rect -81 4301 -47 4335
rect -81 4233 -47 4267
rect -81 4165 -47 4195
rect -81 4097 -47 4123
rect -81 4029 -47 4051
rect -81 3961 -47 3979
rect -81 3893 -47 3907
rect -81 3825 -47 3835
rect -81 3757 -47 3763
rect -81 3689 -47 3691
rect -81 3653 -47 3655
rect -81 3581 -47 3587
rect -81 3509 -47 3519
rect -81 3437 -47 3451
rect -81 3365 -47 3383
rect -81 3293 -47 3315
rect -81 3221 -47 3247
rect -81 3149 -47 3179
rect -81 3077 -47 3111
rect -81 3009 -47 3043
rect -81 2941 -47 2971
rect -81 2873 -47 2899
rect -81 2805 -47 2827
rect -81 2737 -47 2755
rect -81 2669 -47 2683
rect -81 2601 -47 2611
rect -81 2533 -47 2539
rect -81 2465 -47 2467
rect -81 2429 -47 2431
rect -81 2357 -47 2363
rect -81 2285 -47 2295
rect -81 2213 -47 2227
rect -81 2141 -47 2159
rect -81 2069 -47 2091
rect -81 1997 -47 2023
rect -81 1925 -47 1955
rect -81 1853 -47 1887
rect -81 1785 -47 1819
rect -81 1717 -47 1747
rect -81 1649 -47 1675
rect -81 1581 -47 1603
rect -81 1513 -47 1531
rect -81 1445 -47 1459
rect -81 1377 -47 1387
rect -81 1309 -47 1315
rect -81 1241 -47 1243
rect -81 1205 -47 1207
rect -81 1133 -47 1139
rect -81 1061 -47 1071
rect -81 989 -47 1003
rect -81 917 -47 935
rect -81 845 -47 867
rect -81 773 -47 799
rect -81 701 -47 731
rect -81 629 -47 663
rect -81 561 -47 595
rect -81 493 -47 523
rect -81 425 -47 451
rect -81 357 -47 379
rect -81 289 -47 307
rect -81 221 -47 235
rect -81 153 -47 163
rect -81 85 -47 91
rect -81 17 -47 19
rect -81 -19 -47 -17
rect -81 -91 -47 -85
rect -81 -163 -47 -153
rect -81 -235 -47 -221
rect -81 -307 -47 -289
rect -81 -379 -47 -357
rect -81 -451 -47 -425
rect -81 -523 -47 -493
rect -81 -595 -47 -561
rect -81 -663 -47 -629
rect -81 -731 -47 -701
rect -81 -799 -47 -773
rect -81 -867 -47 -845
rect -81 -935 -47 -917
rect -81 -1003 -47 -989
rect -81 -1071 -47 -1061
rect -81 -1139 -47 -1133
rect -81 -1207 -47 -1205
rect -81 -1243 -47 -1241
rect -81 -1315 -47 -1309
rect -81 -1387 -47 -1377
rect -81 -1459 -47 -1445
rect -81 -1531 -47 -1513
rect -81 -1603 -47 -1581
rect -81 -1675 -47 -1649
rect -81 -1747 -47 -1717
rect -81 -1819 -47 -1785
rect -81 -1887 -47 -1853
rect -81 -1955 -47 -1925
rect -81 -2023 -47 -1997
rect -81 -2091 -47 -2069
rect -81 -2159 -47 -2141
rect -81 -2227 -47 -2213
rect -81 -2295 -47 -2285
rect -81 -2363 -47 -2357
rect -81 -2431 -47 -2429
rect -81 -2467 -47 -2465
rect -81 -2539 -47 -2533
rect -81 -2611 -47 -2601
rect -81 -2683 -47 -2669
rect -81 -2755 -47 -2737
rect -81 -2827 -47 -2805
rect -81 -2899 -47 -2873
rect -81 -2971 -47 -2941
rect -81 -3043 -47 -3009
rect -81 -3111 -47 -3077
rect -81 -3179 -47 -3149
rect -81 -3247 -47 -3221
rect -81 -3315 -47 -3293
rect -81 -3383 -47 -3365
rect -81 -3451 -47 -3437
rect -81 -3519 -47 -3509
rect -81 -3587 -47 -3581
rect -81 -3655 -47 -3653
rect -81 -3691 -47 -3689
rect -81 -3763 -47 -3757
rect -81 -3835 -47 -3825
rect -81 -3907 -47 -3893
rect -81 -3979 -47 -3961
rect -81 -4051 -47 -4029
rect -81 -4123 -47 -4097
rect -81 -4195 -47 -4165
rect -81 -4267 -47 -4233
rect -81 -4335 -47 -4301
rect -81 -4403 -47 -4373
rect -81 -4471 -47 -4445
rect -81 -4539 -47 -4517
rect -81 -4607 -47 -4589
rect -81 -4675 -47 -4661
rect -81 -4743 -47 -4733
rect -81 -4811 -47 -4805
rect -81 -4879 -47 -4877
rect -81 -4915 -47 -4913
rect -81 -4987 -47 -4981
rect -81 -5059 -47 -5049
rect -81 -5131 -47 -5117
rect -81 -5203 -47 -5185
rect -81 -5275 -47 -5253
rect -81 -5347 -47 -5321
rect -81 -5419 -47 -5389
rect -81 -5491 -47 -5457
rect -81 -5559 -47 -5525
rect -81 -5627 -47 -5597
rect -81 -5695 -47 -5669
rect -81 -5763 -47 -5741
rect -81 -5831 -47 -5813
rect -81 -5899 -47 -5885
rect -81 -5967 -47 -5957
rect -81 -6035 -47 -6029
rect -81 -6103 -47 -6101
rect -81 -6139 -47 -6137
rect -81 -6211 -47 -6205
rect -81 -6283 -47 -6273
rect -81 -6355 -47 -6341
rect -81 -6427 -47 -6409
rect -81 -6499 -47 -6477
rect -81 -6571 -47 -6545
rect -81 -6643 -47 -6613
rect -81 -6715 -47 -6681
rect -81 -6783 -47 -6749
rect -81 -6851 -47 -6821
rect -81 -6919 -47 -6893
rect -81 -6987 -47 -6965
rect -81 -7055 -47 -7037
rect -81 -7123 -47 -7109
rect -81 -7191 -47 -7181
rect -81 -7259 -47 -7253
rect -81 -7327 -47 -7325
rect -81 -7363 -47 -7361
rect -81 -7435 -47 -7429
rect -81 -7507 -47 -7497
rect -81 -7579 -47 -7565
rect -81 -7651 -47 -7633
rect -81 -7723 -47 -7701
rect -81 -7795 -47 -7769
rect -81 -7867 -47 -7837
rect -81 -7939 -47 -7905
rect -81 -8004 -47 -7973
rect 47 7973 81 8004
rect 47 7905 81 7939
rect 47 7837 81 7867
rect 47 7769 81 7795
rect 47 7701 81 7723
rect 47 7633 81 7651
rect 47 7565 81 7579
rect 47 7497 81 7507
rect 47 7429 81 7435
rect 47 7361 81 7363
rect 47 7325 81 7327
rect 47 7253 81 7259
rect 47 7181 81 7191
rect 47 7109 81 7123
rect 47 7037 81 7055
rect 47 6965 81 6987
rect 47 6893 81 6919
rect 47 6821 81 6851
rect 47 6749 81 6783
rect 47 6681 81 6715
rect 47 6613 81 6643
rect 47 6545 81 6571
rect 47 6477 81 6499
rect 47 6409 81 6427
rect 47 6341 81 6355
rect 47 6273 81 6283
rect 47 6205 81 6211
rect 47 6137 81 6139
rect 47 6101 81 6103
rect 47 6029 81 6035
rect 47 5957 81 5967
rect 47 5885 81 5899
rect 47 5813 81 5831
rect 47 5741 81 5763
rect 47 5669 81 5695
rect 47 5597 81 5627
rect 47 5525 81 5559
rect 47 5457 81 5491
rect 47 5389 81 5419
rect 47 5321 81 5347
rect 47 5253 81 5275
rect 47 5185 81 5203
rect 47 5117 81 5131
rect 47 5049 81 5059
rect 47 4981 81 4987
rect 47 4913 81 4915
rect 47 4877 81 4879
rect 47 4805 81 4811
rect 47 4733 81 4743
rect 47 4661 81 4675
rect 47 4589 81 4607
rect 47 4517 81 4539
rect 47 4445 81 4471
rect 47 4373 81 4403
rect 47 4301 81 4335
rect 47 4233 81 4267
rect 47 4165 81 4195
rect 47 4097 81 4123
rect 47 4029 81 4051
rect 47 3961 81 3979
rect 47 3893 81 3907
rect 47 3825 81 3835
rect 47 3757 81 3763
rect 47 3689 81 3691
rect 47 3653 81 3655
rect 47 3581 81 3587
rect 47 3509 81 3519
rect 47 3437 81 3451
rect 47 3365 81 3383
rect 47 3293 81 3315
rect 47 3221 81 3247
rect 47 3149 81 3179
rect 47 3077 81 3111
rect 47 3009 81 3043
rect 47 2941 81 2971
rect 47 2873 81 2899
rect 47 2805 81 2827
rect 47 2737 81 2755
rect 47 2669 81 2683
rect 47 2601 81 2611
rect 47 2533 81 2539
rect 47 2465 81 2467
rect 47 2429 81 2431
rect 47 2357 81 2363
rect 47 2285 81 2295
rect 47 2213 81 2227
rect 47 2141 81 2159
rect 47 2069 81 2091
rect 47 1997 81 2023
rect 47 1925 81 1955
rect 47 1853 81 1887
rect 47 1785 81 1819
rect 47 1717 81 1747
rect 47 1649 81 1675
rect 47 1581 81 1603
rect 47 1513 81 1531
rect 47 1445 81 1459
rect 47 1377 81 1387
rect 47 1309 81 1315
rect 47 1241 81 1243
rect 47 1205 81 1207
rect 47 1133 81 1139
rect 47 1061 81 1071
rect 47 989 81 1003
rect 47 917 81 935
rect 47 845 81 867
rect 47 773 81 799
rect 47 701 81 731
rect 47 629 81 663
rect 47 561 81 595
rect 47 493 81 523
rect 47 425 81 451
rect 47 357 81 379
rect 47 289 81 307
rect 47 221 81 235
rect 47 153 81 163
rect 47 85 81 91
rect 47 17 81 19
rect 47 -19 81 -17
rect 47 -91 81 -85
rect 47 -163 81 -153
rect 47 -235 81 -221
rect 47 -307 81 -289
rect 47 -379 81 -357
rect 47 -451 81 -425
rect 47 -523 81 -493
rect 47 -595 81 -561
rect 47 -663 81 -629
rect 47 -731 81 -701
rect 47 -799 81 -773
rect 47 -867 81 -845
rect 47 -935 81 -917
rect 47 -1003 81 -989
rect 47 -1071 81 -1061
rect 47 -1139 81 -1133
rect 47 -1207 81 -1205
rect 47 -1243 81 -1241
rect 47 -1315 81 -1309
rect 47 -1387 81 -1377
rect 47 -1459 81 -1445
rect 47 -1531 81 -1513
rect 47 -1603 81 -1581
rect 47 -1675 81 -1649
rect 47 -1747 81 -1717
rect 47 -1819 81 -1785
rect 47 -1887 81 -1853
rect 47 -1955 81 -1925
rect 47 -2023 81 -1997
rect 47 -2091 81 -2069
rect 47 -2159 81 -2141
rect 47 -2227 81 -2213
rect 47 -2295 81 -2285
rect 47 -2363 81 -2357
rect 47 -2431 81 -2429
rect 47 -2467 81 -2465
rect 47 -2539 81 -2533
rect 47 -2611 81 -2601
rect 47 -2683 81 -2669
rect 47 -2755 81 -2737
rect 47 -2827 81 -2805
rect 47 -2899 81 -2873
rect 47 -2971 81 -2941
rect 47 -3043 81 -3009
rect 47 -3111 81 -3077
rect 47 -3179 81 -3149
rect 47 -3247 81 -3221
rect 47 -3315 81 -3293
rect 47 -3383 81 -3365
rect 47 -3451 81 -3437
rect 47 -3519 81 -3509
rect 47 -3587 81 -3581
rect 47 -3655 81 -3653
rect 47 -3691 81 -3689
rect 47 -3763 81 -3757
rect 47 -3835 81 -3825
rect 47 -3907 81 -3893
rect 47 -3979 81 -3961
rect 47 -4051 81 -4029
rect 47 -4123 81 -4097
rect 47 -4195 81 -4165
rect 47 -4267 81 -4233
rect 47 -4335 81 -4301
rect 47 -4403 81 -4373
rect 47 -4471 81 -4445
rect 47 -4539 81 -4517
rect 47 -4607 81 -4589
rect 47 -4675 81 -4661
rect 47 -4743 81 -4733
rect 47 -4811 81 -4805
rect 47 -4879 81 -4877
rect 47 -4915 81 -4913
rect 47 -4987 81 -4981
rect 47 -5059 81 -5049
rect 47 -5131 81 -5117
rect 47 -5203 81 -5185
rect 47 -5275 81 -5253
rect 47 -5347 81 -5321
rect 47 -5419 81 -5389
rect 47 -5491 81 -5457
rect 47 -5559 81 -5525
rect 47 -5627 81 -5597
rect 47 -5695 81 -5669
rect 47 -5763 81 -5741
rect 47 -5831 81 -5813
rect 47 -5899 81 -5885
rect 47 -5967 81 -5957
rect 47 -6035 81 -6029
rect 47 -6103 81 -6101
rect 47 -6139 81 -6137
rect 47 -6211 81 -6205
rect 47 -6283 81 -6273
rect 47 -6355 81 -6341
rect 47 -6427 81 -6409
rect 47 -6499 81 -6477
rect 47 -6571 81 -6545
rect 47 -6643 81 -6613
rect 47 -6715 81 -6681
rect 47 -6783 81 -6749
rect 47 -6851 81 -6821
rect 47 -6919 81 -6893
rect 47 -6987 81 -6965
rect 47 -7055 81 -7037
rect 47 -7123 81 -7109
rect 47 -7191 81 -7181
rect 47 -7259 81 -7253
rect 47 -7327 81 -7325
rect 47 -7363 81 -7361
rect 47 -7435 81 -7429
rect 47 -7507 81 -7497
rect 47 -7579 81 -7565
rect 47 -7651 81 -7633
rect 47 -7723 81 -7701
rect 47 -7795 81 -7769
rect 47 -7867 81 -7837
rect 47 -7939 81 -7905
rect 47 -8004 81 -7973
rect 161 7939 195 7973
rect 161 7871 195 7905
rect 161 7803 195 7837
rect 161 7735 195 7769
rect 161 7667 195 7701
rect 161 7599 195 7633
rect 161 7531 195 7565
rect 161 7463 195 7497
rect 161 7395 195 7429
rect 161 7327 195 7361
rect 161 7259 195 7293
rect 161 7191 195 7225
rect 161 7123 195 7157
rect 161 7055 195 7089
rect 161 6987 195 7021
rect 161 6919 195 6953
rect 161 6851 195 6885
rect 161 6783 195 6817
rect 161 6715 195 6749
rect 161 6647 195 6681
rect 161 6579 195 6613
rect 161 6511 195 6545
rect 161 6443 195 6477
rect 161 6375 195 6409
rect 161 6307 195 6341
rect 161 6239 195 6273
rect 161 6171 195 6205
rect 161 6103 195 6137
rect 161 6035 195 6069
rect 161 5967 195 6001
rect 161 5899 195 5933
rect 161 5831 195 5865
rect 161 5763 195 5797
rect 161 5695 195 5729
rect 161 5627 195 5661
rect 161 5559 195 5593
rect 161 5491 195 5525
rect 161 5423 195 5457
rect 161 5355 195 5389
rect 161 5287 195 5321
rect 161 5219 195 5253
rect 161 5151 195 5185
rect 161 5083 195 5117
rect 161 5015 195 5049
rect 161 4947 195 4981
rect 161 4879 195 4913
rect 161 4811 195 4845
rect 161 4743 195 4777
rect 161 4675 195 4709
rect 161 4607 195 4641
rect 161 4539 195 4573
rect 161 4471 195 4505
rect 161 4403 195 4437
rect 161 4335 195 4369
rect 161 4267 195 4301
rect 161 4199 195 4233
rect 161 4131 195 4165
rect 161 4063 195 4097
rect 161 3995 195 4029
rect 161 3927 195 3961
rect 161 3859 195 3893
rect 161 3791 195 3825
rect 161 3723 195 3757
rect 161 3655 195 3689
rect 161 3587 195 3621
rect 161 3519 195 3553
rect 161 3451 195 3485
rect 161 3383 195 3417
rect 161 3315 195 3349
rect 161 3247 195 3281
rect 161 3179 195 3213
rect 161 3111 195 3145
rect 161 3043 195 3077
rect 161 2975 195 3009
rect 161 2907 195 2941
rect 161 2839 195 2873
rect 161 2771 195 2805
rect 161 2703 195 2737
rect 161 2635 195 2669
rect 161 2567 195 2601
rect 161 2499 195 2533
rect 161 2431 195 2465
rect 161 2363 195 2397
rect 161 2295 195 2329
rect 161 2227 195 2261
rect 161 2159 195 2193
rect 161 2091 195 2125
rect 161 2023 195 2057
rect 161 1955 195 1989
rect 161 1887 195 1921
rect 161 1819 195 1853
rect 161 1751 195 1785
rect 161 1683 195 1717
rect 161 1615 195 1649
rect 161 1547 195 1581
rect 161 1479 195 1513
rect 161 1411 195 1445
rect 161 1343 195 1377
rect 161 1275 195 1309
rect 161 1207 195 1241
rect 161 1139 195 1173
rect 161 1071 195 1105
rect 161 1003 195 1037
rect 161 935 195 969
rect 161 867 195 901
rect 161 799 195 833
rect 161 731 195 765
rect 161 663 195 697
rect 161 595 195 629
rect 161 527 195 561
rect 161 459 195 493
rect 161 391 195 425
rect 161 323 195 357
rect 161 255 195 289
rect 161 187 195 221
rect 161 119 195 153
rect 161 51 195 85
rect 161 -17 195 17
rect 161 -85 195 -51
rect 161 -153 195 -119
rect 161 -221 195 -187
rect 161 -289 195 -255
rect 161 -357 195 -323
rect 161 -425 195 -391
rect 161 -493 195 -459
rect 161 -561 195 -527
rect 161 -629 195 -595
rect 161 -697 195 -663
rect 161 -765 195 -731
rect 161 -833 195 -799
rect 161 -901 195 -867
rect 161 -969 195 -935
rect 161 -1037 195 -1003
rect 161 -1105 195 -1071
rect 161 -1173 195 -1139
rect 161 -1241 195 -1207
rect 161 -1309 195 -1275
rect 161 -1377 195 -1343
rect 161 -1445 195 -1411
rect 161 -1513 195 -1479
rect 161 -1581 195 -1547
rect 161 -1649 195 -1615
rect 161 -1717 195 -1683
rect 161 -1785 195 -1751
rect 161 -1853 195 -1819
rect 161 -1921 195 -1887
rect 161 -1989 195 -1955
rect 161 -2057 195 -2023
rect 161 -2125 195 -2091
rect 161 -2193 195 -2159
rect 161 -2261 195 -2227
rect 161 -2329 195 -2295
rect 161 -2397 195 -2363
rect 161 -2465 195 -2431
rect 161 -2533 195 -2499
rect 161 -2601 195 -2567
rect 161 -2669 195 -2635
rect 161 -2737 195 -2703
rect 161 -2805 195 -2771
rect 161 -2873 195 -2839
rect 161 -2941 195 -2907
rect 161 -3009 195 -2975
rect 161 -3077 195 -3043
rect 161 -3145 195 -3111
rect 161 -3213 195 -3179
rect 161 -3281 195 -3247
rect 161 -3349 195 -3315
rect 161 -3417 195 -3383
rect 161 -3485 195 -3451
rect 161 -3553 195 -3519
rect 161 -3621 195 -3587
rect 161 -3689 195 -3655
rect 161 -3757 195 -3723
rect 161 -3825 195 -3791
rect 161 -3893 195 -3859
rect 161 -3961 195 -3927
rect 161 -4029 195 -3995
rect 161 -4097 195 -4063
rect 161 -4165 195 -4131
rect 161 -4233 195 -4199
rect 161 -4301 195 -4267
rect 161 -4369 195 -4335
rect 161 -4437 195 -4403
rect 161 -4505 195 -4471
rect 161 -4573 195 -4539
rect 161 -4641 195 -4607
rect 161 -4709 195 -4675
rect 161 -4777 195 -4743
rect 161 -4845 195 -4811
rect 161 -4913 195 -4879
rect 161 -4981 195 -4947
rect 161 -5049 195 -5015
rect 161 -5117 195 -5083
rect 161 -5185 195 -5151
rect 161 -5253 195 -5219
rect 161 -5321 195 -5287
rect 161 -5389 195 -5355
rect 161 -5457 195 -5423
rect 161 -5525 195 -5491
rect 161 -5593 195 -5559
rect 161 -5661 195 -5627
rect 161 -5729 195 -5695
rect 161 -5797 195 -5763
rect 161 -5865 195 -5831
rect 161 -5933 195 -5899
rect 161 -6001 195 -5967
rect 161 -6069 195 -6035
rect 161 -6137 195 -6103
rect 161 -6205 195 -6171
rect 161 -6273 195 -6239
rect 161 -6341 195 -6307
rect 161 -6409 195 -6375
rect 161 -6477 195 -6443
rect 161 -6545 195 -6511
rect 161 -6613 195 -6579
rect 161 -6681 195 -6647
rect 161 -6749 195 -6715
rect 161 -6817 195 -6783
rect 161 -6885 195 -6851
rect 161 -6953 195 -6919
rect 161 -7021 195 -6987
rect 161 -7089 195 -7055
rect 161 -7157 195 -7123
rect 161 -7225 195 -7191
rect 161 -7293 195 -7259
rect 161 -7361 195 -7327
rect 161 -7429 195 -7395
rect 161 -7497 195 -7463
rect 161 -7565 195 -7531
rect 161 -7633 195 -7599
rect 161 -7701 195 -7667
rect 161 -7769 195 -7735
rect 161 -7837 195 -7803
rect 161 -7905 195 -7871
rect 161 -7973 195 -7939
rect -195 -8041 -161 -8007
rect -35 -8072 -17 -8038
rect 17 -8072 35 -8038
rect 161 -8041 195 -8007
rect -195 -8140 -161 -8075
rect 161 -8140 195 -8075
rect -195 -8174 -85 -8140
rect -51 -8174 -17 -8140
rect 17 -8174 51 -8140
rect 85 -8174 195 -8140
<< viali >>
rect -17 8038 17 8072
rect -81 7939 -47 7973
rect -81 7871 -47 7901
rect -81 7867 -47 7871
rect -81 7803 -47 7829
rect -81 7795 -47 7803
rect -81 7735 -47 7757
rect -81 7723 -47 7735
rect -81 7667 -47 7685
rect -81 7651 -47 7667
rect -81 7599 -47 7613
rect -81 7579 -47 7599
rect -81 7531 -47 7541
rect -81 7507 -47 7531
rect -81 7463 -47 7469
rect -81 7435 -47 7463
rect -81 7395 -47 7397
rect -81 7363 -47 7395
rect -81 7293 -47 7325
rect -81 7291 -47 7293
rect -81 7225 -47 7253
rect -81 7219 -47 7225
rect -81 7157 -47 7181
rect -81 7147 -47 7157
rect -81 7089 -47 7109
rect -81 7075 -47 7089
rect -81 7021 -47 7037
rect -81 7003 -47 7021
rect -81 6953 -47 6965
rect -81 6931 -47 6953
rect -81 6885 -47 6893
rect -81 6859 -47 6885
rect -81 6817 -47 6821
rect -81 6787 -47 6817
rect -81 6715 -47 6749
rect -81 6647 -47 6677
rect -81 6643 -47 6647
rect -81 6579 -47 6605
rect -81 6571 -47 6579
rect -81 6511 -47 6533
rect -81 6499 -47 6511
rect -81 6443 -47 6461
rect -81 6427 -47 6443
rect -81 6375 -47 6389
rect -81 6355 -47 6375
rect -81 6307 -47 6317
rect -81 6283 -47 6307
rect -81 6239 -47 6245
rect -81 6211 -47 6239
rect -81 6171 -47 6173
rect -81 6139 -47 6171
rect -81 6069 -47 6101
rect -81 6067 -47 6069
rect -81 6001 -47 6029
rect -81 5995 -47 6001
rect -81 5933 -47 5957
rect -81 5923 -47 5933
rect -81 5865 -47 5885
rect -81 5851 -47 5865
rect -81 5797 -47 5813
rect -81 5779 -47 5797
rect -81 5729 -47 5741
rect -81 5707 -47 5729
rect -81 5661 -47 5669
rect -81 5635 -47 5661
rect -81 5593 -47 5597
rect -81 5563 -47 5593
rect -81 5491 -47 5525
rect -81 5423 -47 5453
rect -81 5419 -47 5423
rect -81 5355 -47 5381
rect -81 5347 -47 5355
rect -81 5287 -47 5309
rect -81 5275 -47 5287
rect -81 5219 -47 5237
rect -81 5203 -47 5219
rect -81 5151 -47 5165
rect -81 5131 -47 5151
rect -81 5083 -47 5093
rect -81 5059 -47 5083
rect -81 5015 -47 5021
rect -81 4987 -47 5015
rect -81 4947 -47 4949
rect -81 4915 -47 4947
rect -81 4845 -47 4877
rect -81 4843 -47 4845
rect -81 4777 -47 4805
rect -81 4771 -47 4777
rect -81 4709 -47 4733
rect -81 4699 -47 4709
rect -81 4641 -47 4661
rect -81 4627 -47 4641
rect -81 4573 -47 4589
rect -81 4555 -47 4573
rect -81 4505 -47 4517
rect -81 4483 -47 4505
rect -81 4437 -47 4445
rect -81 4411 -47 4437
rect -81 4369 -47 4373
rect -81 4339 -47 4369
rect -81 4267 -47 4301
rect -81 4199 -47 4229
rect -81 4195 -47 4199
rect -81 4131 -47 4157
rect -81 4123 -47 4131
rect -81 4063 -47 4085
rect -81 4051 -47 4063
rect -81 3995 -47 4013
rect -81 3979 -47 3995
rect -81 3927 -47 3941
rect -81 3907 -47 3927
rect -81 3859 -47 3869
rect -81 3835 -47 3859
rect -81 3791 -47 3797
rect -81 3763 -47 3791
rect -81 3723 -47 3725
rect -81 3691 -47 3723
rect -81 3621 -47 3653
rect -81 3619 -47 3621
rect -81 3553 -47 3581
rect -81 3547 -47 3553
rect -81 3485 -47 3509
rect -81 3475 -47 3485
rect -81 3417 -47 3437
rect -81 3403 -47 3417
rect -81 3349 -47 3365
rect -81 3331 -47 3349
rect -81 3281 -47 3293
rect -81 3259 -47 3281
rect -81 3213 -47 3221
rect -81 3187 -47 3213
rect -81 3145 -47 3149
rect -81 3115 -47 3145
rect -81 3043 -47 3077
rect -81 2975 -47 3005
rect -81 2971 -47 2975
rect -81 2907 -47 2933
rect -81 2899 -47 2907
rect -81 2839 -47 2861
rect -81 2827 -47 2839
rect -81 2771 -47 2789
rect -81 2755 -47 2771
rect -81 2703 -47 2717
rect -81 2683 -47 2703
rect -81 2635 -47 2645
rect -81 2611 -47 2635
rect -81 2567 -47 2573
rect -81 2539 -47 2567
rect -81 2499 -47 2501
rect -81 2467 -47 2499
rect -81 2397 -47 2429
rect -81 2395 -47 2397
rect -81 2329 -47 2357
rect -81 2323 -47 2329
rect -81 2261 -47 2285
rect -81 2251 -47 2261
rect -81 2193 -47 2213
rect -81 2179 -47 2193
rect -81 2125 -47 2141
rect -81 2107 -47 2125
rect -81 2057 -47 2069
rect -81 2035 -47 2057
rect -81 1989 -47 1997
rect -81 1963 -47 1989
rect -81 1921 -47 1925
rect -81 1891 -47 1921
rect -81 1819 -47 1853
rect -81 1751 -47 1781
rect -81 1747 -47 1751
rect -81 1683 -47 1709
rect -81 1675 -47 1683
rect -81 1615 -47 1637
rect -81 1603 -47 1615
rect -81 1547 -47 1565
rect -81 1531 -47 1547
rect -81 1479 -47 1493
rect -81 1459 -47 1479
rect -81 1411 -47 1421
rect -81 1387 -47 1411
rect -81 1343 -47 1349
rect -81 1315 -47 1343
rect -81 1275 -47 1277
rect -81 1243 -47 1275
rect -81 1173 -47 1205
rect -81 1171 -47 1173
rect -81 1105 -47 1133
rect -81 1099 -47 1105
rect -81 1037 -47 1061
rect -81 1027 -47 1037
rect -81 969 -47 989
rect -81 955 -47 969
rect -81 901 -47 917
rect -81 883 -47 901
rect -81 833 -47 845
rect -81 811 -47 833
rect -81 765 -47 773
rect -81 739 -47 765
rect -81 697 -47 701
rect -81 667 -47 697
rect -81 595 -47 629
rect -81 527 -47 557
rect -81 523 -47 527
rect -81 459 -47 485
rect -81 451 -47 459
rect -81 391 -47 413
rect -81 379 -47 391
rect -81 323 -47 341
rect -81 307 -47 323
rect -81 255 -47 269
rect -81 235 -47 255
rect -81 187 -47 197
rect -81 163 -47 187
rect -81 119 -47 125
rect -81 91 -47 119
rect -81 51 -47 53
rect -81 19 -47 51
rect -81 -51 -47 -19
rect -81 -53 -47 -51
rect -81 -119 -47 -91
rect -81 -125 -47 -119
rect -81 -187 -47 -163
rect -81 -197 -47 -187
rect -81 -255 -47 -235
rect -81 -269 -47 -255
rect -81 -323 -47 -307
rect -81 -341 -47 -323
rect -81 -391 -47 -379
rect -81 -413 -47 -391
rect -81 -459 -47 -451
rect -81 -485 -47 -459
rect -81 -527 -47 -523
rect -81 -557 -47 -527
rect -81 -629 -47 -595
rect -81 -697 -47 -667
rect -81 -701 -47 -697
rect -81 -765 -47 -739
rect -81 -773 -47 -765
rect -81 -833 -47 -811
rect -81 -845 -47 -833
rect -81 -901 -47 -883
rect -81 -917 -47 -901
rect -81 -969 -47 -955
rect -81 -989 -47 -969
rect -81 -1037 -47 -1027
rect -81 -1061 -47 -1037
rect -81 -1105 -47 -1099
rect -81 -1133 -47 -1105
rect -81 -1173 -47 -1171
rect -81 -1205 -47 -1173
rect -81 -1275 -47 -1243
rect -81 -1277 -47 -1275
rect -81 -1343 -47 -1315
rect -81 -1349 -47 -1343
rect -81 -1411 -47 -1387
rect -81 -1421 -47 -1411
rect -81 -1479 -47 -1459
rect -81 -1493 -47 -1479
rect -81 -1547 -47 -1531
rect -81 -1565 -47 -1547
rect -81 -1615 -47 -1603
rect -81 -1637 -47 -1615
rect -81 -1683 -47 -1675
rect -81 -1709 -47 -1683
rect -81 -1751 -47 -1747
rect -81 -1781 -47 -1751
rect -81 -1853 -47 -1819
rect -81 -1921 -47 -1891
rect -81 -1925 -47 -1921
rect -81 -1989 -47 -1963
rect -81 -1997 -47 -1989
rect -81 -2057 -47 -2035
rect -81 -2069 -47 -2057
rect -81 -2125 -47 -2107
rect -81 -2141 -47 -2125
rect -81 -2193 -47 -2179
rect -81 -2213 -47 -2193
rect -81 -2261 -47 -2251
rect -81 -2285 -47 -2261
rect -81 -2329 -47 -2323
rect -81 -2357 -47 -2329
rect -81 -2397 -47 -2395
rect -81 -2429 -47 -2397
rect -81 -2499 -47 -2467
rect -81 -2501 -47 -2499
rect -81 -2567 -47 -2539
rect -81 -2573 -47 -2567
rect -81 -2635 -47 -2611
rect -81 -2645 -47 -2635
rect -81 -2703 -47 -2683
rect -81 -2717 -47 -2703
rect -81 -2771 -47 -2755
rect -81 -2789 -47 -2771
rect -81 -2839 -47 -2827
rect -81 -2861 -47 -2839
rect -81 -2907 -47 -2899
rect -81 -2933 -47 -2907
rect -81 -2975 -47 -2971
rect -81 -3005 -47 -2975
rect -81 -3077 -47 -3043
rect -81 -3145 -47 -3115
rect -81 -3149 -47 -3145
rect -81 -3213 -47 -3187
rect -81 -3221 -47 -3213
rect -81 -3281 -47 -3259
rect -81 -3293 -47 -3281
rect -81 -3349 -47 -3331
rect -81 -3365 -47 -3349
rect -81 -3417 -47 -3403
rect -81 -3437 -47 -3417
rect -81 -3485 -47 -3475
rect -81 -3509 -47 -3485
rect -81 -3553 -47 -3547
rect -81 -3581 -47 -3553
rect -81 -3621 -47 -3619
rect -81 -3653 -47 -3621
rect -81 -3723 -47 -3691
rect -81 -3725 -47 -3723
rect -81 -3791 -47 -3763
rect -81 -3797 -47 -3791
rect -81 -3859 -47 -3835
rect -81 -3869 -47 -3859
rect -81 -3927 -47 -3907
rect -81 -3941 -47 -3927
rect -81 -3995 -47 -3979
rect -81 -4013 -47 -3995
rect -81 -4063 -47 -4051
rect -81 -4085 -47 -4063
rect -81 -4131 -47 -4123
rect -81 -4157 -47 -4131
rect -81 -4199 -47 -4195
rect -81 -4229 -47 -4199
rect -81 -4301 -47 -4267
rect -81 -4369 -47 -4339
rect -81 -4373 -47 -4369
rect -81 -4437 -47 -4411
rect -81 -4445 -47 -4437
rect -81 -4505 -47 -4483
rect -81 -4517 -47 -4505
rect -81 -4573 -47 -4555
rect -81 -4589 -47 -4573
rect -81 -4641 -47 -4627
rect -81 -4661 -47 -4641
rect -81 -4709 -47 -4699
rect -81 -4733 -47 -4709
rect -81 -4777 -47 -4771
rect -81 -4805 -47 -4777
rect -81 -4845 -47 -4843
rect -81 -4877 -47 -4845
rect -81 -4947 -47 -4915
rect -81 -4949 -47 -4947
rect -81 -5015 -47 -4987
rect -81 -5021 -47 -5015
rect -81 -5083 -47 -5059
rect -81 -5093 -47 -5083
rect -81 -5151 -47 -5131
rect -81 -5165 -47 -5151
rect -81 -5219 -47 -5203
rect -81 -5237 -47 -5219
rect -81 -5287 -47 -5275
rect -81 -5309 -47 -5287
rect -81 -5355 -47 -5347
rect -81 -5381 -47 -5355
rect -81 -5423 -47 -5419
rect -81 -5453 -47 -5423
rect -81 -5525 -47 -5491
rect -81 -5593 -47 -5563
rect -81 -5597 -47 -5593
rect -81 -5661 -47 -5635
rect -81 -5669 -47 -5661
rect -81 -5729 -47 -5707
rect -81 -5741 -47 -5729
rect -81 -5797 -47 -5779
rect -81 -5813 -47 -5797
rect -81 -5865 -47 -5851
rect -81 -5885 -47 -5865
rect -81 -5933 -47 -5923
rect -81 -5957 -47 -5933
rect -81 -6001 -47 -5995
rect -81 -6029 -47 -6001
rect -81 -6069 -47 -6067
rect -81 -6101 -47 -6069
rect -81 -6171 -47 -6139
rect -81 -6173 -47 -6171
rect -81 -6239 -47 -6211
rect -81 -6245 -47 -6239
rect -81 -6307 -47 -6283
rect -81 -6317 -47 -6307
rect -81 -6375 -47 -6355
rect -81 -6389 -47 -6375
rect -81 -6443 -47 -6427
rect -81 -6461 -47 -6443
rect -81 -6511 -47 -6499
rect -81 -6533 -47 -6511
rect -81 -6579 -47 -6571
rect -81 -6605 -47 -6579
rect -81 -6647 -47 -6643
rect -81 -6677 -47 -6647
rect -81 -6749 -47 -6715
rect -81 -6817 -47 -6787
rect -81 -6821 -47 -6817
rect -81 -6885 -47 -6859
rect -81 -6893 -47 -6885
rect -81 -6953 -47 -6931
rect -81 -6965 -47 -6953
rect -81 -7021 -47 -7003
rect -81 -7037 -47 -7021
rect -81 -7089 -47 -7075
rect -81 -7109 -47 -7089
rect -81 -7157 -47 -7147
rect -81 -7181 -47 -7157
rect -81 -7225 -47 -7219
rect -81 -7253 -47 -7225
rect -81 -7293 -47 -7291
rect -81 -7325 -47 -7293
rect -81 -7395 -47 -7363
rect -81 -7397 -47 -7395
rect -81 -7463 -47 -7435
rect -81 -7469 -47 -7463
rect -81 -7531 -47 -7507
rect -81 -7541 -47 -7531
rect -81 -7599 -47 -7579
rect -81 -7613 -47 -7599
rect -81 -7667 -47 -7651
rect -81 -7685 -47 -7667
rect -81 -7735 -47 -7723
rect -81 -7757 -47 -7735
rect -81 -7803 -47 -7795
rect -81 -7829 -47 -7803
rect -81 -7871 -47 -7867
rect -81 -7901 -47 -7871
rect -81 -7973 -47 -7939
rect 47 7939 81 7973
rect 47 7871 81 7901
rect 47 7867 81 7871
rect 47 7803 81 7829
rect 47 7795 81 7803
rect 47 7735 81 7757
rect 47 7723 81 7735
rect 47 7667 81 7685
rect 47 7651 81 7667
rect 47 7599 81 7613
rect 47 7579 81 7599
rect 47 7531 81 7541
rect 47 7507 81 7531
rect 47 7463 81 7469
rect 47 7435 81 7463
rect 47 7395 81 7397
rect 47 7363 81 7395
rect 47 7293 81 7325
rect 47 7291 81 7293
rect 47 7225 81 7253
rect 47 7219 81 7225
rect 47 7157 81 7181
rect 47 7147 81 7157
rect 47 7089 81 7109
rect 47 7075 81 7089
rect 47 7021 81 7037
rect 47 7003 81 7021
rect 47 6953 81 6965
rect 47 6931 81 6953
rect 47 6885 81 6893
rect 47 6859 81 6885
rect 47 6817 81 6821
rect 47 6787 81 6817
rect 47 6715 81 6749
rect 47 6647 81 6677
rect 47 6643 81 6647
rect 47 6579 81 6605
rect 47 6571 81 6579
rect 47 6511 81 6533
rect 47 6499 81 6511
rect 47 6443 81 6461
rect 47 6427 81 6443
rect 47 6375 81 6389
rect 47 6355 81 6375
rect 47 6307 81 6317
rect 47 6283 81 6307
rect 47 6239 81 6245
rect 47 6211 81 6239
rect 47 6171 81 6173
rect 47 6139 81 6171
rect 47 6069 81 6101
rect 47 6067 81 6069
rect 47 6001 81 6029
rect 47 5995 81 6001
rect 47 5933 81 5957
rect 47 5923 81 5933
rect 47 5865 81 5885
rect 47 5851 81 5865
rect 47 5797 81 5813
rect 47 5779 81 5797
rect 47 5729 81 5741
rect 47 5707 81 5729
rect 47 5661 81 5669
rect 47 5635 81 5661
rect 47 5593 81 5597
rect 47 5563 81 5593
rect 47 5491 81 5525
rect 47 5423 81 5453
rect 47 5419 81 5423
rect 47 5355 81 5381
rect 47 5347 81 5355
rect 47 5287 81 5309
rect 47 5275 81 5287
rect 47 5219 81 5237
rect 47 5203 81 5219
rect 47 5151 81 5165
rect 47 5131 81 5151
rect 47 5083 81 5093
rect 47 5059 81 5083
rect 47 5015 81 5021
rect 47 4987 81 5015
rect 47 4947 81 4949
rect 47 4915 81 4947
rect 47 4845 81 4877
rect 47 4843 81 4845
rect 47 4777 81 4805
rect 47 4771 81 4777
rect 47 4709 81 4733
rect 47 4699 81 4709
rect 47 4641 81 4661
rect 47 4627 81 4641
rect 47 4573 81 4589
rect 47 4555 81 4573
rect 47 4505 81 4517
rect 47 4483 81 4505
rect 47 4437 81 4445
rect 47 4411 81 4437
rect 47 4369 81 4373
rect 47 4339 81 4369
rect 47 4267 81 4301
rect 47 4199 81 4229
rect 47 4195 81 4199
rect 47 4131 81 4157
rect 47 4123 81 4131
rect 47 4063 81 4085
rect 47 4051 81 4063
rect 47 3995 81 4013
rect 47 3979 81 3995
rect 47 3927 81 3941
rect 47 3907 81 3927
rect 47 3859 81 3869
rect 47 3835 81 3859
rect 47 3791 81 3797
rect 47 3763 81 3791
rect 47 3723 81 3725
rect 47 3691 81 3723
rect 47 3621 81 3653
rect 47 3619 81 3621
rect 47 3553 81 3581
rect 47 3547 81 3553
rect 47 3485 81 3509
rect 47 3475 81 3485
rect 47 3417 81 3437
rect 47 3403 81 3417
rect 47 3349 81 3365
rect 47 3331 81 3349
rect 47 3281 81 3293
rect 47 3259 81 3281
rect 47 3213 81 3221
rect 47 3187 81 3213
rect 47 3145 81 3149
rect 47 3115 81 3145
rect 47 3043 81 3077
rect 47 2975 81 3005
rect 47 2971 81 2975
rect 47 2907 81 2933
rect 47 2899 81 2907
rect 47 2839 81 2861
rect 47 2827 81 2839
rect 47 2771 81 2789
rect 47 2755 81 2771
rect 47 2703 81 2717
rect 47 2683 81 2703
rect 47 2635 81 2645
rect 47 2611 81 2635
rect 47 2567 81 2573
rect 47 2539 81 2567
rect 47 2499 81 2501
rect 47 2467 81 2499
rect 47 2397 81 2429
rect 47 2395 81 2397
rect 47 2329 81 2357
rect 47 2323 81 2329
rect 47 2261 81 2285
rect 47 2251 81 2261
rect 47 2193 81 2213
rect 47 2179 81 2193
rect 47 2125 81 2141
rect 47 2107 81 2125
rect 47 2057 81 2069
rect 47 2035 81 2057
rect 47 1989 81 1997
rect 47 1963 81 1989
rect 47 1921 81 1925
rect 47 1891 81 1921
rect 47 1819 81 1853
rect 47 1751 81 1781
rect 47 1747 81 1751
rect 47 1683 81 1709
rect 47 1675 81 1683
rect 47 1615 81 1637
rect 47 1603 81 1615
rect 47 1547 81 1565
rect 47 1531 81 1547
rect 47 1479 81 1493
rect 47 1459 81 1479
rect 47 1411 81 1421
rect 47 1387 81 1411
rect 47 1343 81 1349
rect 47 1315 81 1343
rect 47 1275 81 1277
rect 47 1243 81 1275
rect 47 1173 81 1205
rect 47 1171 81 1173
rect 47 1105 81 1133
rect 47 1099 81 1105
rect 47 1037 81 1061
rect 47 1027 81 1037
rect 47 969 81 989
rect 47 955 81 969
rect 47 901 81 917
rect 47 883 81 901
rect 47 833 81 845
rect 47 811 81 833
rect 47 765 81 773
rect 47 739 81 765
rect 47 697 81 701
rect 47 667 81 697
rect 47 595 81 629
rect 47 527 81 557
rect 47 523 81 527
rect 47 459 81 485
rect 47 451 81 459
rect 47 391 81 413
rect 47 379 81 391
rect 47 323 81 341
rect 47 307 81 323
rect 47 255 81 269
rect 47 235 81 255
rect 47 187 81 197
rect 47 163 81 187
rect 47 119 81 125
rect 47 91 81 119
rect 47 51 81 53
rect 47 19 81 51
rect 47 -51 81 -19
rect 47 -53 81 -51
rect 47 -119 81 -91
rect 47 -125 81 -119
rect 47 -187 81 -163
rect 47 -197 81 -187
rect 47 -255 81 -235
rect 47 -269 81 -255
rect 47 -323 81 -307
rect 47 -341 81 -323
rect 47 -391 81 -379
rect 47 -413 81 -391
rect 47 -459 81 -451
rect 47 -485 81 -459
rect 47 -527 81 -523
rect 47 -557 81 -527
rect 47 -629 81 -595
rect 47 -697 81 -667
rect 47 -701 81 -697
rect 47 -765 81 -739
rect 47 -773 81 -765
rect 47 -833 81 -811
rect 47 -845 81 -833
rect 47 -901 81 -883
rect 47 -917 81 -901
rect 47 -969 81 -955
rect 47 -989 81 -969
rect 47 -1037 81 -1027
rect 47 -1061 81 -1037
rect 47 -1105 81 -1099
rect 47 -1133 81 -1105
rect 47 -1173 81 -1171
rect 47 -1205 81 -1173
rect 47 -1275 81 -1243
rect 47 -1277 81 -1275
rect 47 -1343 81 -1315
rect 47 -1349 81 -1343
rect 47 -1411 81 -1387
rect 47 -1421 81 -1411
rect 47 -1479 81 -1459
rect 47 -1493 81 -1479
rect 47 -1547 81 -1531
rect 47 -1565 81 -1547
rect 47 -1615 81 -1603
rect 47 -1637 81 -1615
rect 47 -1683 81 -1675
rect 47 -1709 81 -1683
rect 47 -1751 81 -1747
rect 47 -1781 81 -1751
rect 47 -1853 81 -1819
rect 47 -1921 81 -1891
rect 47 -1925 81 -1921
rect 47 -1989 81 -1963
rect 47 -1997 81 -1989
rect 47 -2057 81 -2035
rect 47 -2069 81 -2057
rect 47 -2125 81 -2107
rect 47 -2141 81 -2125
rect 47 -2193 81 -2179
rect 47 -2213 81 -2193
rect 47 -2261 81 -2251
rect 47 -2285 81 -2261
rect 47 -2329 81 -2323
rect 47 -2357 81 -2329
rect 47 -2397 81 -2395
rect 47 -2429 81 -2397
rect 47 -2499 81 -2467
rect 47 -2501 81 -2499
rect 47 -2567 81 -2539
rect 47 -2573 81 -2567
rect 47 -2635 81 -2611
rect 47 -2645 81 -2635
rect 47 -2703 81 -2683
rect 47 -2717 81 -2703
rect 47 -2771 81 -2755
rect 47 -2789 81 -2771
rect 47 -2839 81 -2827
rect 47 -2861 81 -2839
rect 47 -2907 81 -2899
rect 47 -2933 81 -2907
rect 47 -2975 81 -2971
rect 47 -3005 81 -2975
rect 47 -3077 81 -3043
rect 47 -3145 81 -3115
rect 47 -3149 81 -3145
rect 47 -3213 81 -3187
rect 47 -3221 81 -3213
rect 47 -3281 81 -3259
rect 47 -3293 81 -3281
rect 47 -3349 81 -3331
rect 47 -3365 81 -3349
rect 47 -3417 81 -3403
rect 47 -3437 81 -3417
rect 47 -3485 81 -3475
rect 47 -3509 81 -3485
rect 47 -3553 81 -3547
rect 47 -3581 81 -3553
rect 47 -3621 81 -3619
rect 47 -3653 81 -3621
rect 47 -3723 81 -3691
rect 47 -3725 81 -3723
rect 47 -3791 81 -3763
rect 47 -3797 81 -3791
rect 47 -3859 81 -3835
rect 47 -3869 81 -3859
rect 47 -3927 81 -3907
rect 47 -3941 81 -3927
rect 47 -3995 81 -3979
rect 47 -4013 81 -3995
rect 47 -4063 81 -4051
rect 47 -4085 81 -4063
rect 47 -4131 81 -4123
rect 47 -4157 81 -4131
rect 47 -4199 81 -4195
rect 47 -4229 81 -4199
rect 47 -4301 81 -4267
rect 47 -4369 81 -4339
rect 47 -4373 81 -4369
rect 47 -4437 81 -4411
rect 47 -4445 81 -4437
rect 47 -4505 81 -4483
rect 47 -4517 81 -4505
rect 47 -4573 81 -4555
rect 47 -4589 81 -4573
rect 47 -4641 81 -4627
rect 47 -4661 81 -4641
rect 47 -4709 81 -4699
rect 47 -4733 81 -4709
rect 47 -4777 81 -4771
rect 47 -4805 81 -4777
rect 47 -4845 81 -4843
rect 47 -4877 81 -4845
rect 47 -4947 81 -4915
rect 47 -4949 81 -4947
rect 47 -5015 81 -4987
rect 47 -5021 81 -5015
rect 47 -5083 81 -5059
rect 47 -5093 81 -5083
rect 47 -5151 81 -5131
rect 47 -5165 81 -5151
rect 47 -5219 81 -5203
rect 47 -5237 81 -5219
rect 47 -5287 81 -5275
rect 47 -5309 81 -5287
rect 47 -5355 81 -5347
rect 47 -5381 81 -5355
rect 47 -5423 81 -5419
rect 47 -5453 81 -5423
rect 47 -5525 81 -5491
rect 47 -5593 81 -5563
rect 47 -5597 81 -5593
rect 47 -5661 81 -5635
rect 47 -5669 81 -5661
rect 47 -5729 81 -5707
rect 47 -5741 81 -5729
rect 47 -5797 81 -5779
rect 47 -5813 81 -5797
rect 47 -5865 81 -5851
rect 47 -5885 81 -5865
rect 47 -5933 81 -5923
rect 47 -5957 81 -5933
rect 47 -6001 81 -5995
rect 47 -6029 81 -6001
rect 47 -6069 81 -6067
rect 47 -6101 81 -6069
rect 47 -6171 81 -6139
rect 47 -6173 81 -6171
rect 47 -6239 81 -6211
rect 47 -6245 81 -6239
rect 47 -6307 81 -6283
rect 47 -6317 81 -6307
rect 47 -6375 81 -6355
rect 47 -6389 81 -6375
rect 47 -6443 81 -6427
rect 47 -6461 81 -6443
rect 47 -6511 81 -6499
rect 47 -6533 81 -6511
rect 47 -6579 81 -6571
rect 47 -6605 81 -6579
rect 47 -6647 81 -6643
rect 47 -6677 81 -6647
rect 47 -6749 81 -6715
rect 47 -6817 81 -6787
rect 47 -6821 81 -6817
rect 47 -6885 81 -6859
rect 47 -6893 81 -6885
rect 47 -6953 81 -6931
rect 47 -6965 81 -6953
rect 47 -7021 81 -7003
rect 47 -7037 81 -7021
rect 47 -7089 81 -7075
rect 47 -7109 81 -7089
rect 47 -7157 81 -7147
rect 47 -7181 81 -7157
rect 47 -7225 81 -7219
rect 47 -7253 81 -7225
rect 47 -7293 81 -7291
rect 47 -7325 81 -7293
rect 47 -7395 81 -7363
rect 47 -7397 81 -7395
rect 47 -7463 81 -7435
rect 47 -7469 81 -7463
rect 47 -7531 81 -7507
rect 47 -7541 81 -7531
rect 47 -7599 81 -7579
rect 47 -7613 81 -7599
rect 47 -7667 81 -7651
rect 47 -7685 81 -7667
rect 47 -7735 81 -7723
rect 47 -7757 81 -7735
rect 47 -7803 81 -7795
rect 47 -7829 81 -7803
rect 47 -7871 81 -7867
rect 47 -7901 81 -7871
rect 47 -7973 81 -7939
rect -17 -8072 17 -8038
<< metal1 >>
rect -31 8072 31 8078
rect -31 8038 -17 8072
rect 17 8038 31 8072
rect -31 8032 31 8038
rect -87 7973 -41 8000
rect -87 7939 -81 7973
rect -47 7939 -41 7973
rect -87 7901 -41 7939
rect -87 7867 -81 7901
rect -47 7867 -41 7901
rect -87 7829 -41 7867
rect -87 7795 -81 7829
rect -47 7795 -41 7829
rect -87 7757 -41 7795
rect -87 7723 -81 7757
rect -47 7723 -41 7757
rect -87 7685 -41 7723
rect -87 7651 -81 7685
rect -47 7651 -41 7685
rect -87 7613 -41 7651
rect -87 7579 -81 7613
rect -47 7579 -41 7613
rect -87 7541 -41 7579
rect -87 7507 -81 7541
rect -47 7507 -41 7541
rect -87 7469 -41 7507
rect -87 7435 -81 7469
rect -47 7435 -41 7469
rect -87 7397 -41 7435
rect -87 7363 -81 7397
rect -47 7363 -41 7397
rect -87 7325 -41 7363
rect -87 7291 -81 7325
rect -47 7291 -41 7325
rect -87 7253 -41 7291
rect -87 7219 -81 7253
rect -47 7219 -41 7253
rect -87 7181 -41 7219
rect -87 7147 -81 7181
rect -47 7147 -41 7181
rect -87 7109 -41 7147
rect -87 7075 -81 7109
rect -47 7075 -41 7109
rect -87 7037 -41 7075
rect -87 7003 -81 7037
rect -47 7003 -41 7037
rect -87 6965 -41 7003
rect -87 6931 -81 6965
rect -47 6931 -41 6965
rect -87 6893 -41 6931
rect -87 6859 -81 6893
rect -47 6859 -41 6893
rect -87 6821 -41 6859
rect -87 6787 -81 6821
rect -47 6787 -41 6821
rect -87 6749 -41 6787
rect -87 6715 -81 6749
rect -47 6715 -41 6749
rect -87 6677 -41 6715
rect -87 6643 -81 6677
rect -47 6643 -41 6677
rect -87 6605 -41 6643
rect -87 6571 -81 6605
rect -47 6571 -41 6605
rect -87 6533 -41 6571
rect -87 6499 -81 6533
rect -47 6499 -41 6533
rect -87 6461 -41 6499
rect -87 6427 -81 6461
rect -47 6427 -41 6461
rect -87 6389 -41 6427
rect -87 6355 -81 6389
rect -47 6355 -41 6389
rect -87 6317 -41 6355
rect -87 6283 -81 6317
rect -47 6283 -41 6317
rect -87 6245 -41 6283
rect -87 6211 -81 6245
rect -47 6211 -41 6245
rect -87 6173 -41 6211
rect -87 6139 -81 6173
rect -47 6139 -41 6173
rect -87 6101 -41 6139
rect -87 6067 -81 6101
rect -47 6067 -41 6101
rect -87 6029 -41 6067
rect -87 5995 -81 6029
rect -47 5995 -41 6029
rect -87 5957 -41 5995
rect -87 5923 -81 5957
rect -47 5923 -41 5957
rect -87 5885 -41 5923
rect -87 5851 -81 5885
rect -47 5851 -41 5885
rect -87 5813 -41 5851
rect -87 5779 -81 5813
rect -47 5779 -41 5813
rect -87 5741 -41 5779
rect -87 5707 -81 5741
rect -47 5707 -41 5741
rect -87 5669 -41 5707
rect -87 5635 -81 5669
rect -47 5635 -41 5669
rect -87 5597 -41 5635
rect -87 5563 -81 5597
rect -47 5563 -41 5597
rect -87 5525 -41 5563
rect -87 5491 -81 5525
rect -47 5491 -41 5525
rect -87 5453 -41 5491
rect -87 5419 -81 5453
rect -47 5419 -41 5453
rect -87 5381 -41 5419
rect -87 5347 -81 5381
rect -47 5347 -41 5381
rect -87 5309 -41 5347
rect -87 5275 -81 5309
rect -47 5275 -41 5309
rect -87 5237 -41 5275
rect -87 5203 -81 5237
rect -47 5203 -41 5237
rect -87 5165 -41 5203
rect -87 5131 -81 5165
rect -47 5131 -41 5165
rect -87 5093 -41 5131
rect -87 5059 -81 5093
rect -47 5059 -41 5093
rect -87 5021 -41 5059
rect -87 4987 -81 5021
rect -47 4987 -41 5021
rect -87 4949 -41 4987
rect -87 4915 -81 4949
rect -47 4915 -41 4949
rect -87 4877 -41 4915
rect -87 4843 -81 4877
rect -47 4843 -41 4877
rect -87 4805 -41 4843
rect -87 4771 -81 4805
rect -47 4771 -41 4805
rect -87 4733 -41 4771
rect -87 4699 -81 4733
rect -47 4699 -41 4733
rect -87 4661 -41 4699
rect -87 4627 -81 4661
rect -47 4627 -41 4661
rect -87 4589 -41 4627
rect -87 4555 -81 4589
rect -47 4555 -41 4589
rect -87 4517 -41 4555
rect -87 4483 -81 4517
rect -47 4483 -41 4517
rect -87 4445 -41 4483
rect -87 4411 -81 4445
rect -47 4411 -41 4445
rect -87 4373 -41 4411
rect -87 4339 -81 4373
rect -47 4339 -41 4373
rect -87 4301 -41 4339
rect -87 4267 -81 4301
rect -47 4267 -41 4301
rect -87 4229 -41 4267
rect -87 4195 -81 4229
rect -47 4195 -41 4229
rect -87 4157 -41 4195
rect -87 4123 -81 4157
rect -47 4123 -41 4157
rect -87 4085 -41 4123
rect -87 4051 -81 4085
rect -47 4051 -41 4085
rect -87 4013 -41 4051
rect -87 3979 -81 4013
rect -47 3979 -41 4013
rect -87 3941 -41 3979
rect -87 3907 -81 3941
rect -47 3907 -41 3941
rect -87 3869 -41 3907
rect -87 3835 -81 3869
rect -47 3835 -41 3869
rect -87 3797 -41 3835
rect -87 3763 -81 3797
rect -47 3763 -41 3797
rect -87 3725 -41 3763
rect -87 3691 -81 3725
rect -47 3691 -41 3725
rect -87 3653 -41 3691
rect -87 3619 -81 3653
rect -47 3619 -41 3653
rect -87 3581 -41 3619
rect -87 3547 -81 3581
rect -47 3547 -41 3581
rect -87 3509 -41 3547
rect -87 3475 -81 3509
rect -47 3475 -41 3509
rect -87 3437 -41 3475
rect -87 3403 -81 3437
rect -47 3403 -41 3437
rect -87 3365 -41 3403
rect -87 3331 -81 3365
rect -47 3331 -41 3365
rect -87 3293 -41 3331
rect -87 3259 -81 3293
rect -47 3259 -41 3293
rect -87 3221 -41 3259
rect -87 3187 -81 3221
rect -47 3187 -41 3221
rect -87 3149 -41 3187
rect -87 3115 -81 3149
rect -47 3115 -41 3149
rect -87 3077 -41 3115
rect -87 3043 -81 3077
rect -47 3043 -41 3077
rect -87 3005 -41 3043
rect -87 2971 -81 3005
rect -47 2971 -41 3005
rect -87 2933 -41 2971
rect -87 2899 -81 2933
rect -47 2899 -41 2933
rect -87 2861 -41 2899
rect -87 2827 -81 2861
rect -47 2827 -41 2861
rect -87 2789 -41 2827
rect -87 2755 -81 2789
rect -47 2755 -41 2789
rect -87 2717 -41 2755
rect -87 2683 -81 2717
rect -47 2683 -41 2717
rect -87 2645 -41 2683
rect -87 2611 -81 2645
rect -47 2611 -41 2645
rect -87 2573 -41 2611
rect -87 2539 -81 2573
rect -47 2539 -41 2573
rect -87 2501 -41 2539
rect -87 2467 -81 2501
rect -47 2467 -41 2501
rect -87 2429 -41 2467
rect -87 2395 -81 2429
rect -47 2395 -41 2429
rect -87 2357 -41 2395
rect -87 2323 -81 2357
rect -47 2323 -41 2357
rect -87 2285 -41 2323
rect -87 2251 -81 2285
rect -47 2251 -41 2285
rect -87 2213 -41 2251
rect -87 2179 -81 2213
rect -47 2179 -41 2213
rect -87 2141 -41 2179
rect -87 2107 -81 2141
rect -47 2107 -41 2141
rect -87 2069 -41 2107
rect -87 2035 -81 2069
rect -47 2035 -41 2069
rect -87 1997 -41 2035
rect -87 1963 -81 1997
rect -47 1963 -41 1997
rect -87 1925 -41 1963
rect -87 1891 -81 1925
rect -47 1891 -41 1925
rect -87 1853 -41 1891
rect -87 1819 -81 1853
rect -47 1819 -41 1853
rect -87 1781 -41 1819
rect -87 1747 -81 1781
rect -47 1747 -41 1781
rect -87 1709 -41 1747
rect -87 1675 -81 1709
rect -47 1675 -41 1709
rect -87 1637 -41 1675
rect -87 1603 -81 1637
rect -47 1603 -41 1637
rect -87 1565 -41 1603
rect -87 1531 -81 1565
rect -47 1531 -41 1565
rect -87 1493 -41 1531
rect -87 1459 -81 1493
rect -47 1459 -41 1493
rect -87 1421 -41 1459
rect -87 1387 -81 1421
rect -47 1387 -41 1421
rect -87 1349 -41 1387
rect -87 1315 -81 1349
rect -47 1315 -41 1349
rect -87 1277 -41 1315
rect -87 1243 -81 1277
rect -47 1243 -41 1277
rect -87 1205 -41 1243
rect -87 1171 -81 1205
rect -47 1171 -41 1205
rect -87 1133 -41 1171
rect -87 1099 -81 1133
rect -47 1099 -41 1133
rect -87 1061 -41 1099
rect -87 1027 -81 1061
rect -47 1027 -41 1061
rect -87 989 -41 1027
rect -87 955 -81 989
rect -47 955 -41 989
rect -87 917 -41 955
rect -87 883 -81 917
rect -47 883 -41 917
rect -87 845 -41 883
rect -87 811 -81 845
rect -47 811 -41 845
rect -87 773 -41 811
rect -87 739 -81 773
rect -47 739 -41 773
rect -87 701 -41 739
rect -87 667 -81 701
rect -47 667 -41 701
rect -87 629 -41 667
rect -87 595 -81 629
rect -47 595 -41 629
rect -87 557 -41 595
rect -87 523 -81 557
rect -47 523 -41 557
rect -87 485 -41 523
rect -87 451 -81 485
rect -47 451 -41 485
rect -87 413 -41 451
rect -87 379 -81 413
rect -47 379 -41 413
rect -87 341 -41 379
rect -87 307 -81 341
rect -47 307 -41 341
rect -87 269 -41 307
rect -87 235 -81 269
rect -47 235 -41 269
rect -87 197 -41 235
rect -87 163 -81 197
rect -47 163 -41 197
rect -87 125 -41 163
rect -87 91 -81 125
rect -47 91 -41 125
rect -87 53 -41 91
rect -87 19 -81 53
rect -47 19 -41 53
rect -87 -19 -41 19
rect -87 -53 -81 -19
rect -47 -53 -41 -19
rect -87 -91 -41 -53
rect -87 -125 -81 -91
rect -47 -125 -41 -91
rect -87 -163 -41 -125
rect -87 -197 -81 -163
rect -47 -197 -41 -163
rect -87 -235 -41 -197
rect -87 -269 -81 -235
rect -47 -269 -41 -235
rect -87 -307 -41 -269
rect -87 -341 -81 -307
rect -47 -341 -41 -307
rect -87 -379 -41 -341
rect -87 -413 -81 -379
rect -47 -413 -41 -379
rect -87 -451 -41 -413
rect -87 -485 -81 -451
rect -47 -485 -41 -451
rect -87 -523 -41 -485
rect -87 -557 -81 -523
rect -47 -557 -41 -523
rect -87 -595 -41 -557
rect -87 -629 -81 -595
rect -47 -629 -41 -595
rect -87 -667 -41 -629
rect -87 -701 -81 -667
rect -47 -701 -41 -667
rect -87 -739 -41 -701
rect -87 -773 -81 -739
rect -47 -773 -41 -739
rect -87 -811 -41 -773
rect -87 -845 -81 -811
rect -47 -845 -41 -811
rect -87 -883 -41 -845
rect -87 -917 -81 -883
rect -47 -917 -41 -883
rect -87 -955 -41 -917
rect -87 -989 -81 -955
rect -47 -989 -41 -955
rect -87 -1027 -41 -989
rect -87 -1061 -81 -1027
rect -47 -1061 -41 -1027
rect -87 -1099 -41 -1061
rect -87 -1133 -81 -1099
rect -47 -1133 -41 -1099
rect -87 -1171 -41 -1133
rect -87 -1205 -81 -1171
rect -47 -1205 -41 -1171
rect -87 -1243 -41 -1205
rect -87 -1277 -81 -1243
rect -47 -1277 -41 -1243
rect -87 -1315 -41 -1277
rect -87 -1349 -81 -1315
rect -47 -1349 -41 -1315
rect -87 -1387 -41 -1349
rect -87 -1421 -81 -1387
rect -47 -1421 -41 -1387
rect -87 -1459 -41 -1421
rect -87 -1493 -81 -1459
rect -47 -1493 -41 -1459
rect -87 -1531 -41 -1493
rect -87 -1565 -81 -1531
rect -47 -1565 -41 -1531
rect -87 -1603 -41 -1565
rect -87 -1637 -81 -1603
rect -47 -1637 -41 -1603
rect -87 -1675 -41 -1637
rect -87 -1709 -81 -1675
rect -47 -1709 -41 -1675
rect -87 -1747 -41 -1709
rect -87 -1781 -81 -1747
rect -47 -1781 -41 -1747
rect -87 -1819 -41 -1781
rect -87 -1853 -81 -1819
rect -47 -1853 -41 -1819
rect -87 -1891 -41 -1853
rect -87 -1925 -81 -1891
rect -47 -1925 -41 -1891
rect -87 -1963 -41 -1925
rect -87 -1997 -81 -1963
rect -47 -1997 -41 -1963
rect -87 -2035 -41 -1997
rect -87 -2069 -81 -2035
rect -47 -2069 -41 -2035
rect -87 -2107 -41 -2069
rect -87 -2141 -81 -2107
rect -47 -2141 -41 -2107
rect -87 -2179 -41 -2141
rect -87 -2213 -81 -2179
rect -47 -2213 -41 -2179
rect -87 -2251 -41 -2213
rect -87 -2285 -81 -2251
rect -47 -2285 -41 -2251
rect -87 -2323 -41 -2285
rect -87 -2357 -81 -2323
rect -47 -2357 -41 -2323
rect -87 -2395 -41 -2357
rect -87 -2429 -81 -2395
rect -47 -2429 -41 -2395
rect -87 -2467 -41 -2429
rect -87 -2501 -81 -2467
rect -47 -2501 -41 -2467
rect -87 -2539 -41 -2501
rect -87 -2573 -81 -2539
rect -47 -2573 -41 -2539
rect -87 -2611 -41 -2573
rect -87 -2645 -81 -2611
rect -47 -2645 -41 -2611
rect -87 -2683 -41 -2645
rect -87 -2717 -81 -2683
rect -47 -2717 -41 -2683
rect -87 -2755 -41 -2717
rect -87 -2789 -81 -2755
rect -47 -2789 -41 -2755
rect -87 -2827 -41 -2789
rect -87 -2861 -81 -2827
rect -47 -2861 -41 -2827
rect -87 -2899 -41 -2861
rect -87 -2933 -81 -2899
rect -47 -2933 -41 -2899
rect -87 -2971 -41 -2933
rect -87 -3005 -81 -2971
rect -47 -3005 -41 -2971
rect -87 -3043 -41 -3005
rect -87 -3077 -81 -3043
rect -47 -3077 -41 -3043
rect -87 -3115 -41 -3077
rect -87 -3149 -81 -3115
rect -47 -3149 -41 -3115
rect -87 -3187 -41 -3149
rect -87 -3221 -81 -3187
rect -47 -3221 -41 -3187
rect -87 -3259 -41 -3221
rect -87 -3293 -81 -3259
rect -47 -3293 -41 -3259
rect -87 -3331 -41 -3293
rect -87 -3365 -81 -3331
rect -47 -3365 -41 -3331
rect -87 -3403 -41 -3365
rect -87 -3437 -81 -3403
rect -47 -3437 -41 -3403
rect -87 -3475 -41 -3437
rect -87 -3509 -81 -3475
rect -47 -3509 -41 -3475
rect -87 -3547 -41 -3509
rect -87 -3581 -81 -3547
rect -47 -3581 -41 -3547
rect -87 -3619 -41 -3581
rect -87 -3653 -81 -3619
rect -47 -3653 -41 -3619
rect -87 -3691 -41 -3653
rect -87 -3725 -81 -3691
rect -47 -3725 -41 -3691
rect -87 -3763 -41 -3725
rect -87 -3797 -81 -3763
rect -47 -3797 -41 -3763
rect -87 -3835 -41 -3797
rect -87 -3869 -81 -3835
rect -47 -3869 -41 -3835
rect -87 -3907 -41 -3869
rect -87 -3941 -81 -3907
rect -47 -3941 -41 -3907
rect -87 -3979 -41 -3941
rect -87 -4013 -81 -3979
rect -47 -4013 -41 -3979
rect -87 -4051 -41 -4013
rect -87 -4085 -81 -4051
rect -47 -4085 -41 -4051
rect -87 -4123 -41 -4085
rect -87 -4157 -81 -4123
rect -47 -4157 -41 -4123
rect -87 -4195 -41 -4157
rect -87 -4229 -81 -4195
rect -47 -4229 -41 -4195
rect -87 -4267 -41 -4229
rect -87 -4301 -81 -4267
rect -47 -4301 -41 -4267
rect -87 -4339 -41 -4301
rect -87 -4373 -81 -4339
rect -47 -4373 -41 -4339
rect -87 -4411 -41 -4373
rect -87 -4445 -81 -4411
rect -47 -4445 -41 -4411
rect -87 -4483 -41 -4445
rect -87 -4517 -81 -4483
rect -47 -4517 -41 -4483
rect -87 -4555 -41 -4517
rect -87 -4589 -81 -4555
rect -47 -4589 -41 -4555
rect -87 -4627 -41 -4589
rect -87 -4661 -81 -4627
rect -47 -4661 -41 -4627
rect -87 -4699 -41 -4661
rect -87 -4733 -81 -4699
rect -47 -4733 -41 -4699
rect -87 -4771 -41 -4733
rect -87 -4805 -81 -4771
rect -47 -4805 -41 -4771
rect -87 -4843 -41 -4805
rect -87 -4877 -81 -4843
rect -47 -4877 -41 -4843
rect -87 -4915 -41 -4877
rect -87 -4949 -81 -4915
rect -47 -4949 -41 -4915
rect -87 -4987 -41 -4949
rect -87 -5021 -81 -4987
rect -47 -5021 -41 -4987
rect -87 -5059 -41 -5021
rect -87 -5093 -81 -5059
rect -47 -5093 -41 -5059
rect -87 -5131 -41 -5093
rect -87 -5165 -81 -5131
rect -47 -5165 -41 -5131
rect -87 -5203 -41 -5165
rect -87 -5237 -81 -5203
rect -47 -5237 -41 -5203
rect -87 -5275 -41 -5237
rect -87 -5309 -81 -5275
rect -47 -5309 -41 -5275
rect -87 -5347 -41 -5309
rect -87 -5381 -81 -5347
rect -47 -5381 -41 -5347
rect -87 -5419 -41 -5381
rect -87 -5453 -81 -5419
rect -47 -5453 -41 -5419
rect -87 -5491 -41 -5453
rect -87 -5525 -81 -5491
rect -47 -5525 -41 -5491
rect -87 -5563 -41 -5525
rect -87 -5597 -81 -5563
rect -47 -5597 -41 -5563
rect -87 -5635 -41 -5597
rect -87 -5669 -81 -5635
rect -47 -5669 -41 -5635
rect -87 -5707 -41 -5669
rect -87 -5741 -81 -5707
rect -47 -5741 -41 -5707
rect -87 -5779 -41 -5741
rect -87 -5813 -81 -5779
rect -47 -5813 -41 -5779
rect -87 -5851 -41 -5813
rect -87 -5885 -81 -5851
rect -47 -5885 -41 -5851
rect -87 -5923 -41 -5885
rect -87 -5957 -81 -5923
rect -47 -5957 -41 -5923
rect -87 -5995 -41 -5957
rect -87 -6029 -81 -5995
rect -47 -6029 -41 -5995
rect -87 -6067 -41 -6029
rect -87 -6101 -81 -6067
rect -47 -6101 -41 -6067
rect -87 -6139 -41 -6101
rect -87 -6173 -81 -6139
rect -47 -6173 -41 -6139
rect -87 -6211 -41 -6173
rect -87 -6245 -81 -6211
rect -47 -6245 -41 -6211
rect -87 -6283 -41 -6245
rect -87 -6317 -81 -6283
rect -47 -6317 -41 -6283
rect -87 -6355 -41 -6317
rect -87 -6389 -81 -6355
rect -47 -6389 -41 -6355
rect -87 -6427 -41 -6389
rect -87 -6461 -81 -6427
rect -47 -6461 -41 -6427
rect -87 -6499 -41 -6461
rect -87 -6533 -81 -6499
rect -47 -6533 -41 -6499
rect -87 -6571 -41 -6533
rect -87 -6605 -81 -6571
rect -47 -6605 -41 -6571
rect -87 -6643 -41 -6605
rect -87 -6677 -81 -6643
rect -47 -6677 -41 -6643
rect -87 -6715 -41 -6677
rect -87 -6749 -81 -6715
rect -47 -6749 -41 -6715
rect -87 -6787 -41 -6749
rect -87 -6821 -81 -6787
rect -47 -6821 -41 -6787
rect -87 -6859 -41 -6821
rect -87 -6893 -81 -6859
rect -47 -6893 -41 -6859
rect -87 -6931 -41 -6893
rect -87 -6965 -81 -6931
rect -47 -6965 -41 -6931
rect -87 -7003 -41 -6965
rect -87 -7037 -81 -7003
rect -47 -7037 -41 -7003
rect -87 -7075 -41 -7037
rect -87 -7109 -81 -7075
rect -47 -7109 -41 -7075
rect -87 -7147 -41 -7109
rect -87 -7181 -81 -7147
rect -47 -7181 -41 -7147
rect -87 -7219 -41 -7181
rect -87 -7253 -81 -7219
rect -47 -7253 -41 -7219
rect -87 -7291 -41 -7253
rect -87 -7325 -81 -7291
rect -47 -7325 -41 -7291
rect -87 -7363 -41 -7325
rect -87 -7397 -81 -7363
rect -47 -7397 -41 -7363
rect -87 -7435 -41 -7397
rect -87 -7469 -81 -7435
rect -47 -7469 -41 -7435
rect -87 -7507 -41 -7469
rect -87 -7541 -81 -7507
rect -47 -7541 -41 -7507
rect -87 -7579 -41 -7541
rect -87 -7613 -81 -7579
rect -47 -7613 -41 -7579
rect -87 -7651 -41 -7613
rect -87 -7685 -81 -7651
rect -47 -7685 -41 -7651
rect -87 -7723 -41 -7685
rect -87 -7757 -81 -7723
rect -47 -7757 -41 -7723
rect -87 -7795 -41 -7757
rect -87 -7829 -81 -7795
rect -47 -7829 -41 -7795
rect -87 -7867 -41 -7829
rect -87 -7901 -81 -7867
rect -47 -7901 -41 -7867
rect -87 -7939 -41 -7901
rect -87 -7973 -81 -7939
rect -47 -7973 -41 -7939
rect -87 -8000 -41 -7973
rect 41 7973 87 8000
rect 41 7939 47 7973
rect 81 7939 87 7973
rect 41 7901 87 7939
rect 41 7867 47 7901
rect 81 7867 87 7901
rect 41 7829 87 7867
rect 41 7795 47 7829
rect 81 7795 87 7829
rect 41 7757 87 7795
rect 41 7723 47 7757
rect 81 7723 87 7757
rect 41 7685 87 7723
rect 41 7651 47 7685
rect 81 7651 87 7685
rect 41 7613 87 7651
rect 41 7579 47 7613
rect 81 7579 87 7613
rect 41 7541 87 7579
rect 41 7507 47 7541
rect 81 7507 87 7541
rect 41 7469 87 7507
rect 41 7435 47 7469
rect 81 7435 87 7469
rect 41 7397 87 7435
rect 41 7363 47 7397
rect 81 7363 87 7397
rect 41 7325 87 7363
rect 41 7291 47 7325
rect 81 7291 87 7325
rect 41 7253 87 7291
rect 41 7219 47 7253
rect 81 7219 87 7253
rect 41 7181 87 7219
rect 41 7147 47 7181
rect 81 7147 87 7181
rect 41 7109 87 7147
rect 41 7075 47 7109
rect 81 7075 87 7109
rect 41 7037 87 7075
rect 41 7003 47 7037
rect 81 7003 87 7037
rect 41 6965 87 7003
rect 41 6931 47 6965
rect 81 6931 87 6965
rect 41 6893 87 6931
rect 41 6859 47 6893
rect 81 6859 87 6893
rect 41 6821 87 6859
rect 41 6787 47 6821
rect 81 6787 87 6821
rect 41 6749 87 6787
rect 41 6715 47 6749
rect 81 6715 87 6749
rect 41 6677 87 6715
rect 41 6643 47 6677
rect 81 6643 87 6677
rect 41 6605 87 6643
rect 41 6571 47 6605
rect 81 6571 87 6605
rect 41 6533 87 6571
rect 41 6499 47 6533
rect 81 6499 87 6533
rect 41 6461 87 6499
rect 41 6427 47 6461
rect 81 6427 87 6461
rect 41 6389 87 6427
rect 41 6355 47 6389
rect 81 6355 87 6389
rect 41 6317 87 6355
rect 41 6283 47 6317
rect 81 6283 87 6317
rect 41 6245 87 6283
rect 41 6211 47 6245
rect 81 6211 87 6245
rect 41 6173 87 6211
rect 41 6139 47 6173
rect 81 6139 87 6173
rect 41 6101 87 6139
rect 41 6067 47 6101
rect 81 6067 87 6101
rect 41 6029 87 6067
rect 41 5995 47 6029
rect 81 5995 87 6029
rect 41 5957 87 5995
rect 41 5923 47 5957
rect 81 5923 87 5957
rect 41 5885 87 5923
rect 41 5851 47 5885
rect 81 5851 87 5885
rect 41 5813 87 5851
rect 41 5779 47 5813
rect 81 5779 87 5813
rect 41 5741 87 5779
rect 41 5707 47 5741
rect 81 5707 87 5741
rect 41 5669 87 5707
rect 41 5635 47 5669
rect 81 5635 87 5669
rect 41 5597 87 5635
rect 41 5563 47 5597
rect 81 5563 87 5597
rect 41 5525 87 5563
rect 41 5491 47 5525
rect 81 5491 87 5525
rect 41 5453 87 5491
rect 41 5419 47 5453
rect 81 5419 87 5453
rect 41 5381 87 5419
rect 41 5347 47 5381
rect 81 5347 87 5381
rect 41 5309 87 5347
rect 41 5275 47 5309
rect 81 5275 87 5309
rect 41 5237 87 5275
rect 41 5203 47 5237
rect 81 5203 87 5237
rect 41 5165 87 5203
rect 41 5131 47 5165
rect 81 5131 87 5165
rect 41 5093 87 5131
rect 41 5059 47 5093
rect 81 5059 87 5093
rect 41 5021 87 5059
rect 41 4987 47 5021
rect 81 4987 87 5021
rect 41 4949 87 4987
rect 41 4915 47 4949
rect 81 4915 87 4949
rect 41 4877 87 4915
rect 41 4843 47 4877
rect 81 4843 87 4877
rect 41 4805 87 4843
rect 41 4771 47 4805
rect 81 4771 87 4805
rect 41 4733 87 4771
rect 41 4699 47 4733
rect 81 4699 87 4733
rect 41 4661 87 4699
rect 41 4627 47 4661
rect 81 4627 87 4661
rect 41 4589 87 4627
rect 41 4555 47 4589
rect 81 4555 87 4589
rect 41 4517 87 4555
rect 41 4483 47 4517
rect 81 4483 87 4517
rect 41 4445 87 4483
rect 41 4411 47 4445
rect 81 4411 87 4445
rect 41 4373 87 4411
rect 41 4339 47 4373
rect 81 4339 87 4373
rect 41 4301 87 4339
rect 41 4267 47 4301
rect 81 4267 87 4301
rect 41 4229 87 4267
rect 41 4195 47 4229
rect 81 4195 87 4229
rect 41 4157 87 4195
rect 41 4123 47 4157
rect 81 4123 87 4157
rect 41 4085 87 4123
rect 41 4051 47 4085
rect 81 4051 87 4085
rect 41 4013 87 4051
rect 41 3979 47 4013
rect 81 3979 87 4013
rect 41 3941 87 3979
rect 41 3907 47 3941
rect 81 3907 87 3941
rect 41 3869 87 3907
rect 41 3835 47 3869
rect 81 3835 87 3869
rect 41 3797 87 3835
rect 41 3763 47 3797
rect 81 3763 87 3797
rect 41 3725 87 3763
rect 41 3691 47 3725
rect 81 3691 87 3725
rect 41 3653 87 3691
rect 41 3619 47 3653
rect 81 3619 87 3653
rect 41 3581 87 3619
rect 41 3547 47 3581
rect 81 3547 87 3581
rect 41 3509 87 3547
rect 41 3475 47 3509
rect 81 3475 87 3509
rect 41 3437 87 3475
rect 41 3403 47 3437
rect 81 3403 87 3437
rect 41 3365 87 3403
rect 41 3331 47 3365
rect 81 3331 87 3365
rect 41 3293 87 3331
rect 41 3259 47 3293
rect 81 3259 87 3293
rect 41 3221 87 3259
rect 41 3187 47 3221
rect 81 3187 87 3221
rect 41 3149 87 3187
rect 41 3115 47 3149
rect 81 3115 87 3149
rect 41 3077 87 3115
rect 41 3043 47 3077
rect 81 3043 87 3077
rect 41 3005 87 3043
rect 41 2971 47 3005
rect 81 2971 87 3005
rect 41 2933 87 2971
rect 41 2899 47 2933
rect 81 2899 87 2933
rect 41 2861 87 2899
rect 41 2827 47 2861
rect 81 2827 87 2861
rect 41 2789 87 2827
rect 41 2755 47 2789
rect 81 2755 87 2789
rect 41 2717 87 2755
rect 41 2683 47 2717
rect 81 2683 87 2717
rect 41 2645 87 2683
rect 41 2611 47 2645
rect 81 2611 87 2645
rect 41 2573 87 2611
rect 41 2539 47 2573
rect 81 2539 87 2573
rect 41 2501 87 2539
rect 41 2467 47 2501
rect 81 2467 87 2501
rect 41 2429 87 2467
rect 41 2395 47 2429
rect 81 2395 87 2429
rect 41 2357 87 2395
rect 41 2323 47 2357
rect 81 2323 87 2357
rect 41 2285 87 2323
rect 41 2251 47 2285
rect 81 2251 87 2285
rect 41 2213 87 2251
rect 41 2179 47 2213
rect 81 2179 87 2213
rect 41 2141 87 2179
rect 41 2107 47 2141
rect 81 2107 87 2141
rect 41 2069 87 2107
rect 41 2035 47 2069
rect 81 2035 87 2069
rect 41 1997 87 2035
rect 41 1963 47 1997
rect 81 1963 87 1997
rect 41 1925 87 1963
rect 41 1891 47 1925
rect 81 1891 87 1925
rect 41 1853 87 1891
rect 41 1819 47 1853
rect 81 1819 87 1853
rect 41 1781 87 1819
rect 41 1747 47 1781
rect 81 1747 87 1781
rect 41 1709 87 1747
rect 41 1675 47 1709
rect 81 1675 87 1709
rect 41 1637 87 1675
rect 41 1603 47 1637
rect 81 1603 87 1637
rect 41 1565 87 1603
rect 41 1531 47 1565
rect 81 1531 87 1565
rect 41 1493 87 1531
rect 41 1459 47 1493
rect 81 1459 87 1493
rect 41 1421 87 1459
rect 41 1387 47 1421
rect 81 1387 87 1421
rect 41 1349 87 1387
rect 41 1315 47 1349
rect 81 1315 87 1349
rect 41 1277 87 1315
rect 41 1243 47 1277
rect 81 1243 87 1277
rect 41 1205 87 1243
rect 41 1171 47 1205
rect 81 1171 87 1205
rect 41 1133 87 1171
rect 41 1099 47 1133
rect 81 1099 87 1133
rect 41 1061 87 1099
rect 41 1027 47 1061
rect 81 1027 87 1061
rect 41 989 87 1027
rect 41 955 47 989
rect 81 955 87 989
rect 41 917 87 955
rect 41 883 47 917
rect 81 883 87 917
rect 41 845 87 883
rect 41 811 47 845
rect 81 811 87 845
rect 41 773 87 811
rect 41 739 47 773
rect 81 739 87 773
rect 41 701 87 739
rect 41 667 47 701
rect 81 667 87 701
rect 41 629 87 667
rect 41 595 47 629
rect 81 595 87 629
rect 41 557 87 595
rect 41 523 47 557
rect 81 523 87 557
rect 41 485 87 523
rect 41 451 47 485
rect 81 451 87 485
rect 41 413 87 451
rect 41 379 47 413
rect 81 379 87 413
rect 41 341 87 379
rect 41 307 47 341
rect 81 307 87 341
rect 41 269 87 307
rect 41 235 47 269
rect 81 235 87 269
rect 41 197 87 235
rect 41 163 47 197
rect 81 163 87 197
rect 41 125 87 163
rect 41 91 47 125
rect 81 91 87 125
rect 41 53 87 91
rect 41 19 47 53
rect 81 19 87 53
rect 41 -19 87 19
rect 41 -53 47 -19
rect 81 -53 87 -19
rect 41 -91 87 -53
rect 41 -125 47 -91
rect 81 -125 87 -91
rect 41 -163 87 -125
rect 41 -197 47 -163
rect 81 -197 87 -163
rect 41 -235 87 -197
rect 41 -269 47 -235
rect 81 -269 87 -235
rect 41 -307 87 -269
rect 41 -341 47 -307
rect 81 -341 87 -307
rect 41 -379 87 -341
rect 41 -413 47 -379
rect 81 -413 87 -379
rect 41 -451 87 -413
rect 41 -485 47 -451
rect 81 -485 87 -451
rect 41 -523 87 -485
rect 41 -557 47 -523
rect 81 -557 87 -523
rect 41 -595 87 -557
rect 41 -629 47 -595
rect 81 -629 87 -595
rect 41 -667 87 -629
rect 41 -701 47 -667
rect 81 -701 87 -667
rect 41 -739 87 -701
rect 41 -773 47 -739
rect 81 -773 87 -739
rect 41 -811 87 -773
rect 41 -845 47 -811
rect 81 -845 87 -811
rect 41 -883 87 -845
rect 41 -917 47 -883
rect 81 -917 87 -883
rect 41 -955 87 -917
rect 41 -989 47 -955
rect 81 -989 87 -955
rect 41 -1027 87 -989
rect 41 -1061 47 -1027
rect 81 -1061 87 -1027
rect 41 -1099 87 -1061
rect 41 -1133 47 -1099
rect 81 -1133 87 -1099
rect 41 -1171 87 -1133
rect 41 -1205 47 -1171
rect 81 -1205 87 -1171
rect 41 -1243 87 -1205
rect 41 -1277 47 -1243
rect 81 -1277 87 -1243
rect 41 -1315 87 -1277
rect 41 -1349 47 -1315
rect 81 -1349 87 -1315
rect 41 -1387 87 -1349
rect 41 -1421 47 -1387
rect 81 -1421 87 -1387
rect 41 -1459 87 -1421
rect 41 -1493 47 -1459
rect 81 -1493 87 -1459
rect 41 -1531 87 -1493
rect 41 -1565 47 -1531
rect 81 -1565 87 -1531
rect 41 -1603 87 -1565
rect 41 -1637 47 -1603
rect 81 -1637 87 -1603
rect 41 -1675 87 -1637
rect 41 -1709 47 -1675
rect 81 -1709 87 -1675
rect 41 -1747 87 -1709
rect 41 -1781 47 -1747
rect 81 -1781 87 -1747
rect 41 -1819 87 -1781
rect 41 -1853 47 -1819
rect 81 -1853 87 -1819
rect 41 -1891 87 -1853
rect 41 -1925 47 -1891
rect 81 -1925 87 -1891
rect 41 -1963 87 -1925
rect 41 -1997 47 -1963
rect 81 -1997 87 -1963
rect 41 -2035 87 -1997
rect 41 -2069 47 -2035
rect 81 -2069 87 -2035
rect 41 -2107 87 -2069
rect 41 -2141 47 -2107
rect 81 -2141 87 -2107
rect 41 -2179 87 -2141
rect 41 -2213 47 -2179
rect 81 -2213 87 -2179
rect 41 -2251 87 -2213
rect 41 -2285 47 -2251
rect 81 -2285 87 -2251
rect 41 -2323 87 -2285
rect 41 -2357 47 -2323
rect 81 -2357 87 -2323
rect 41 -2395 87 -2357
rect 41 -2429 47 -2395
rect 81 -2429 87 -2395
rect 41 -2467 87 -2429
rect 41 -2501 47 -2467
rect 81 -2501 87 -2467
rect 41 -2539 87 -2501
rect 41 -2573 47 -2539
rect 81 -2573 87 -2539
rect 41 -2611 87 -2573
rect 41 -2645 47 -2611
rect 81 -2645 87 -2611
rect 41 -2683 87 -2645
rect 41 -2717 47 -2683
rect 81 -2717 87 -2683
rect 41 -2755 87 -2717
rect 41 -2789 47 -2755
rect 81 -2789 87 -2755
rect 41 -2827 87 -2789
rect 41 -2861 47 -2827
rect 81 -2861 87 -2827
rect 41 -2899 87 -2861
rect 41 -2933 47 -2899
rect 81 -2933 87 -2899
rect 41 -2971 87 -2933
rect 41 -3005 47 -2971
rect 81 -3005 87 -2971
rect 41 -3043 87 -3005
rect 41 -3077 47 -3043
rect 81 -3077 87 -3043
rect 41 -3115 87 -3077
rect 41 -3149 47 -3115
rect 81 -3149 87 -3115
rect 41 -3187 87 -3149
rect 41 -3221 47 -3187
rect 81 -3221 87 -3187
rect 41 -3259 87 -3221
rect 41 -3293 47 -3259
rect 81 -3293 87 -3259
rect 41 -3331 87 -3293
rect 41 -3365 47 -3331
rect 81 -3365 87 -3331
rect 41 -3403 87 -3365
rect 41 -3437 47 -3403
rect 81 -3437 87 -3403
rect 41 -3475 87 -3437
rect 41 -3509 47 -3475
rect 81 -3509 87 -3475
rect 41 -3547 87 -3509
rect 41 -3581 47 -3547
rect 81 -3581 87 -3547
rect 41 -3619 87 -3581
rect 41 -3653 47 -3619
rect 81 -3653 87 -3619
rect 41 -3691 87 -3653
rect 41 -3725 47 -3691
rect 81 -3725 87 -3691
rect 41 -3763 87 -3725
rect 41 -3797 47 -3763
rect 81 -3797 87 -3763
rect 41 -3835 87 -3797
rect 41 -3869 47 -3835
rect 81 -3869 87 -3835
rect 41 -3907 87 -3869
rect 41 -3941 47 -3907
rect 81 -3941 87 -3907
rect 41 -3979 87 -3941
rect 41 -4013 47 -3979
rect 81 -4013 87 -3979
rect 41 -4051 87 -4013
rect 41 -4085 47 -4051
rect 81 -4085 87 -4051
rect 41 -4123 87 -4085
rect 41 -4157 47 -4123
rect 81 -4157 87 -4123
rect 41 -4195 87 -4157
rect 41 -4229 47 -4195
rect 81 -4229 87 -4195
rect 41 -4267 87 -4229
rect 41 -4301 47 -4267
rect 81 -4301 87 -4267
rect 41 -4339 87 -4301
rect 41 -4373 47 -4339
rect 81 -4373 87 -4339
rect 41 -4411 87 -4373
rect 41 -4445 47 -4411
rect 81 -4445 87 -4411
rect 41 -4483 87 -4445
rect 41 -4517 47 -4483
rect 81 -4517 87 -4483
rect 41 -4555 87 -4517
rect 41 -4589 47 -4555
rect 81 -4589 87 -4555
rect 41 -4627 87 -4589
rect 41 -4661 47 -4627
rect 81 -4661 87 -4627
rect 41 -4699 87 -4661
rect 41 -4733 47 -4699
rect 81 -4733 87 -4699
rect 41 -4771 87 -4733
rect 41 -4805 47 -4771
rect 81 -4805 87 -4771
rect 41 -4843 87 -4805
rect 41 -4877 47 -4843
rect 81 -4877 87 -4843
rect 41 -4915 87 -4877
rect 41 -4949 47 -4915
rect 81 -4949 87 -4915
rect 41 -4987 87 -4949
rect 41 -5021 47 -4987
rect 81 -5021 87 -4987
rect 41 -5059 87 -5021
rect 41 -5093 47 -5059
rect 81 -5093 87 -5059
rect 41 -5131 87 -5093
rect 41 -5165 47 -5131
rect 81 -5165 87 -5131
rect 41 -5203 87 -5165
rect 41 -5237 47 -5203
rect 81 -5237 87 -5203
rect 41 -5275 87 -5237
rect 41 -5309 47 -5275
rect 81 -5309 87 -5275
rect 41 -5347 87 -5309
rect 41 -5381 47 -5347
rect 81 -5381 87 -5347
rect 41 -5419 87 -5381
rect 41 -5453 47 -5419
rect 81 -5453 87 -5419
rect 41 -5491 87 -5453
rect 41 -5525 47 -5491
rect 81 -5525 87 -5491
rect 41 -5563 87 -5525
rect 41 -5597 47 -5563
rect 81 -5597 87 -5563
rect 41 -5635 87 -5597
rect 41 -5669 47 -5635
rect 81 -5669 87 -5635
rect 41 -5707 87 -5669
rect 41 -5741 47 -5707
rect 81 -5741 87 -5707
rect 41 -5779 87 -5741
rect 41 -5813 47 -5779
rect 81 -5813 87 -5779
rect 41 -5851 87 -5813
rect 41 -5885 47 -5851
rect 81 -5885 87 -5851
rect 41 -5923 87 -5885
rect 41 -5957 47 -5923
rect 81 -5957 87 -5923
rect 41 -5995 87 -5957
rect 41 -6029 47 -5995
rect 81 -6029 87 -5995
rect 41 -6067 87 -6029
rect 41 -6101 47 -6067
rect 81 -6101 87 -6067
rect 41 -6139 87 -6101
rect 41 -6173 47 -6139
rect 81 -6173 87 -6139
rect 41 -6211 87 -6173
rect 41 -6245 47 -6211
rect 81 -6245 87 -6211
rect 41 -6283 87 -6245
rect 41 -6317 47 -6283
rect 81 -6317 87 -6283
rect 41 -6355 87 -6317
rect 41 -6389 47 -6355
rect 81 -6389 87 -6355
rect 41 -6427 87 -6389
rect 41 -6461 47 -6427
rect 81 -6461 87 -6427
rect 41 -6499 87 -6461
rect 41 -6533 47 -6499
rect 81 -6533 87 -6499
rect 41 -6571 87 -6533
rect 41 -6605 47 -6571
rect 81 -6605 87 -6571
rect 41 -6643 87 -6605
rect 41 -6677 47 -6643
rect 81 -6677 87 -6643
rect 41 -6715 87 -6677
rect 41 -6749 47 -6715
rect 81 -6749 87 -6715
rect 41 -6787 87 -6749
rect 41 -6821 47 -6787
rect 81 -6821 87 -6787
rect 41 -6859 87 -6821
rect 41 -6893 47 -6859
rect 81 -6893 87 -6859
rect 41 -6931 87 -6893
rect 41 -6965 47 -6931
rect 81 -6965 87 -6931
rect 41 -7003 87 -6965
rect 41 -7037 47 -7003
rect 81 -7037 87 -7003
rect 41 -7075 87 -7037
rect 41 -7109 47 -7075
rect 81 -7109 87 -7075
rect 41 -7147 87 -7109
rect 41 -7181 47 -7147
rect 81 -7181 87 -7147
rect 41 -7219 87 -7181
rect 41 -7253 47 -7219
rect 81 -7253 87 -7219
rect 41 -7291 87 -7253
rect 41 -7325 47 -7291
rect 81 -7325 87 -7291
rect 41 -7363 87 -7325
rect 41 -7397 47 -7363
rect 81 -7397 87 -7363
rect 41 -7435 87 -7397
rect 41 -7469 47 -7435
rect 81 -7469 87 -7435
rect 41 -7507 87 -7469
rect 41 -7541 47 -7507
rect 81 -7541 87 -7507
rect 41 -7579 87 -7541
rect 41 -7613 47 -7579
rect 81 -7613 87 -7579
rect 41 -7651 87 -7613
rect 41 -7685 47 -7651
rect 81 -7685 87 -7651
rect 41 -7723 87 -7685
rect 41 -7757 47 -7723
rect 81 -7757 87 -7723
rect 41 -7795 87 -7757
rect 41 -7829 47 -7795
rect 81 -7829 87 -7795
rect 41 -7867 87 -7829
rect 41 -7901 47 -7867
rect 81 -7901 87 -7867
rect 41 -7939 87 -7901
rect 41 -7973 47 -7939
rect 81 -7973 87 -7939
rect 41 -8000 87 -7973
rect -31 -8038 31 -8032
rect -31 -8072 -17 -8038
rect 17 -8072 31 -8038
rect -31 -8078 31 -8072
<< properties >>
string FIXED_BBOX -178 -8157 178 8157
<< end >>
