magic
tech sky130A
magscale 1 2
timestamp 1635855079
<< locali >>
rect -18 16312 9156 16348
rect -18 -18 9150 18
<< metal1 >>
rect 144 16252 9216 16344
rect 142 16240 9216 16252
rect 142 16214 8992 16240
rect 142 16208 672 16214
rect -238 16168 132 16172
rect 946 16168 1050 16176
rect -238 16116 38 16168
rect 90 16116 132 16168
rect -238 16100 132 16116
rect 482 16164 586 16168
rect 482 16112 494 16164
rect 546 16112 586 16164
rect 946 16116 956 16168
rect 1008 16116 1050 16168
rect 946 16112 1050 16116
rect 1402 16164 1506 16172
rect 1402 16112 1414 16164
rect 1466 16112 1506 16164
rect 1868 16170 1972 16176
rect 1868 16118 1878 16170
rect 1930 16118 1972 16170
rect 1868 16112 1972 16118
rect 2328 16174 2432 16180
rect 2328 16122 2336 16174
rect 2388 16122 2432 16174
rect 2328 16116 2432 16122
rect 2796 16174 2900 16182
rect 2796 16122 2806 16174
rect 2858 16122 2900 16174
rect 3254 16176 3358 16186
rect 3254 16124 3264 16176
rect 3316 16124 3358 16176
rect 3254 16122 3358 16124
rect 3716 16176 3820 16184
rect 3716 16124 3728 16176
rect 3780 16124 3820 16176
rect 2796 16118 2900 16122
rect 3716 16120 3820 16124
rect 4178 16176 4282 16184
rect 4178 16124 4190 16176
rect 4242 16124 4282 16176
rect 4178 16120 4282 16124
rect 4640 16176 4744 16182
rect 4640 16124 4652 16176
rect 4704 16124 4744 16176
rect 4640 16118 4744 16124
rect 5100 16176 5204 16186
rect 5100 16124 5112 16176
rect 5164 16124 5204 16176
rect 5100 16122 5204 16124
rect 5564 16176 5668 16184
rect 5564 16124 5576 16176
rect 5628 16124 5668 16176
rect 5564 16120 5668 16124
rect 6026 16180 6130 16186
rect 6026 16128 6036 16180
rect 6088 16128 6130 16180
rect 6026 16122 6130 16128
rect 6484 16174 6588 16184
rect 6484 16122 6502 16174
rect 6554 16122 6588 16174
rect 6948 16176 7052 16186
rect 6948 16124 6960 16176
rect 7012 16124 7052 16176
rect 6948 16122 7052 16124
rect 7408 16178 7512 16186
rect 7408 16126 7426 16178
rect 7478 16126 7512 16178
rect 7408 16122 7512 16126
rect 7872 16178 7976 16186
rect 7872 16126 7888 16178
rect 7940 16126 7976 16178
rect 7872 16122 7976 16126
rect 8334 16178 8438 16186
rect 8334 16126 8348 16178
rect 8400 16126 8438 16178
rect 8334 16122 8438 16126
rect 8794 16172 8898 16180
rect 6484 16120 6588 16122
rect 8794 16120 8810 16172
rect 8862 16120 8898 16172
rect 8794 16116 8898 16120
rect 482 16104 586 16112
rect 1402 16108 1506 16112
rect 224 229 340 236
rect 224 177 274 229
rect 326 177 340 229
rect 224 162 340 177
rect 684 231 800 240
rect 684 179 732 231
rect 784 179 800 231
rect 684 166 800 179
rect 1142 235 1258 240
rect 1142 183 1198 235
rect 1250 183 1258 235
rect 1142 166 1258 183
rect 1606 233 1722 240
rect 1606 181 1654 233
rect 1706 181 1722 233
rect 1606 166 1722 181
rect 2066 231 2182 240
rect 2066 179 2114 231
rect 2166 179 2182 231
rect 2066 166 2182 179
rect 2528 235 2644 240
rect 2528 183 2582 235
rect 2634 183 2644 235
rect 2528 166 2644 183
rect 2990 229 3106 240
rect 2990 177 3046 229
rect 3098 177 3106 229
rect 2990 166 3106 177
rect 3452 231 3568 240
rect 3452 179 3508 231
rect 3560 179 3568 231
rect 3452 166 3568 179
rect 3914 233 4030 240
rect 3914 181 3968 233
rect 4020 181 4030 233
rect 3914 166 4030 181
rect 4376 233 4492 240
rect 4376 181 4428 233
rect 4480 181 4492 233
rect 4376 166 4492 181
rect 4840 229 4956 240
rect 4840 177 4888 229
rect 4940 177 4956 229
rect 4840 166 4956 177
rect 5302 231 5418 240
rect 5302 179 5352 231
rect 5404 179 5418 231
rect 5302 166 5418 179
rect 5762 229 5878 236
rect 5762 177 5814 229
rect 5866 177 5878 229
rect 5762 162 5878 177
rect 6224 231 6340 240
rect 6224 179 6276 231
rect 6328 179 6340 231
rect 6224 166 6340 179
rect 6688 233 6804 242
rect 6688 181 6742 233
rect 6794 181 6804 233
rect 6688 168 6804 181
rect 7150 233 7266 238
rect 7150 181 7202 233
rect 7254 181 7266 233
rect 7150 164 7266 181
rect 7612 233 7728 238
rect 7612 181 7664 233
rect 7716 181 7728 233
rect 7612 164 7728 181
rect 8070 231 8186 238
rect 8070 179 8126 231
rect 8178 179 8186 231
rect 8070 164 8186 179
rect 8536 231 8652 240
rect 8536 179 8586 231
rect 8638 179 8652 231
rect 8536 166 8652 179
rect 8996 231 9112 238
rect 8996 179 9056 231
rect 9108 179 9112 231
rect 8996 164 9112 179
rect 140 -278 9006 126
<< via1 >>
rect 38 16116 90 16168
rect 494 16112 546 16164
rect 956 16116 1008 16168
rect 1414 16112 1466 16164
rect 1878 16118 1930 16170
rect 2336 16122 2388 16174
rect 2806 16122 2858 16174
rect 3264 16124 3316 16176
rect 3728 16124 3780 16176
rect 4190 16124 4242 16176
rect 4652 16124 4704 16176
rect 5112 16124 5164 16176
rect 5576 16124 5628 16176
rect 6036 16128 6088 16180
rect 6502 16122 6554 16174
rect 6960 16124 7012 16176
rect 7426 16126 7478 16178
rect 7888 16126 7940 16178
rect 8348 16126 8400 16178
rect 8810 16120 8862 16172
rect 274 177 326 229
rect 732 179 784 231
rect 1198 183 1250 235
rect 1654 181 1706 233
rect 2114 179 2166 231
rect 2582 183 2634 235
rect 3046 177 3098 229
rect 3508 179 3560 231
rect 3968 181 4020 233
rect 4428 181 4480 233
rect 4888 177 4940 229
rect 5352 179 5404 231
rect 5814 177 5866 229
rect 6276 179 6328 231
rect 6742 181 6794 233
rect 7202 181 7254 233
rect 7664 181 7716 233
rect 8126 179 8178 231
rect 8586 179 8638 231
rect 9056 179 9108 231
<< metal2 >>
rect 22 16176 6036 16180
rect 22 16174 3264 16176
rect 22 16170 2336 16174
rect 22 16168 1878 16170
rect 22 16116 38 16168
rect 90 16164 956 16168
rect 90 16116 494 16164
rect 22 16112 494 16116
rect 546 16116 956 16164
rect 1008 16164 1878 16168
rect 1008 16116 1414 16164
rect 546 16112 1414 16116
rect 1466 16118 1878 16164
rect 1930 16122 2336 16170
rect 2388 16122 2806 16174
rect 2858 16124 3264 16174
rect 3316 16124 3728 16176
rect 3780 16124 4190 16176
rect 4242 16124 4652 16176
rect 4704 16124 5112 16176
rect 5164 16124 5576 16176
rect 5628 16128 6036 16176
rect 6088 16178 8918 16180
rect 6088 16176 7426 16178
rect 6088 16174 6960 16176
rect 6088 16128 6502 16174
rect 5628 16124 6502 16128
rect 2858 16122 6502 16124
rect 6554 16124 6960 16174
rect 7012 16126 7426 16176
rect 7478 16126 7888 16178
rect 7940 16126 8348 16178
rect 8400 16172 8918 16178
rect 8400 16126 8810 16172
rect 7012 16124 8810 16126
rect 6554 16122 8810 16124
rect 1930 16120 8810 16122
rect 8862 16120 8918 16172
rect 1930 16118 8918 16120
rect 1466 16112 8918 16118
rect 22 16102 8918 16112
rect -154 235 9114 240
rect -154 231 1198 235
rect -154 229 732 231
rect -154 177 274 229
rect 326 179 732 229
rect 784 183 1198 231
rect 1250 233 2582 235
rect 1250 183 1654 233
rect 784 181 1654 183
rect 1706 231 2582 233
rect 1706 181 2114 231
rect 784 179 2114 181
rect 2166 183 2582 231
rect 2634 233 9114 235
rect 2634 231 3968 233
rect 2634 229 3508 231
rect 2634 183 3046 229
rect 2166 179 3046 183
rect 326 177 3046 179
rect 3098 179 3508 229
rect 3560 181 3968 231
rect 4020 181 4428 233
rect 4480 231 6742 233
rect 4480 229 5352 231
rect 4480 181 4888 229
rect 3560 179 4888 181
rect 3098 177 4888 179
rect 4940 179 5352 229
rect 5404 229 6276 231
rect 5404 179 5814 229
rect 4940 177 5814 179
rect 5866 179 6276 229
rect 6328 181 6742 231
rect 6794 181 7202 233
rect 7254 181 7664 233
rect 7716 231 9114 233
rect 7716 181 8126 231
rect 6328 179 8126 181
rect 8178 179 8586 231
rect 8638 179 9056 231
rect 9108 179 9114 231
rect 5866 177 9114 179
rect -154 166 9114 177
rect -154 162 342 166
use sky130_fd_pr__pfet_01v8_lvt_4QDPGG  sky130_fd_pr__pfet_01v8_lvt_4QDPGG_0
array 19 0 462 0 0 16438
timestamp 1635855079
transform 1 0 178 0 1 8166
box -231 -8219 231 8219
<< labels >>
rlabel metal1 s -216 16116 -216 16116 4 D
port 1 nsew
rlabel metal2 s -132 200 -132 200 4 S
port 2 nsew
rlabel locali s 9120 -6 9120 -6 4 B
port 3 nsew
rlabel metal1 s 504 -162 504 -162 4 G
port 4 nsew
<< end >>
