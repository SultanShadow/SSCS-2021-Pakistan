magic
tech sky130A
magscale 1 2
timestamp 1637060811
<< poly >>
rect 1404 1180 1550 1252
rect 3294 1184 3394 1264
rect 224 980 370 1046
<< locali >>
rect 2045 2435 2079 2466
rect 2045 2363 2079 2401
rect 2045 2291 2079 2329
rect 2045 2219 2079 2257
rect 2045 2147 2079 2185
rect 2045 2083 2079 2113
rect 1304 1861 1824 1862
rect 1303 1750 2216 1861
rect 868 1749 2216 1750
rect 868 1494 1824 1749
rect -614 1337 -590 1371
rect -556 1337 -518 1371
rect -484 1337 -446 1371
rect -412 1337 -374 1371
rect -340 1337 -302 1371
rect -268 1337 -244 1371
rect 868 1292 1287 1494
rect -580 963 6 1224
rect 502 80 622 1034
rect 3438 378 3584 872
rect 876 -12 895 22
rect 929 -12 967 22
rect 1001 -12 1039 22
rect 1073 -12 1111 22
rect 1145 -12 1164 22
rect 761 -89 912 -88
rect 761 -416 914 -89
rect 1346 -753 1972 -385
<< viali >>
rect 2045 2401 2079 2435
rect 2045 2329 2079 2363
rect 2045 2257 2079 2291
rect 2045 2185 2079 2219
rect 2045 2113 2079 2147
rect -590 1337 -556 1371
rect -518 1337 -484 1371
rect -446 1337 -412 1371
rect -374 1337 -340 1371
rect -302 1337 -268 1371
rect 895 -12 929 22
rect 967 -12 1001 22
rect 1039 -12 1073 22
rect 1111 -12 1145 22
<< metal1 >>
rect 2030 2435 4228 2491
rect 2030 2401 2045 2435
rect 2079 2401 4228 2435
rect 2030 2397 4228 2401
rect 821 2300 1054 2375
rect 166 2090 402 2130
rect 166 1674 195 2090
rect -308 1450 195 1674
rect -670 1371 -206 1386
rect -670 1337 -590 1371
rect -556 1337 -518 1371
rect -484 1337 -446 1371
rect -412 1337 -374 1371
rect -340 1337 -302 1371
rect -268 1337 -206 1371
rect -3199 856 -2566 865
rect -3199 812 -2445 856
rect -3199 696 -3135 812
rect -2635 696 -2445 812
rect -3199 651 -2445 696
rect -670 814 -206 1337
rect 166 1014 195 1450
rect 375 1014 402 2090
rect 821 1250 842 2300
rect 816 1224 842 1250
rect 1022 2234 1054 2300
rect 2030 2363 3761 2397
rect 2030 2329 2045 2363
rect 2079 2329 3761 2363
rect 2030 2291 3761 2329
rect 2030 2257 2045 2291
rect 2079 2257 3761 2291
rect 1022 2090 1694 2234
rect 2030 2219 3761 2257
rect 2030 2185 2045 2219
rect 2079 2185 3761 2219
rect 2030 2153 3761 2185
rect 4133 2153 4228 2397
rect 2030 2147 4228 2153
rect 2030 2113 2045 2147
rect 2079 2113 4228 2147
rect 1022 1250 1054 2090
rect 2030 2066 4228 2113
rect 1917 1266 2345 1626
rect 5321 1557 5794 6376
rect 5350 1555 5791 1557
rect 1022 1224 1476 1250
rect 816 1192 1476 1224
rect 1917 1210 3454 1266
rect 1917 1209 2345 1210
rect 166 1000 402 1014
rect 694 1036 764 1054
rect 206 987 371 1000
rect 694 984 707 1036
rect 759 984 764 1036
rect 694 972 764 984
rect 694 920 707 972
rect 759 920 764 972
rect 694 902 764 920
rect 880 1036 948 1062
rect 880 984 891 1036
rect 943 984 948 1036
rect 880 972 948 984
rect 880 920 891 972
rect 943 920 948 972
rect 880 900 948 920
rect 1068 1034 1136 1062
rect 1068 982 1075 1034
rect 1127 982 1136 1034
rect 1068 970 1136 982
rect 1068 918 1075 970
rect 1127 918 1136 970
rect 1068 900 1136 918
rect 1258 1034 1326 1060
rect 1258 982 1269 1034
rect 1321 982 1326 1034
rect 1258 970 1326 982
rect 1258 918 1269 970
rect 1321 918 1326 970
rect 1258 898 1326 918
rect 1458 1034 1526 1054
rect 1458 982 1463 1034
rect 1515 982 1526 1034
rect 1458 970 1526 982
rect 1458 918 1463 970
rect 1515 918 1526 970
rect 1458 892 1526 918
rect 1972 1036 2058 1060
rect 1972 984 1989 1036
rect 2041 984 2058 1036
rect 1972 972 2058 984
rect 1972 920 1989 972
rect 2041 920 2058 972
rect 1972 894 2058 920
rect 2162 1034 2248 1062
rect 2162 982 2177 1034
rect 2229 982 2248 1034
rect 2162 970 2248 982
rect 2162 918 2177 970
rect 2229 918 2248 970
rect 2162 896 2248 918
rect 2356 1036 2442 1062
rect 2356 984 2373 1036
rect 2425 984 2442 1036
rect 2356 972 2442 984
rect 2356 920 2373 972
rect 2425 920 2442 972
rect 2356 896 2442 920
rect 2548 1034 2634 1060
rect 2548 982 2563 1034
rect 2615 982 2634 1034
rect 2548 970 2634 982
rect 2548 918 2563 970
rect 2615 918 2634 970
rect 2548 894 2634 918
rect 2736 1036 2822 1060
rect 2736 984 2751 1036
rect 2803 984 2822 1036
rect 2736 972 2822 984
rect 2736 920 2751 972
rect 2803 920 2822 972
rect 2736 894 2822 920
rect 2930 1040 3016 1062
rect 2930 988 2947 1040
rect 2999 988 3016 1040
rect 2930 976 3016 988
rect 2930 924 2947 976
rect 2999 924 3016 976
rect 2930 896 3016 924
rect 3120 1060 3196 1064
rect 3120 1038 3206 1060
rect 3120 986 3137 1038
rect 3189 986 3206 1038
rect 3120 974 3206 986
rect 3120 922 3137 974
rect 3189 922 3206 974
rect 3120 894 3206 922
rect 3312 1036 3388 1060
rect 3312 984 3321 1036
rect 3373 984 3388 1036
rect 3312 972 3388 984
rect 3312 920 3321 972
rect 3373 920 3388 972
rect 3312 890 3388 920
rect -670 698 -585 814
rect -277 698 -206 814
rect 96 833 156 854
rect 286 846 350 858
rect 148 781 156 833
rect 96 762 156 781
rect 284 833 350 846
rect 336 781 350 833
rect 284 768 350 781
rect 286 758 350 768
rect -3199 -294 -2566 651
rect -670 648 -206 698
rect 184 348 252 360
rect 390 358 732 762
rect 1884 498 1956 508
rect 1884 446 1895 498
rect 1947 446 1956 498
rect 1884 434 1956 446
rect 1884 382 1895 434
rect 1947 382 1956 434
rect 1884 374 1956 382
rect 2078 498 2140 506
rect 2078 446 2083 498
rect 2135 446 2140 498
rect 2078 434 2140 446
rect 2078 382 2083 434
rect 2135 382 2140 434
rect 2078 374 2140 382
rect 2260 504 2322 510
rect 2260 502 2324 504
rect 2260 450 2271 502
rect 2323 450 2324 502
rect 2260 438 2324 450
rect 2260 386 2271 438
rect 2323 386 2324 438
rect 2260 384 2324 386
rect 2458 498 2528 508
rect 2458 446 2467 498
rect 2519 446 2528 498
rect 2458 434 2528 446
rect 2260 378 2322 384
rect 2458 382 2467 434
rect 2519 382 2528 434
rect 2458 376 2528 382
rect 2650 500 2712 508
rect 2650 448 2657 500
rect 2709 448 2712 500
rect 2650 436 2712 448
rect 2650 384 2657 436
rect 2709 384 2712 436
rect 2650 376 2712 384
rect 2846 502 2916 508
rect 2846 450 2853 502
rect 2905 450 2916 502
rect 2846 438 2916 450
rect 2846 386 2853 438
rect 2905 386 2916 438
rect 2846 376 2916 386
rect 3038 498 3108 508
rect 3038 446 3045 498
rect 3097 446 3108 498
rect 3038 434 3108 446
rect 3038 382 3045 434
rect 3097 382 3108 434
rect 3038 376 3108 382
rect 3228 498 3298 506
rect 3228 446 3235 498
rect 3287 446 3298 498
rect 3228 434 3298 446
rect 3228 382 3235 434
rect 3287 382 3298 434
rect 3228 374 3298 382
rect 3416 500 3486 510
rect 3416 448 3427 500
rect 3479 448 3486 500
rect 3416 436 3486 448
rect 3416 384 3427 436
rect 3479 384 3486 436
rect 3416 378 3486 384
rect 184 296 193 348
rect 245 296 252 348
rect 184 284 252 296
rect 184 232 193 284
rect 245 232 252 284
rect 184 222 252 232
rect 364 348 732 358
rect 364 296 372 348
rect 424 344 732 348
rect 424 296 426 344
rect 364 284 426 296
rect 364 232 372 284
rect 424 232 426 284
rect 364 222 426 232
rect 784 303 858 324
rect 784 251 795 303
rect 847 251 858 303
rect 784 230 858 251
rect 972 318 1046 322
rect 972 303 1048 318
rect 972 251 985 303
rect 1037 251 1048 303
rect 972 228 1048 251
rect 1162 303 1236 324
rect 1162 251 1173 303
rect 1225 251 1236 303
rect 1162 230 1236 251
rect 1356 322 1368 326
rect 1544 322 1618 324
rect 1356 305 1434 322
rect 1356 253 1369 305
rect 1421 253 1434 305
rect 1356 236 1434 253
rect 1542 307 1618 322
rect 1542 255 1553 307
rect 1605 255 1618 307
rect 1542 240 1618 255
rect 1360 228 1434 236
rect 1544 230 1618 240
rect 126 120 386 124
rect 126 68 389 120
rect 726 70 1584 128
rect 129 -287 389 68
rect 874 36 1164 42
rect 874 28 897 36
rect 862 22 897 28
rect 862 -12 895 22
rect 862 -16 897 -12
rect 949 -16 961 36
rect 1013 -16 1025 36
rect 1077 -16 1089 36
rect 1141 28 1164 36
rect 1141 22 1210 28
rect 1145 -12 1210 22
rect 1141 -16 1210 -12
rect 862 -42 1210 -16
rect 1263 -288 1432 70
rect 1916 68 3356 126
rect -3196 -673 -2759 -294
rect 3021 -889 3469 -217
<< via1 >>
rect -3135 696 -2635 812
rect 195 1014 375 2090
rect 842 1224 1022 2300
rect 3761 2153 4133 2397
rect 707 984 759 1036
rect 707 920 759 972
rect 891 984 943 1036
rect 891 920 943 972
rect 1075 982 1127 1034
rect 1075 918 1127 970
rect 1269 982 1321 1034
rect 1269 918 1321 970
rect 1463 982 1515 1034
rect 1463 918 1515 970
rect 1989 984 2041 1036
rect 1989 920 2041 972
rect 2177 982 2229 1034
rect 2177 918 2229 970
rect 2373 984 2425 1036
rect 2373 920 2425 972
rect 2563 982 2615 1034
rect 2563 918 2615 970
rect 2751 984 2803 1036
rect 2751 920 2803 972
rect 2947 988 2999 1040
rect 2947 924 2999 976
rect 3137 986 3189 1038
rect 3137 922 3189 974
rect 3321 984 3373 1036
rect 3321 920 3373 972
rect -585 698 -277 814
rect 96 781 148 833
rect 284 781 336 833
rect 1895 446 1947 498
rect 1895 382 1947 434
rect 2083 446 2135 498
rect 2083 382 2135 434
rect 2271 450 2323 502
rect 2271 386 2323 438
rect 2467 446 2519 498
rect 2467 382 2519 434
rect 2657 448 2709 500
rect 2657 384 2709 436
rect 2853 450 2905 502
rect 2853 386 2905 438
rect 3045 446 3097 498
rect 3045 382 3097 434
rect 3235 446 3287 498
rect 3235 382 3287 434
rect 3427 448 3479 500
rect 3427 384 3479 436
rect 193 296 245 348
rect 193 232 245 284
rect 372 296 424 348
rect 372 232 424 284
rect 795 251 847 303
rect 985 251 1037 303
rect 1173 251 1225 303
rect 1369 253 1421 305
rect 1553 255 1605 307
rect 897 22 949 36
rect 897 -12 929 22
rect 929 -12 949 22
rect 897 -16 949 -12
rect 961 22 1013 36
rect 961 -12 967 22
rect 967 -12 1001 22
rect 1001 -12 1013 22
rect 961 -16 1013 -12
rect 1025 22 1077 36
rect 1025 -12 1039 22
rect 1039 -12 1073 22
rect 1073 -12 1077 22
rect 1025 -16 1077 -12
rect 1089 22 1141 36
rect 1089 -12 1111 22
rect 1111 -12 1141 22
rect 1089 -16 1141 -12
<< metal2 >>
rect 120 5768 440 5770
rect -1428 5557 444 5768
rect -1428 4941 -1284 5557
rect 132 4941 444 5557
rect -1428 4822 444 4941
rect 120 2090 440 4822
rect 822 3317 1040 3996
rect 822 2376 864 3317
rect 120 2080 195 2090
rect 166 1014 195 2080
rect 375 2080 440 2090
rect 816 2300 864 2376
rect 1000 2376 1040 3317
rect 1000 2300 1054 2376
rect 375 1014 402 2080
rect 816 1224 842 2300
rect 1022 1224 1054 2300
rect 2775 2071 3380 6301
rect 816 1212 1054 1224
rect 821 1192 1054 1212
rect 2776 1060 3380 2071
rect 3662 2397 4227 2491
rect 3662 2153 3761 2397
rect 4133 2153 4227 2397
rect 166 999 402 1014
rect 694 1040 3388 1060
rect 694 1036 2947 1040
rect 208 994 362 999
rect 694 984 707 1036
rect 759 984 891 1036
rect 943 1034 1989 1036
rect 943 984 1075 1034
rect 694 982 1075 984
rect 1127 982 1269 1034
rect 1321 982 1463 1034
rect 1515 984 1989 1034
rect 2041 1034 2373 1036
rect 2041 984 2177 1034
rect 1515 982 2177 984
rect 2229 984 2373 1034
rect 2425 1034 2751 1036
rect 2425 984 2563 1034
rect 2229 982 2563 984
rect 2615 984 2751 1034
rect 2803 988 2947 1036
rect 2999 1038 3388 1040
rect 2999 988 3137 1038
rect 2803 986 3137 988
rect 3189 1036 3388 1038
rect 3189 986 3321 1036
rect 2803 984 3321 986
rect 3373 984 3388 1036
rect 2615 982 3388 984
rect 694 976 3388 982
rect 694 972 2947 976
rect 694 920 707 972
rect 759 920 891 972
rect 943 970 1989 972
rect 943 920 1075 970
rect 694 918 1075 920
rect 1127 918 1269 970
rect 1321 918 1463 970
rect 1515 920 1989 970
rect 2041 970 2373 972
rect 2041 920 2177 970
rect 1515 918 2177 920
rect 2229 920 2373 970
rect 2425 970 2751 972
rect 2425 920 2563 970
rect 2229 918 2563 920
rect 2615 920 2751 970
rect 2803 924 2947 972
rect 2999 974 3388 976
rect 2999 924 3137 974
rect 2803 922 3137 924
rect 3189 972 3388 974
rect 3189 922 3321 972
rect 2803 920 3321 922
rect 3373 920 3388 972
rect 2615 918 3388 920
rect 694 894 3388 918
rect 1454 892 3388 894
rect 3312 890 3388 892
rect -3178 833 353 860
rect -3178 814 96 833
rect -3178 812 -585 814
rect -3178 696 -3135 812
rect -2635 698 -585 812
rect -277 781 96 814
rect 148 781 284 833
rect 336 781 353 833
rect -277 744 353 781
rect -277 698 2844 744
rect -2635 696 2844 698
rect -3178 644 2844 696
rect 98 508 2844 644
rect 3662 508 4227 2153
rect 98 502 4227 508
rect 98 498 2271 502
rect 98 463 1895 498
rect 1888 446 1895 463
rect 1947 446 2083 498
rect 2135 450 2271 498
rect 2323 500 2853 502
rect 2323 498 2657 500
rect 2323 450 2467 498
rect 2135 446 2467 450
rect 2519 448 2657 498
rect 2709 450 2853 500
rect 2905 500 4227 502
rect 2905 498 3427 500
rect 2905 450 3045 498
rect 2709 448 3045 450
rect 2519 446 3045 448
rect 3097 446 3235 498
rect 3287 448 3427 498
rect 3479 448 4227 500
rect 3287 446 4227 448
rect 1888 438 4227 446
rect 1888 434 2271 438
rect 1888 382 1895 434
rect 1947 382 2083 434
rect 2135 386 2271 434
rect 2323 436 2853 438
rect 2323 434 2657 436
rect 2323 386 2467 434
rect 2135 382 2467 386
rect 2519 384 2657 434
rect 2709 386 2853 436
rect 2905 436 4227 438
rect 2905 434 3427 436
rect 2905 386 3045 434
rect 2709 384 3045 386
rect 2519 382 3045 384
rect 3097 382 3235 434
rect 3287 384 3427 434
rect 3479 384 4227 436
rect 3287 382 4227 384
rect 1888 376 4227 382
rect 182 348 432 362
rect 182 296 193 348
rect 245 296 372 348
rect 424 296 432 348
rect 182 284 432 296
rect 182 232 193 284
rect 245 232 372 284
rect 424 232 432 284
rect 182 220 432 232
rect 786 307 1616 328
rect 786 305 1553 307
rect 786 303 1369 305
rect 786 251 795 303
rect 847 251 985 303
rect 1037 251 1173 303
rect 1225 253 1369 303
rect 1421 255 1553 305
rect 1605 255 1616 307
rect 1421 253 1616 255
rect 1225 251 1616 253
rect 786 228 1616 251
rect 868 36 1176 228
rect 868 -16 897 36
rect 949 -16 961 36
rect 1013 -16 1025 36
rect 1077 -16 1089 36
rect 1141 -16 1176 36
rect 868 -18 1176 -16
<< via2 >>
rect -1284 4941 132 5557
rect 864 2300 1000 3317
rect 864 2221 1000 2300
<< metal3 >>
rect -1440 6972 -194 7084
rect -1440 6028 -1296 6972
rect -352 6028 -194 6972
rect 386 6987 1566 7062
rect 386 6203 524 6987
rect 1388 6203 1566 6987
rect 386 6092 1566 6203
rect -1440 5768 -194 6028
rect -1440 5557 444 5768
rect -1440 5496 -1284 5557
rect -1428 4941 -1284 5496
rect 132 4941 444 5557
rect -1428 4822 444 4941
rect 764 3348 1112 6092
rect 774 3317 1106 3348
rect 774 2221 864 3317
rect 1000 2221 1106 3317
rect 774 2012 1106 2221
<< via3 >>
rect -1296 6028 -352 6972
rect 524 6203 1388 6987
<< metal4 >>
rect -1440 6972 -194 7084
rect -1440 6028 -1296 6972
rect -352 6028 -194 6972
rect 386 6987 1566 7062
rect 386 6203 524 6987
rect 1388 6203 1566 6987
rect 386 6092 1566 6203
rect -1440 5496 -194 6028
rect 774 5496 1098 6092
rect 178 1008 392 2096
rect 838 1212 1026 2313
<< metal5 >>
rect -4557 5180 -1647 6084
rect 3790 5420 4920 6326
use sky130_fd_pr__diode_pd2nw_05v5_WW7YB9  sky130_fd_pr__diode_pd2nw_05v5_WW7YB9_1
timestamp 1637060811
transform 1 0 -434 0 1 1639
box -466 -466 466 466
use sky130_fd_pr__nfet_01v8_lvt_EN8PG3  sky130_fd_pr__nfet_01v8_lvt_EN8PG3_0
timestamp 1637060811
transform 1 0 258 0 1 557
box -301 -600 301 600
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_1
timestamp 1637060811
transform 1 0 -2929 0 1 2664
box -3351 -3101 3373 3101
use sky130_fd_pr__res_high_po_0p35_MGFMH8  sky130_fd_pr__res_high_po_0p35_MGFMH8_1
timestamp 1637060811
transform 0 -1 -1263 1 0 -251
box -191 -2088 191 2088
use sky130_fd_pr__diode_pd2nw_05v5_WW7YB9  sky130_fd_pr__diode_pd2nw_05v5_WW7YB9_0
timestamp 1637060811
transform 1 0 1777 0 1 2260
box -466 -466 466 466
use sky130_fd_pr__nfet_01v8_lvt_USGZYX  sky130_fd_pr__nfet_01v8_lvt_USGZYX_0
timestamp 1637060811
transform 1 0 1151 0 1 658
box -589 -700 589 700
use sky130_fd_pr__pfet_01v8_VCU74W  sky130_fd_pr__pfet_01v8_VCU74W_0
timestamp 1637060811
transform 1 0 2685 0 1 667
box -935 -719 935 719
use sky130_fd_pr__res_high_po_0p35_V3QVRN  sky130_fd_pr__res_high_po_0p35_V3QVRN_0
timestamp 1637060811
transform 0 1 2230 -1 0 -253
box -191 -1388 191 1388
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1637060811
transform -1 0 4150 0 -1 2663
box -3351 -3101 3373 3101
use sky130_fd_pr__res_high_po_0p35_MGFMH8  sky130_fd_pr__res_high_po_0p35_MGFMH8_0
timestamp 1637060811
transform 0 -1 3847 1 0 1590
box -191 -2088 191 2088
<< labels >>
rlabel metal1 s 3272 -840 3272 -840 4 VCASC10
port 1 nsew
rlabel metal1 s 5535 6329 5535 6329 4 VDD9
port 2 nsew
rlabel metal2 s 2982 6299 2982 6299 4 Vo2
port 3 nsew
rlabel metal5 s -3234 6049 -3234 6049 4 Vo1p
port 4 nsew
rlabel metal5 s 4301 6316 4301 6316 4 Vo1n
port 5 nsew
rlabel metal1 s -2964 -669 -2964 -669 4 VDD
port 6 nsew
rlabel locali s 1598 -750 1598 -750 4 VSS
port 7 nsew
<< end >>
