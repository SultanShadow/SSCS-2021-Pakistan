magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< pwell >>
rect -255 956 2546 1142
rect -255 -2 -89 956
rect 2380 -2 2546 956
rect -255 -854 2546 -2
rect -255 -1026 -89 -854
rect 2380 -1026 2546 -854
rect -255 -1212 2546 -1026
<< nmoslvt >>
rect 58 -828 88 -28
rect 146 -828 176 -28
rect 234 -828 264 -28
rect 322 -828 352 -28
rect 410 -828 440 -28
rect 498 -828 528 -28
rect 586 -828 616 -28
rect 674 -828 704 -28
rect 762 -828 792 -28
rect 850 -828 880 -28
rect 938 -828 968 -28
rect 1026 -828 1056 -28
rect 1114 -828 1144 -28
rect 1202 -828 1232 -28
rect 1290 -828 1320 -28
rect 1378 -828 1408 -28
rect 1466 -828 1496 -28
rect 1554 -828 1584 -28
rect 1642 -828 1672 -28
rect 1730 -828 1760 -28
rect 1818 -828 1848 -28
rect 1906 -828 1936 -28
rect 1994 -828 2024 -28
rect 2082 -828 2112 -28
rect 2170 -828 2200 -28
<< ndiff >>
rect 0 -71 58 -28
rect 0 -105 12 -71
rect 46 -105 58 -71
rect 0 -139 58 -105
rect 0 -173 12 -139
rect 46 -173 58 -139
rect 0 -207 58 -173
rect 0 -241 12 -207
rect 46 -241 58 -207
rect 0 -275 58 -241
rect 0 -309 12 -275
rect 46 -309 58 -275
rect 0 -343 58 -309
rect 0 -377 12 -343
rect 46 -377 58 -343
rect 0 -411 58 -377
rect 0 -445 12 -411
rect 46 -445 58 -411
rect 0 -479 58 -445
rect 0 -513 12 -479
rect 46 -513 58 -479
rect 0 -547 58 -513
rect 0 -581 12 -547
rect 46 -581 58 -547
rect 0 -615 58 -581
rect 0 -649 12 -615
rect 46 -649 58 -615
rect 0 -683 58 -649
rect 0 -717 12 -683
rect 46 -717 58 -683
rect 0 -751 58 -717
rect 0 -785 12 -751
rect 46 -785 58 -751
rect 0 -828 58 -785
rect 88 -71 146 -28
rect 88 -105 100 -71
rect 134 -105 146 -71
rect 88 -139 146 -105
rect 88 -173 100 -139
rect 134 -173 146 -139
rect 88 -207 146 -173
rect 88 -241 100 -207
rect 134 -241 146 -207
rect 88 -275 146 -241
rect 88 -309 100 -275
rect 134 -309 146 -275
rect 88 -343 146 -309
rect 88 -377 100 -343
rect 134 -377 146 -343
rect 88 -411 146 -377
rect 88 -445 100 -411
rect 134 -445 146 -411
rect 88 -479 146 -445
rect 88 -513 100 -479
rect 134 -513 146 -479
rect 88 -547 146 -513
rect 88 -581 100 -547
rect 134 -581 146 -547
rect 88 -615 146 -581
rect 88 -649 100 -615
rect 134 -649 146 -615
rect 88 -683 146 -649
rect 88 -717 100 -683
rect 134 -717 146 -683
rect 88 -751 146 -717
rect 88 -785 100 -751
rect 134 -785 146 -751
rect 88 -828 146 -785
rect 176 -71 234 -28
rect 176 -105 188 -71
rect 222 -105 234 -71
rect 176 -139 234 -105
rect 176 -173 188 -139
rect 222 -173 234 -139
rect 176 -207 234 -173
rect 176 -241 188 -207
rect 222 -241 234 -207
rect 176 -275 234 -241
rect 176 -309 188 -275
rect 222 -309 234 -275
rect 176 -343 234 -309
rect 176 -377 188 -343
rect 222 -377 234 -343
rect 176 -411 234 -377
rect 176 -445 188 -411
rect 222 -445 234 -411
rect 176 -479 234 -445
rect 176 -513 188 -479
rect 222 -513 234 -479
rect 176 -547 234 -513
rect 176 -581 188 -547
rect 222 -581 234 -547
rect 176 -615 234 -581
rect 176 -649 188 -615
rect 222 -649 234 -615
rect 176 -683 234 -649
rect 176 -717 188 -683
rect 222 -717 234 -683
rect 176 -751 234 -717
rect 176 -785 188 -751
rect 222 -785 234 -751
rect 176 -828 234 -785
rect 264 -71 322 -28
rect 264 -105 276 -71
rect 310 -105 322 -71
rect 264 -139 322 -105
rect 264 -173 276 -139
rect 310 -173 322 -139
rect 264 -207 322 -173
rect 264 -241 276 -207
rect 310 -241 322 -207
rect 264 -275 322 -241
rect 264 -309 276 -275
rect 310 -309 322 -275
rect 264 -343 322 -309
rect 264 -377 276 -343
rect 310 -377 322 -343
rect 264 -411 322 -377
rect 264 -445 276 -411
rect 310 -445 322 -411
rect 264 -479 322 -445
rect 264 -513 276 -479
rect 310 -513 322 -479
rect 264 -547 322 -513
rect 264 -581 276 -547
rect 310 -581 322 -547
rect 264 -615 322 -581
rect 264 -649 276 -615
rect 310 -649 322 -615
rect 264 -683 322 -649
rect 264 -717 276 -683
rect 310 -717 322 -683
rect 264 -751 322 -717
rect 264 -785 276 -751
rect 310 -785 322 -751
rect 264 -828 322 -785
rect 352 -71 410 -28
rect 352 -105 364 -71
rect 398 -105 410 -71
rect 352 -139 410 -105
rect 352 -173 364 -139
rect 398 -173 410 -139
rect 352 -207 410 -173
rect 352 -241 364 -207
rect 398 -241 410 -207
rect 352 -275 410 -241
rect 352 -309 364 -275
rect 398 -309 410 -275
rect 352 -343 410 -309
rect 352 -377 364 -343
rect 398 -377 410 -343
rect 352 -411 410 -377
rect 352 -445 364 -411
rect 398 -445 410 -411
rect 352 -479 410 -445
rect 352 -513 364 -479
rect 398 -513 410 -479
rect 352 -547 410 -513
rect 352 -581 364 -547
rect 398 -581 410 -547
rect 352 -615 410 -581
rect 352 -649 364 -615
rect 398 -649 410 -615
rect 352 -683 410 -649
rect 352 -717 364 -683
rect 398 -717 410 -683
rect 352 -751 410 -717
rect 352 -785 364 -751
rect 398 -785 410 -751
rect 352 -828 410 -785
rect 440 -71 498 -28
rect 440 -105 452 -71
rect 486 -105 498 -71
rect 440 -139 498 -105
rect 440 -173 452 -139
rect 486 -173 498 -139
rect 440 -207 498 -173
rect 440 -241 452 -207
rect 486 -241 498 -207
rect 440 -275 498 -241
rect 440 -309 452 -275
rect 486 -309 498 -275
rect 440 -343 498 -309
rect 440 -377 452 -343
rect 486 -377 498 -343
rect 440 -411 498 -377
rect 440 -445 452 -411
rect 486 -445 498 -411
rect 440 -479 498 -445
rect 440 -513 452 -479
rect 486 -513 498 -479
rect 440 -547 498 -513
rect 440 -581 452 -547
rect 486 -581 498 -547
rect 440 -615 498 -581
rect 440 -649 452 -615
rect 486 -649 498 -615
rect 440 -683 498 -649
rect 440 -717 452 -683
rect 486 -717 498 -683
rect 440 -751 498 -717
rect 440 -785 452 -751
rect 486 -785 498 -751
rect 440 -828 498 -785
rect 528 -71 586 -28
rect 528 -105 540 -71
rect 574 -105 586 -71
rect 528 -139 586 -105
rect 528 -173 540 -139
rect 574 -173 586 -139
rect 528 -207 586 -173
rect 528 -241 540 -207
rect 574 -241 586 -207
rect 528 -275 586 -241
rect 528 -309 540 -275
rect 574 -309 586 -275
rect 528 -343 586 -309
rect 528 -377 540 -343
rect 574 -377 586 -343
rect 528 -411 586 -377
rect 528 -445 540 -411
rect 574 -445 586 -411
rect 528 -479 586 -445
rect 528 -513 540 -479
rect 574 -513 586 -479
rect 528 -547 586 -513
rect 528 -581 540 -547
rect 574 -581 586 -547
rect 528 -615 586 -581
rect 528 -649 540 -615
rect 574 -649 586 -615
rect 528 -683 586 -649
rect 528 -717 540 -683
rect 574 -717 586 -683
rect 528 -751 586 -717
rect 528 -785 540 -751
rect 574 -785 586 -751
rect 528 -828 586 -785
rect 616 -71 674 -28
rect 616 -105 628 -71
rect 662 -105 674 -71
rect 616 -139 674 -105
rect 616 -173 628 -139
rect 662 -173 674 -139
rect 616 -207 674 -173
rect 616 -241 628 -207
rect 662 -241 674 -207
rect 616 -275 674 -241
rect 616 -309 628 -275
rect 662 -309 674 -275
rect 616 -343 674 -309
rect 616 -377 628 -343
rect 662 -377 674 -343
rect 616 -411 674 -377
rect 616 -445 628 -411
rect 662 -445 674 -411
rect 616 -479 674 -445
rect 616 -513 628 -479
rect 662 -513 674 -479
rect 616 -547 674 -513
rect 616 -581 628 -547
rect 662 -581 674 -547
rect 616 -615 674 -581
rect 616 -649 628 -615
rect 662 -649 674 -615
rect 616 -683 674 -649
rect 616 -717 628 -683
rect 662 -717 674 -683
rect 616 -751 674 -717
rect 616 -785 628 -751
rect 662 -785 674 -751
rect 616 -828 674 -785
rect 704 -71 762 -28
rect 704 -105 716 -71
rect 750 -105 762 -71
rect 704 -139 762 -105
rect 704 -173 716 -139
rect 750 -173 762 -139
rect 704 -207 762 -173
rect 704 -241 716 -207
rect 750 -241 762 -207
rect 704 -275 762 -241
rect 704 -309 716 -275
rect 750 -309 762 -275
rect 704 -343 762 -309
rect 704 -377 716 -343
rect 750 -377 762 -343
rect 704 -411 762 -377
rect 704 -445 716 -411
rect 750 -445 762 -411
rect 704 -479 762 -445
rect 704 -513 716 -479
rect 750 -513 762 -479
rect 704 -547 762 -513
rect 704 -581 716 -547
rect 750 -581 762 -547
rect 704 -615 762 -581
rect 704 -649 716 -615
rect 750 -649 762 -615
rect 704 -683 762 -649
rect 704 -717 716 -683
rect 750 -717 762 -683
rect 704 -751 762 -717
rect 704 -785 716 -751
rect 750 -785 762 -751
rect 704 -828 762 -785
rect 792 -71 850 -28
rect 792 -105 804 -71
rect 838 -105 850 -71
rect 792 -139 850 -105
rect 792 -173 804 -139
rect 838 -173 850 -139
rect 792 -207 850 -173
rect 792 -241 804 -207
rect 838 -241 850 -207
rect 792 -275 850 -241
rect 792 -309 804 -275
rect 838 -309 850 -275
rect 792 -343 850 -309
rect 792 -377 804 -343
rect 838 -377 850 -343
rect 792 -411 850 -377
rect 792 -445 804 -411
rect 838 -445 850 -411
rect 792 -479 850 -445
rect 792 -513 804 -479
rect 838 -513 850 -479
rect 792 -547 850 -513
rect 792 -581 804 -547
rect 838 -581 850 -547
rect 792 -615 850 -581
rect 792 -649 804 -615
rect 838 -649 850 -615
rect 792 -683 850 -649
rect 792 -717 804 -683
rect 838 -717 850 -683
rect 792 -751 850 -717
rect 792 -785 804 -751
rect 838 -785 850 -751
rect 792 -828 850 -785
rect 880 -71 938 -28
rect 880 -105 892 -71
rect 926 -105 938 -71
rect 880 -139 938 -105
rect 880 -173 892 -139
rect 926 -173 938 -139
rect 880 -207 938 -173
rect 880 -241 892 -207
rect 926 -241 938 -207
rect 880 -275 938 -241
rect 880 -309 892 -275
rect 926 -309 938 -275
rect 880 -343 938 -309
rect 880 -377 892 -343
rect 926 -377 938 -343
rect 880 -411 938 -377
rect 880 -445 892 -411
rect 926 -445 938 -411
rect 880 -479 938 -445
rect 880 -513 892 -479
rect 926 -513 938 -479
rect 880 -547 938 -513
rect 880 -581 892 -547
rect 926 -581 938 -547
rect 880 -615 938 -581
rect 880 -649 892 -615
rect 926 -649 938 -615
rect 880 -683 938 -649
rect 880 -717 892 -683
rect 926 -717 938 -683
rect 880 -751 938 -717
rect 880 -785 892 -751
rect 926 -785 938 -751
rect 880 -828 938 -785
rect 968 -71 1026 -28
rect 968 -105 980 -71
rect 1014 -105 1026 -71
rect 968 -139 1026 -105
rect 968 -173 980 -139
rect 1014 -173 1026 -139
rect 968 -207 1026 -173
rect 968 -241 980 -207
rect 1014 -241 1026 -207
rect 968 -275 1026 -241
rect 968 -309 980 -275
rect 1014 -309 1026 -275
rect 968 -343 1026 -309
rect 968 -377 980 -343
rect 1014 -377 1026 -343
rect 968 -411 1026 -377
rect 968 -445 980 -411
rect 1014 -445 1026 -411
rect 968 -479 1026 -445
rect 968 -513 980 -479
rect 1014 -513 1026 -479
rect 968 -547 1026 -513
rect 968 -581 980 -547
rect 1014 -581 1026 -547
rect 968 -615 1026 -581
rect 968 -649 980 -615
rect 1014 -649 1026 -615
rect 968 -683 1026 -649
rect 968 -717 980 -683
rect 1014 -717 1026 -683
rect 968 -751 1026 -717
rect 968 -785 980 -751
rect 1014 -785 1026 -751
rect 968 -828 1026 -785
rect 1056 -71 1114 -28
rect 1056 -105 1068 -71
rect 1102 -105 1114 -71
rect 1056 -139 1114 -105
rect 1056 -173 1068 -139
rect 1102 -173 1114 -139
rect 1056 -207 1114 -173
rect 1056 -241 1068 -207
rect 1102 -241 1114 -207
rect 1056 -275 1114 -241
rect 1056 -309 1068 -275
rect 1102 -309 1114 -275
rect 1056 -343 1114 -309
rect 1056 -377 1068 -343
rect 1102 -377 1114 -343
rect 1056 -411 1114 -377
rect 1056 -445 1068 -411
rect 1102 -445 1114 -411
rect 1056 -479 1114 -445
rect 1056 -513 1068 -479
rect 1102 -513 1114 -479
rect 1056 -547 1114 -513
rect 1056 -581 1068 -547
rect 1102 -581 1114 -547
rect 1056 -615 1114 -581
rect 1056 -649 1068 -615
rect 1102 -649 1114 -615
rect 1056 -683 1114 -649
rect 1056 -717 1068 -683
rect 1102 -717 1114 -683
rect 1056 -751 1114 -717
rect 1056 -785 1068 -751
rect 1102 -785 1114 -751
rect 1056 -828 1114 -785
rect 1144 -71 1202 -28
rect 1144 -105 1156 -71
rect 1190 -105 1202 -71
rect 1144 -139 1202 -105
rect 1144 -173 1156 -139
rect 1190 -173 1202 -139
rect 1144 -207 1202 -173
rect 1144 -241 1156 -207
rect 1190 -241 1202 -207
rect 1144 -275 1202 -241
rect 1144 -309 1156 -275
rect 1190 -309 1202 -275
rect 1144 -343 1202 -309
rect 1144 -377 1156 -343
rect 1190 -377 1202 -343
rect 1144 -411 1202 -377
rect 1144 -445 1156 -411
rect 1190 -445 1202 -411
rect 1144 -479 1202 -445
rect 1144 -513 1156 -479
rect 1190 -513 1202 -479
rect 1144 -547 1202 -513
rect 1144 -581 1156 -547
rect 1190 -581 1202 -547
rect 1144 -615 1202 -581
rect 1144 -649 1156 -615
rect 1190 -649 1202 -615
rect 1144 -683 1202 -649
rect 1144 -717 1156 -683
rect 1190 -717 1202 -683
rect 1144 -751 1202 -717
rect 1144 -785 1156 -751
rect 1190 -785 1202 -751
rect 1144 -828 1202 -785
rect 1232 -71 1290 -28
rect 1232 -105 1244 -71
rect 1278 -105 1290 -71
rect 1232 -139 1290 -105
rect 1232 -173 1244 -139
rect 1278 -173 1290 -139
rect 1232 -207 1290 -173
rect 1232 -241 1244 -207
rect 1278 -241 1290 -207
rect 1232 -275 1290 -241
rect 1232 -309 1244 -275
rect 1278 -309 1290 -275
rect 1232 -343 1290 -309
rect 1232 -377 1244 -343
rect 1278 -377 1290 -343
rect 1232 -411 1290 -377
rect 1232 -445 1244 -411
rect 1278 -445 1290 -411
rect 1232 -479 1290 -445
rect 1232 -513 1244 -479
rect 1278 -513 1290 -479
rect 1232 -547 1290 -513
rect 1232 -581 1244 -547
rect 1278 -581 1290 -547
rect 1232 -615 1290 -581
rect 1232 -649 1244 -615
rect 1278 -649 1290 -615
rect 1232 -683 1290 -649
rect 1232 -717 1244 -683
rect 1278 -717 1290 -683
rect 1232 -751 1290 -717
rect 1232 -785 1244 -751
rect 1278 -785 1290 -751
rect 1232 -828 1290 -785
rect 1320 -71 1378 -28
rect 1320 -105 1332 -71
rect 1366 -105 1378 -71
rect 1320 -139 1378 -105
rect 1320 -173 1332 -139
rect 1366 -173 1378 -139
rect 1320 -207 1378 -173
rect 1320 -241 1332 -207
rect 1366 -241 1378 -207
rect 1320 -275 1378 -241
rect 1320 -309 1332 -275
rect 1366 -309 1378 -275
rect 1320 -343 1378 -309
rect 1320 -377 1332 -343
rect 1366 -377 1378 -343
rect 1320 -411 1378 -377
rect 1320 -445 1332 -411
rect 1366 -445 1378 -411
rect 1320 -479 1378 -445
rect 1320 -513 1332 -479
rect 1366 -513 1378 -479
rect 1320 -547 1378 -513
rect 1320 -581 1332 -547
rect 1366 -581 1378 -547
rect 1320 -615 1378 -581
rect 1320 -649 1332 -615
rect 1366 -649 1378 -615
rect 1320 -683 1378 -649
rect 1320 -717 1332 -683
rect 1366 -717 1378 -683
rect 1320 -751 1378 -717
rect 1320 -785 1332 -751
rect 1366 -785 1378 -751
rect 1320 -828 1378 -785
rect 1408 -71 1466 -28
rect 1408 -105 1420 -71
rect 1454 -105 1466 -71
rect 1408 -139 1466 -105
rect 1408 -173 1420 -139
rect 1454 -173 1466 -139
rect 1408 -207 1466 -173
rect 1408 -241 1420 -207
rect 1454 -241 1466 -207
rect 1408 -275 1466 -241
rect 1408 -309 1420 -275
rect 1454 -309 1466 -275
rect 1408 -343 1466 -309
rect 1408 -377 1420 -343
rect 1454 -377 1466 -343
rect 1408 -411 1466 -377
rect 1408 -445 1420 -411
rect 1454 -445 1466 -411
rect 1408 -479 1466 -445
rect 1408 -513 1420 -479
rect 1454 -513 1466 -479
rect 1408 -547 1466 -513
rect 1408 -581 1420 -547
rect 1454 -581 1466 -547
rect 1408 -615 1466 -581
rect 1408 -649 1420 -615
rect 1454 -649 1466 -615
rect 1408 -683 1466 -649
rect 1408 -717 1420 -683
rect 1454 -717 1466 -683
rect 1408 -751 1466 -717
rect 1408 -785 1420 -751
rect 1454 -785 1466 -751
rect 1408 -828 1466 -785
rect 1496 -71 1554 -28
rect 1496 -105 1508 -71
rect 1542 -105 1554 -71
rect 1496 -139 1554 -105
rect 1496 -173 1508 -139
rect 1542 -173 1554 -139
rect 1496 -207 1554 -173
rect 1496 -241 1508 -207
rect 1542 -241 1554 -207
rect 1496 -275 1554 -241
rect 1496 -309 1508 -275
rect 1542 -309 1554 -275
rect 1496 -343 1554 -309
rect 1496 -377 1508 -343
rect 1542 -377 1554 -343
rect 1496 -411 1554 -377
rect 1496 -445 1508 -411
rect 1542 -445 1554 -411
rect 1496 -479 1554 -445
rect 1496 -513 1508 -479
rect 1542 -513 1554 -479
rect 1496 -547 1554 -513
rect 1496 -581 1508 -547
rect 1542 -581 1554 -547
rect 1496 -615 1554 -581
rect 1496 -649 1508 -615
rect 1542 -649 1554 -615
rect 1496 -683 1554 -649
rect 1496 -717 1508 -683
rect 1542 -717 1554 -683
rect 1496 -751 1554 -717
rect 1496 -785 1508 -751
rect 1542 -785 1554 -751
rect 1496 -828 1554 -785
rect 1584 -71 1642 -28
rect 1584 -105 1596 -71
rect 1630 -105 1642 -71
rect 1584 -139 1642 -105
rect 1584 -173 1596 -139
rect 1630 -173 1642 -139
rect 1584 -207 1642 -173
rect 1584 -241 1596 -207
rect 1630 -241 1642 -207
rect 1584 -275 1642 -241
rect 1584 -309 1596 -275
rect 1630 -309 1642 -275
rect 1584 -343 1642 -309
rect 1584 -377 1596 -343
rect 1630 -377 1642 -343
rect 1584 -411 1642 -377
rect 1584 -445 1596 -411
rect 1630 -445 1642 -411
rect 1584 -479 1642 -445
rect 1584 -513 1596 -479
rect 1630 -513 1642 -479
rect 1584 -547 1642 -513
rect 1584 -581 1596 -547
rect 1630 -581 1642 -547
rect 1584 -615 1642 -581
rect 1584 -649 1596 -615
rect 1630 -649 1642 -615
rect 1584 -683 1642 -649
rect 1584 -717 1596 -683
rect 1630 -717 1642 -683
rect 1584 -751 1642 -717
rect 1584 -785 1596 -751
rect 1630 -785 1642 -751
rect 1584 -828 1642 -785
rect 1672 -71 1730 -28
rect 1672 -105 1684 -71
rect 1718 -105 1730 -71
rect 1672 -139 1730 -105
rect 1672 -173 1684 -139
rect 1718 -173 1730 -139
rect 1672 -207 1730 -173
rect 1672 -241 1684 -207
rect 1718 -241 1730 -207
rect 1672 -275 1730 -241
rect 1672 -309 1684 -275
rect 1718 -309 1730 -275
rect 1672 -343 1730 -309
rect 1672 -377 1684 -343
rect 1718 -377 1730 -343
rect 1672 -411 1730 -377
rect 1672 -445 1684 -411
rect 1718 -445 1730 -411
rect 1672 -479 1730 -445
rect 1672 -513 1684 -479
rect 1718 -513 1730 -479
rect 1672 -547 1730 -513
rect 1672 -581 1684 -547
rect 1718 -581 1730 -547
rect 1672 -615 1730 -581
rect 1672 -649 1684 -615
rect 1718 -649 1730 -615
rect 1672 -683 1730 -649
rect 1672 -717 1684 -683
rect 1718 -717 1730 -683
rect 1672 -751 1730 -717
rect 1672 -785 1684 -751
rect 1718 -785 1730 -751
rect 1672 -828 1730 -785
rect 1760 -71 1818 -28
rect 1760 -105 1772 -71
rect 1806 -105 1818 -71
rect 1760 -139 1818 -105
rect 1760 -173 1772 -139
rect 1806 -173 1818 -139
rect 1760 -207 1818 -173
rect 1760 -241 1772 -207
rect 1806 -241 1818 -207
rect 1760 -275 1818 -241
rect 1760 -309 1772 -275
rect 1806 -309 1818 -275
rect 1760 -343 1818 -309
rect 1760 -377 1772 -343
rect 1806 -377 1818 -343
rect 1760 -411 1818 -377
rect 1760 -445 1772 -411
rect 1806 -445 1818 -411
rect 1760 -479 1818 -445
rect 1760 -513 1772 -479
rect 1806 -513 1818 -479
rect 1760 -547 1818 -513
rect 1760 -581 1772 -547
rect 1806 -581 1818 -547
rect 1760 -615 1818 -581
rect 1760 -649 1772 -615
rect 1806 -649 1818 -615
rect 1760 -683 1818 -649
rect 1760 -717 1772 -683
rect 1806 -717 1818 -683
rect 1760 -751 1818 -717
rect 1760 -785 1772 -751
rect 1806 -785 1818 -751
rect 1760 -828 1818 -785
rect 1848 -71 1906 -28
rect 1848 -105 1860 -71
rect 1894 -105 1906 -71
rect 1848 -139 1906 -105
rect 1848 -173 1860 -139
rect 1894 -173 1906 -139
rect 1848 -207 1906 -173
rect 1848 -241 1860 -207
rect 1894 -241 1906 -207
rect 1848 -275 1906 -241
rect 1848 -309 1860 -275
rect 1894 -309 1906 -275
rect 1848 -343 1906 -309
rect 1848 -377 1860 -343
rect 1894 -377 1906 -343
rect 1848 -411 1906 -377
rect 1848 -445 1860 -411
rect 1894 -445 1906 -411
rect 1848 -479 1906 -445
rect 1848 -513 1860 -479
rect 1894 -513 1906 -479
rect 1848 -547 1906 -513
rect 1848 -581 1860 -547
rect 1894 -581 1906 -547
rect 1848 -615 1906 -581
rect 1848 -649 1860 -615
rect 1894 -649 1906 -615
rect 1848 -683 1906 -649
rect 1848 -717 1860 -683
rect 1894 -717 1906 -683
rect 1848 -751 1906 -717
rect 1848 -785 1860 -751
rect 1894 -785 1906 -751
rect 1848 -828 1906 -785
rect 1936 -71 1994 -28
rect 1936 -105 1948 -71
rect 1982 -105 1994 -71
rect 1936 -139 1994 -105
rect 1936 -173 1948 -139
rect 1982 -173 1994 -139
rect 1936 -207 1994 -173
rect 1936 -241 1948 -207
rect 1982 -241 1994 -207
rect 1936 -275 1994 -241
rect 1936 -309 1948 -275
rect 1982 -309 1994 -275
rect 1936 -343 1994 -309
rect 1936 -377 1948 -343
rect 1982 -377 1994 -343
rect 1936 -411 1994 -377
rect 1936 -445 1948 -411
rect 1982 -445 1994 -411
rect 1936 -479 1994 -445
rect 1936 -513 1948 -479
rect 1982 -513 1994 -479
rect 1936 -547 1994 -513
rect 1936 -581 1948 -547
rect 1982 -581 1994 -547
rect 1936 -615 1994 -581
rect 1936 -649 1948 -615
rect 1982 -649 1994 -615
rect 1936 -683 1994 -649
rect 1936 -717 1948 -683
rect 1982 -717 1994 -683
rect 1936 -751 1994 -717
rect 1936 -785 1948 -751
rect 1982 -785 1994 -751
rect 1936 -828 1994 -785
rect 2024 -71 2082 -28
rect 2024 -105 2036 -71
rect 2070 -105 2082 -71
rect 2024 -139 2082 -105
rect 2024 -173 2036 -139
rect 2070 -173 2082 -139
rect 2024 -207 2082 -173
rect 2024 -241 2036 -207
rect 2070 -241 2082 -207
rect 2024 -275 2082 -241
rect 2024 -309 2036 -275
rect 2070 -309 2082 -275
rect 2024 -343 2082 -309
rect 2024 -377 2036 -343
rect 2070 -377 2082 -343
rect 2024 -411 2082 -377
rect 2024 -445 2036 -411
rect 2070 -445 2082 -411
rect 2024 -479 2082 -445
rect 2024 -513 2036 -479
rect 2070 -513 2082 -479
rect 2024 -547 2082 -513
rect 2024 -581 2036 -547
rect 2070 -581 2082 -547
rect 2024 -615 2082 -581
rect 2024 -649 2036 -615
rect 2070 -649 2082 -615
rect 2024 -683 2082 -649
rect 2024 -717 2036 -683
rect 2070 -717 2082 -683
rect 2024 -751 2082 -717
rect 2024 -785 2036 -751
rect 2070 -785 2082 -751
rect 2024 -828 2082 -785
rect 2112 -71 2170 -28
rect 2112 -105 2124 -71
rect 2158 -105 2170 -71
rect 2112 -139 2170 -105
rect 2112 -173 2124 -139
rect 2158 -173 2170 -139
rect 2112 -207 2170 -173
rect 2112 -241 2124 -207
rect 2158 -241 2170 -207
rect 2112 -275 2170 -241
rect 2112 -309 2124 -275
rect 2158 -309 2170 -275
rect 2112 -343 2170 -309
rect 2112 -377 2124 -343
rect 2158 -377 2170 -343
rect 2112 -411 2170 -377
rect 2112 -445 2124 -411
rect 2158 -445 2170 -411
rect 2112 -479 2170 -445
rect 2112 -513 2124 -479
rect 2158 -513 2170 -479
rect 2112 -547 2170 -513
rect 2112 -581 2124 -547
rect 2158 -581 2170 -547
rect 2112 -615 2170 -581
rect 2112 -649 2124 -615
rect 2158 -649 2170 -615
rect 2112 -683 2170 -649
rect 2112 -717 2124 -683
rect 2158 -717 2170 -683
rect 2112 -751 2170 -717
rect 2112 -785 2124 -751
rect 2158 -785 2170 -751
rect 2112 -828 2170 -785
rect 2200 -71 2257 -28
rect 2200 -105 2212 -71
rect 2246 -105 2257 -71
rect 2200 -139 2257 -105
rect 2200 -173 2212 -139
rect 2246 -173 2257 -139
rect 2200 -207 2257 -173
rect 2200 -241 2212 -207
rect 2246 -241 2257 -207
rect 2200 -275 2257 -241
rect 2200 -309 2212 -275
rect 2246 -309 2257 -275
rect 2200 -343 2257 -309
rect 2200 -377 2212 -343
rect 2246 -377 2257 -343
rect 2200 -411 2257 -377
rect 2200 -445 2212 -411
rect 2246 -445 2257 -411
rect 2200 -479 2257 -445
rect 2200 -513 2212 -479
rect 2246 -513 2257 -479
rect 2200 -547 2257 -513
rect 2200 -581 2212 -547
rect 2246 -581 2257 -547
rect 2200 -615 2257 -581
rect 2200 -649 2212 -615
rect 2246 -649 2257 -615
rect 2200 -683 2257 -649
rect 2200 -717 2212 -683
rect 2246 -717 2257 -683
rect 2200 -751 2257 -717
rect 2200 -785 2212 -751
rect 2246 -785 2257 -751
rect 2200 -828 2257 -785
<< ndiffc >>
rect 12 -105 46 -71
rect 12 -173 46 -139
rect 12 -241 46 -207
rect 12 -309 46 -275
rect 12 -377 46 -343
rect 12 -445 46 -411
rect 12 -513 46 -479
rect 12 -581 46 -547
rect 12 -649 46 -615
rect 12 -717 46 -683
rect 12 -785 46 -751
rect 100 -105 134 -71
rect 100 -173 134 -139
rect 100 -241 134 -207
rect 100 -309 134 -275
rect 100 -377 134 -343
rect 100 -445 134 -411
rect 100 -513 134 -479
rect 100 -581 134 -547
rect 100 -649 134 -615
rect 100 -717 134 -683
rect 100 -785 134 -751
rect 188 -105 222 -71
rect 188 -173 222 -139
rect 188 -241 222 -207
rect 188 -309 222 -275
rect 188 -377 222 -343
rect 188 -445 222 -411
rect 188 -513 222 -479
rect 188 -581 222 -547
rect 188 -649 222 -615
rect 188 -717 222 -683
rect 188 -785 222 -751
rect 276 -105 310 -71
rect 276 -173 310 -139
rect 276 -241 310 -207
rect 276 -309 310 -275
rect 276 -377 310 -343
rect 276 -445 310 -411
rect 276 -513 310 -479
rect 276 -581 310 -547
rect 276 -649 310 -615
rect 276 -717 310 -683
rect 276 -785 310 -751
rect 364 -105 398 -71
rect 364 -173 398 -139
rect 364 -241 398 -207
rect 364 -309 398 -275
rect 364 -377 398 -343
rect 364 -445 398 -411
rect 364 -513 398 -479
rect 364 -581 398 -547
rect 364 -649 398 -615
rect 364 -717 398 -683
rect 364 -785 398 -751
rect 452 -105 486 -71
rect 452 -173 486 -139
rect 452 -241 486 -207
rect 452 -309 486 -275
rect 452 -377 486 -343
rect 452 -445 486 -411
rect 452 -513 486 -479
rect 452 -581 486 -547
rect 452 -649 486 -615
rect 452 -717 486 -683
rect 452 -785 486 -751
rect 540 -105 574 -71
rect 540 -173 574 -139
rect 540 -241 574 -207
rect 540 -309 574 -275
rect 540 -377 574 -343
rect 540 -445 574 -411
rect 540 -513 574 -479
rect 540 -581 574 -547
rect 540 -649 574 -615
rect 540 -717 574 -683
rect 540 -785 574 -751
rect 628 -105 662 -71
rect 628 -173 662 -139
rect 628 -241 662 -207
rect 628 -309 662 -275
rect 628 -377 662 -343
rect 628 -445 662 -411
rect 628 -513 662 -479
rect 628 -581 662 -547
rect 628 -649 662 -615
rect 628 -717 662 -683
rect 628 -785 662 -751
rect 716 -105 750 -71
rect 716 -173 750 -139
rect 716 -241 750 -207
rect 716 -309 750 -275
rect 716 -377 750 -343
rect 716 -445 750 -411
rect 716 -513 750 -479
rect 716 -581 750 -547
rect 716 -649 750 -615
rect 716 -717 750 -683
rect 716 -785 750 -751
rect 804 -105 838 -71
rect 804 -173 838 -139
rect 804 -241 838 -207
rect 804 -309 838 -275
rect 804 -377 838 -343
rect 804 -445 838 -411
rect 804 -513 838 -479
rect 804 -581 838 -547
rect 804 -649 838 -615
rect 804 -717 838 -683
rect 804 -785 838 -751
rect 892 -105 926 -71
rect 892 -173 926 -139
rect 892 -241 926 -207
rect 892 -309 926 -275
rect 892 -377 926 -343
rect 892 -445 926 -411
rect 892 -513 926 -479
rect 892 -581 926 -547
rect 892 -649 926 -615
rect 892 -717 926 -683
rect 892 -785 926 -751
rect 980 -105 1014 -71
rect 980 -173 1014 -139
rect 980 -241 1014 -207
rect 980 -309 1014 -275
rect 980 -377 1014 -343
rect 980 -445 1014 -411
rect 980 -513 1014 -479
rect 980 -581 1014 -547
rect 980 -649 1014 -615
rect 980 -717 1014 -683
rect 980 -785 1014 -751
rect 1068 -105 1102 -71
rect 1068 -173 1102 -139
rect 1068 -241 1102 -207
rect 1068 -309 1102 -275
rect 1068 -377 1102 -343
rect 1068 -445 1102 -411
rect 1068 -513 1102 -479
rect 1068 -581 1102 -547
rect 1068 -649 1102 -615
rect 1068 -717 1102 -683
rect 1068 -785 1102 -751
rect 1156 -105 1190 -71
rect 1156 -173 1190 -139
rect 1156 -241 1190 -207
rect 1156 -309 1190 -275
rect 1156 -377 1190 -343
rect 1156 -445 1190 -411
rect 1156 -513 1190 -479
rect 1156 -581 1190 -547
rect 1156 -649 1190 -615
rect 1156 -717 1190 -683
rect 1156 -785 1190 -751
rect 1244 -105 1278 -71
rect 1244 -173 1278 -139
rect 1244 -241 1278 -207
rect 1244 -309 1278 -275
rect 1244 -377 1278 -343
rect 1244 -445 1278 -411
rect 1244 -513 1278 -479
rect 1244 -581 1278 -547
rect 1244 -649 1278 -615
rect 1244 -717 1278 -683
rect 1244 -785 1278 -751
rect 1332 -105 1366 -71
rect 1332 -173 1366 -139
rect 1332 -241 1366 -207
rect 1332 -309 1366 -275
rect 1332 -377 1366 -343
rect 1332 -445 1366 -411
rect 1332 -513 1366 -479
rect 1332 -581 1366 -547
rect 1332 -649 1366 -615
rect 1332 -717 1366 -683
rect 1332 -785 1366 -751
rect 1420 -105 1454 -71
rect 1420 -173 1454 -139
rect 1420 -241 1454 -207
rect 1420 -309 1454 -275
rect 1420 -377 1454 -343
rect 1420 -445 1454 -411
rect 1420 -513 1454 -479
rect 1420 -581 1454 -547
rect 1420 -649 1454 -615
rect 1420 -717 1454 -683
rect 1420 -785 1454 -751
rect 1508 -105 1542 -71
rect 1508 -173 1542 -139
rect 1508 -241 1542 -207
rect 1508 -309 1542 -275
rect 1508 -377 1542 -343
rect 1508 -445 1542 -411
rect 1508 -513 1542 -479
rect 1508 -581 1542 -547
rect 1508 -649 1542 -615
rect 1508 -717 1542 -683
rect 1508 -785 1542 -751
rect 1596 -105 1630 -71
rect 1596 -173 1630 -139
rect 1596 -241 1630 -207
rect 1596 -309 1630 -275
rect 1596 -377 1630 -343
rect 1596 -445 1630 -411
rect 1596 -513 1630 -479
rect 1596 -581 1630 -547
rect 1596 -649 1630 -615
rect 1596 -717 1630 -683
rect 1596 -785 1630 -751
rect 1684 -105 1718 -71
rect 1684 -173 1718 -139
rect 1684 -241 1718 -207
rect 1684 -309 1718 -275
rect 1684 -377 1718 -343
rect 1684 -445 1718 -411
rect 1684 -513 1718 -479
rect 1684 -581 1718 -547
rect 1684 -649 1718 -615
rect 1684 -717 1718 -683
rect 1684 -785 1718 -751
rect 1772 -105 1806 -71
rect 1772 -173 1806 -139
rect 1772 -241 1806 -207
rect 1772 -309 1806 -275
rect 1772 -377 1806 -343
rect 1772 -445 1806 -411
rect 1772 -513 1806 -479
rect 1772 -581 1806 -547
rect 1772 -649 1806 -615
rect 1772 -717 1806 -683
rect 1772 -785 1806 -751
rect 1860 -105 1894 -71
rect 1860 -173 1894 -139
rect 1860 -241 1894 -207
rect 1860 -309 1894 -275
rect 1860 -377 1894 -343
rect 1860 -445 1894 -411
rect 1860 -513 1894 -479
rect 1860 -581 1894 -547
rect 1860 -649 1894 -615
rect 1860 -717 1894 -683
rect 1860 -785 1894 -751
rect 1948 -105 1982 -71
rect 1948 -173 1982 -139
rect 1948 -241 1982 -207
rect 1948 -309 1982 -275
rect 1948 -377 1982 -343
rect 1948 -445 1982 -411
rect 1948 -513 1982 -479
rect 1948 -581 1982 -547
rect 1948 -649 1982 -615
rect 1948 -717 1982 -683
rect 1948 -785 1982 -751
rect 2036 -105 2070 -71
rect 2036 -173 2070 -139
rect 2036 -241 2070 -207
rect 2036 -309 2070 -275
rect 2036 -377 2070 -343
rect 2036 -445 2070 -411
rect 2036 -513 2070 -479
rect 2036 -581 2070 -547
rect 2036 -649 2070 -615
rect 2036 -717 2070 -683
rect 2036 -785 2070 -751
rect 2124 -105 2158 -71
rect 2124 -173 2158 -139
rect 2124 -241 2158 -207
rect 2124 -309 2158 -275
rect 2124 -377 2158 -343
rect 2124 -445 2158 -411
rect 2124 -513 2158 -479
rect 2124 -581 2158 -547
rect 2124 -649 2158 -615
rect 2124 -717 2158 -683
rect 2124 -785 2158 -751
rect 2212 -105 2246 -71
rect 2212 -173 2246 -139
rect 2212 -241 2246 -207
rect 2212 -309 2246 -275
rect 2212 -377 2246 -343
rect 2212 -445 2246 -411
rect 2212 -513 2246 -479
rect 2212 -581 2246 -547
rect 2212 -649 2246 -615
rect 2212 -717 2246 -683
rect 2212 -785 2246 -751
<< psubdiff >>
rect -229 1100 2520 1116
rect -229 998 78 1100
rect 2356 998 2520 1100
rect -229 982 2520 998
rect -229 881 -115 982
rect -229 -785 -223 881
rect -121 -785 -115 881
rect 2406 857 2520 982
rect -229 -1052 -115 -785
rect 2406 -809 2412 857
rect 2514 -809 2520 857
rect 2406 -1052 2520 -809
rect -229 -1068 2520 -1052
rect -229 -1170 3 -1068
rect 2281 -1170 2520 -1068
rect -229 -1186 2520 -1170
<< psubdiffcont >>
rect 78 998 2356 1100
rect -223 -785 -121 881
rect 2412 -809 2514 857
rect 3 -1170 2281 -1068
<< poly >>
rect 58 914 2200 924
rect 58 880 91 914
rect 125 880 159 914
rect 193 880 227 914
rect 261 880 295 914
rect 329 880 363 914
rect 397 880 431 914
rect 465 880 499 914
rect 533 880 567 914
rect 601 880 635 914
rect 669 880 703 914
rect 737 880 771 914
rect 805 880 839 914
rect 873 880 907 914
rect 941 880 975 914
rect 1009 880 1043 914
rect 1077 880 1111 914
rect 1145 880 1179 914
rect 1213 880 1247 914
rect 1281 880 1315 914
rect 1349 880 1383 914
rect 1417 880 1451 914
rect 1485 880 1519 914
rect 1553 880 1587 914
rect 1621 880 1655 914
rect 1689 880 1723 914
rect 1757 880 1791 914
rect 1825 880 1859 914
rect 1893 880 1927 914
rect 1961 880 1995 914
rect 2029 880 2063 914
rect 2097 880 2131 914
rect 2165 880 2200 914
rect 58 864 2200 880
rect 58 851 88 864
rect 146 826 176 864
rect 234 826 264 864
rect 322 826 352 864
rect 410 826 440 864
rect 498 826 528 864
rect 586 826 616 864
rect 674 826 704 864
rect 762 826 792 864
rect 850 826 880 864
rect 938 826 968 864
rect 1026 826 1056 864
rect 1114 826 1144 864
rect 1202 826 1232 864
rect 1290 826 1320 864
rect 1378 826 1408 864
rect 1466 826 1496 864
rect 1554 826 1584 864
rect 1642 826 1672 864
rect 1730 826 1760 864
rect 1818 826 1848 864
rect 1906 826 1936 864
rect 1994 826 2024 864
rect 2082 826 2112 864
rect 2170 826 2200 864
rect 58 -28 88 11
rect 146 -28 176 26
rect 234 -28 264 26
rect 322 -28 352 26
rect 410 -28 440 26
rect 498 -28 528 26
rect 586 -28 616 26
rect 674 -28 704 26
rect 762 -28 792 26
rect 850 -28 880 26
rect 938 -28 968 26
rect 1026 -28 1056 26
rect 1114 -28 1144 26
rect 1202 -28 1232 26
rect 1290 -28 1320 26
rect 1378 -28 1408 26
rect 1466 -28 1496 26
rect 1554 -28 1584 26
rect 1642 -28 1672 26
rect 1730 -28 1760 26
rect 1818 -28 1848 26
rect 1906 -28 1936 26
rect 1994 -28 2024 26
rect 2082 -28 2112 26
rect 2170 -28 2200 26
rect 58 -866 88 -828
rect 146 -866 176 -828
rect 234 -866 264 -828
rect 322 -866 352 -828
rect 410 -866 440 -828
rect 498 -866 528 -828
rect 586 -866 616 -828
rect 674 -866 704 -828
rect 762 -866 792 -828
rect 850 -866 880 -828
rect 938 -866 968 -828
rect 1026 -866 1056 -828
rect 1114 -866 1144 -828
rect 1202 -866 1232 -828
rect 1290 -866 1320 -828
rect 1378 -866 1408 -828
rect 1466 -866 1496 -828
rect 1554 -866 1584 -828
rect 1642 -866 1672 -828
rect 1730 -866 1760 -828
rect 1818 -866 1848 -828
rect 1906 -866 1936 -828
rect 1994 -866 2024 -828
rect 2082 -866 2112 -828
rect 2170 -866 2200 -828
rect 58 -881 2200 -866
rect 58 -915 91 -881
rect 125 -915 159 -881
rect 193 -915 227 -881
rect 261 -915 295 -881
rect 329 -915 363 -881
rect 397 -915 431 -881
rect 465 -915 499 -881
rect 533 -915 567 -881
rect 601 -915 635 -881
rect 669 -915 703 -881
rect 737 -915 771 -881
rect 805 -915 839 -881
rect 873 -915 907 -881
rect 941 -915 975 -881
rect 1009 -915 1043 -881
rect 1077 -915 1111 -881
rect 1145 -915 1179 -881
rect 1213 -915 1247 -881
rect 1281 -915 1315 -881
rect 1349 -915 1383 -881
rect 1417 -915 1451 -881
rect 1485 -915 1519 -881
rect 1553 -915 1587 -881
rect 1621 -915 1655 -881
rect 1689 -915 1723 -881
rect 1757 -915 1791 -881
rect 1825 -915 1859 -881
rect 1893 -915 1927 -881
rect 1961 -915 1995 -881
rect 2029 -915 2063 -881
rect 2097 -915 2131 -881
rect 2165 -915 2200 -881
rect 58 -926 2200 -915
<< polycont >>
rect 91 880 125 914
rect 159 880 193 914
rect 227 880 261 914
rect 295 880 329 914
rect 363 880 397 914
rect 431 880 465 914
rect 499 880 533 914
rect 567 880 601 914
rect 635 880 669 914
rect 703 880 737 914
rect 771 880 805 914
rect 839 880 873 914
rect 907 880 941 914
rect 975 880 1009 914
rect 1043 880 1077 914
rect 1111 880 1145 914
rect 1179 880 1213 914
rect 1247 880 1281 914
rect 1315 880 1349 914
rect 1383 880 1417 914
rect 1451 880 1485 914
rect 1519 880 1553 914
rect 1587 880 1621 914
rect 1655 880 1689 914
rect 1723 880 1757 914
rect 1791 880 1825 914
rect 1859 880 1893 914
rect 1927 880 1961 914
rect 1995 880 2029 914
rect 2063 880 2097 914
rect 2131 880 2165 914
rect 91 -915 125 -881
rect 159 -915 193 -881
rect 227 -915 261 -881
rect 295 -915 329 -881
rect 363 -915 397 -881
rect 431 -915 465 -881
rect 499 -915 533 -881
rect 567 -915 601 -881
rect 635 -915 669 -881
rect 703 -915 737 -881
rect 771 -915 805 -881
rect 839 -915 873 -881
rect 907 -915 941 -881
rect 975 -915 1009 -881
rect 1043 -915 1077 -881
rect 1111 -915 1145 -881
rect 1179 -915 1213 -881
rect 1247 -915 1281 -881
rect 1315 -915 1349 -881
rect 1383 -915 1417 -881
rect 1451 -915 1485 -881
rect 1519 -915 1553 -881
rect 1587 -915 1621 -881
rect 1655 -915 1689 -881
rect 1723 -915 1757 -881
rect 1791 -915 1825 -881
rect 1859 -915 1893 -881
rect 1927 -915 1961 -881
rect 1995 -915 2029 -881
rect 2063 -915 2097 -881
rect 2131 -915 2165 -881
<< locali >>
rect -229 1100 2520 1116
rect -229 998 78 1100
rect 2356 998 2520 1100
rect -229 982 2520 998
rect -229 881 -115 982
rect -229 -785 -223 881
rect -121 -785 -115 881
rect 58 914 2200 924
rect 58 880 91 914
rect 137 880 159 914
rect 209 880 227 914
rect 281 880 295 914
rect 353 880 363 914
rect 425 880 431 914
rect 497 880 499 914
rect 533 880 535 914
rect 601 880 607 914
rect 669 880 679 914
rect 737 880 751 914
rect 805 880 823 914
rect 873 880 895 914
rect 941 880 967 914
rect 1009 880 1039 914
rect 1077 880 1111 914
rect 1145 880 1179 914
rect 1217 880 1247 914
rect 1289 880 1315 914
rect 1361 880 1383 914
rect 1433 880 1451 914
rect 1505 880 1519 914
rect 1577 880 1587 914
rect 1649 880 1655 914
rect 1721 880 1723 914
rect 1757 880 1759 914
rect 1825 880 1831 914
rect 1893 880 1903 914
rect 1961 880 1975 914
rect 2029 880 2047 914
rect 2097 880 2119 914
rect 2165 880 2200 914
rect 58 864 2200 880
rect 2406 857 2520 982
rect -229 -1052 -115 -785
rect 12 -51 46 26
rect 12 -123 46 -105
rect 12 -195 46 -173
rect 12 -267 46 -241
rect 12 -339 46 -309
rect 12 -411 46 -377
rect 12 -479 46 -445
rect 12 -547 46 -517
rect 12 -615 46 -589
rect 12 -683 46 -661
rect 12 -751 46 -733
rect 12 -832 46 -805
rect 100 -51 134 26
rect 100 -123 134 -105
rect 100 -195 134 -173
rect 100 -267 134 -241
rect 100 -339 134 -309
rect 100 -411 134 -377
rect 100 -479 134 -445
rect 100 -547 134 -517
rect 100 -615 134 -589
rect 100 -683 134 -661
rect 100 -751 134 -733
rect 100 -832 134 -805
rect 188 -51 222 26
rect 188 -123 222 -105
rect 188 -195 222 -173
rect 188 -267 222 -241
rect 188 -339 222 -309
rect 188 -411 222 -377
rect 188 -479 222 -445
rect 188 -547 222 -517
rect 188 -615 222 -589
rect 188 -683 222 -661
rect 188 -751 222 -733
rect 188 -832 222 -805
rect 276 -51 310 26
rect 276 -123 310 -105
rect 276 -195 310 -173
rect 276 -267 310 -241
rect 276 -339 310 -309
rect 276 -411 310 -377
rect 276 -479 310 -445
rect 276 -547 310 -517
rect 276 -615 310 -589
rect 276 -683 310 -661
rect 276 -751 310 -733
rect 276 -832 310 -805
rect 364 -51 398 26
rect 364 -123 398 -105
rect 364 -195 398 -173
rect 364 -267 398 -241
rect 364 -339 398 -309
rect 364 -411 398 -377
rect 364 -479 398 -445
rect 364 -547 398 -517
rect 364 -615 398 -589
rect 364 -683 398 -661
rect 364 -751 398 -733
rect 364 -832 398 -805
rect 452 -51 486 26
rect 452 -123 486 -105
rect 452 -195 486 -173
rect 452 -267 486 -241
rect 452 -339 486 -309
rect 452 -411 486 -377
rect 452 -479 486 -445
rect 452 -547 486 -517
rect 452 -615 486 -589
rect 452 -683 486 -661
rect 452 -751 486 -733
rect 452 -832 486 -805
rect 540 -51 574 26
rect 540 -123 574 -105
rect 540 -195 574 -173
rect 540 -267 574 -241
rect 540 -339 574 -309
rect 540 -411 574 -377
rect 540 -479 574 -445
rect 540 -547 574 -517
rect 540 -615 574 -589
rect 540 -683 574 -661
rect 540 -751 574 -733
rect 540 -832 574 -805
rect 628 -51 662 26
rect 628 -123 662 -105
rect 628 -195 662 -173
rect 628 -267 662 -241
rect 628 -339 662 -309
rect 628 -411 662 -377
rect 628 -479 662 -445
rect 628 -547 662 -517
rect 628 -615 662 -589
rect 628 -683 662 -661
rect 628 -751 662 -733
rect 628 -832 662 -805
rect 716 -51 750 26
rect 716 -123 750 -105
rect 716 -195 750 -173
rect 716 -267 750 -241
rect 716 -339 750 -309
rect 716 -411 750 -377
rect 716 -479 750 -445
rect 716 -547 750 -517
rect 716 -615 750 -589
rect 716 -683 750 -661
rect 716 -751 750 -733
rect 716 -832 750 -805
rect 804 -51 838 26
rect 804 -123 838 -105
rect 804 -195 838 -173
rect 804 -267 838 -241
rect 804 -339 838 -309
rect 804 -411 838 -377
rect 804 -479 838 -445
rect 804 -547 838 -517
rect 804 -615 838 -589
rect 804 -683 838 -661
rect 804 -751 838 -733
rect 804 -832 838 -805
rect 892 -51 926 26
rect 892 -123 926 -105
rect 892 -195 926 -173
rect 892 -267 926 -241
rect 892 -339 926 -309
rect 892 -411 926 -377
rect 892 -479 926 -445
rect 892 -547 926 -517
rect 892 -615 926 -589
rect 892 -683 926 -661
rect 892 -751 926 -733
rect 892 -832 926 -805
rect 980 -51 1014 26
rect 980 -123 1014 -105
rect 980 -195 1014 -173
rect 980 -267 1014 -241
rect 980 -339 1014 -309
rect 980 -411 1014 -377
rect 980 -479 1014 -445
rect 980 -547 1014 -517
rect 980 -615 1014 -589
rect 980 -683 1014 -661
rect 980 -751 1014 -733
rect 980 -832 1014 -805
rect 1068 -51 1102 26
rect 1068 -123 1102 -105
rect 1068 -195 1102 -173
rect 1068 -267 1102 -241
rect 1068 -339 1102 -309
rect 1068 -411 1102 -377
rect 1068 -479 1102 -445
rect 1068 -547 1102 -517
rect 1068 -615 1102 -589
rect 1068 -683 1102 -661
rect 1068 -751 1102 -733
rect 1068 -832 1102 -805
rect 1156 -51 1190 26
rect 1156 -123 1190 -105
rect 1156 -195 1190 -173
rect 1156 -267 1190 -241
rect 1156 -339 1190 -309
rect 1156 -411 1190 -377
rect 1156 -479 1190 -445
rect 1156 -547 1190 -517
rect 1156 -615 1190 -589
rect 1156 -683 1190 -661
rect 1156 -751 1190 -733
rect 1156 -832 1190 -805
rect 1244 -51 1278 26
rect 1244 -123 1278 -105
rect 1244 -195 1278 -173
rect 1244 -267 1278 -241
rect 1244 -339 1278 -309
rect 1244 -411 1278 -377
rect 1244 -479 1278 -445
rect 1244 -547 1278 -517
rect 1244 -615 1278 -589
rect 1244 -683 1278 -661
rect 1244 -751 1278 -733
rect 1244 -832 1278 -805
rect 1332 -51 1366 26
rect 1332 -123 1366 -105
rect 1332 -195 1366 -173
rect 1332 -267 1366 -241
rect 1332 -339 1366 -309
rect 1332 -411 1366 -377
rect 1332 -479 1366 -445
rect 1332 -547 1366 -517
rect 1332 -615 1366 -589
rect 1332 -683 1366 -661
rect 1332 -751 1366 -733
rect 1332 -832 1366 -805
rect 1420 -51 1454 26
rect 1420 -123 1454 -105
rect 1420 -195 1454 -173
rect 1420 -267 1454 -241
rect 1420 -339 1454 -309
rect 1420 -411 1454 -377
rect 1420 -479 1454 -445
rect 1420 -547 1454 -517
rect 1420 -615 1454 -589
rect 1420 -683 1454 -661
rect 1420 -751 1454 -733
rect 1420 -832 1454 -805
rect 1508 -51 1542 26
rect 1508 -123 1542 -105
rect 1508 -195 1542 -173
rect 1508 -267 1542 -241
rect 1508 -339 1542 -309
rect 1508 -411 1542 -377
rect 1508 -479 1542 -445
rect 1508 -547 1542 -517
rect 1508 -615 1542 -589
rect 1508 -683 1542 -661
rect 1508 -751 1542 -733
rect 1508 -832 1542 -805
rect 1596 -51 1630 26
rect 1596 -123 1630 -105
rect 1596 -195 1630 -173
rect 1596 -267 1630 -241
rect 1596 -339 1630 -309
rect 1596 -411 1630 -377
rect 1596 -479 1630 -445
rect 1596 -547 1630 -517
rect 1596 -615 1630 -589
rect 1596 -683 1630 -661
rect 1596 -751 1630 -733
rect 1596 -832 1630 -805
rect 1684 -51 1718 26
rect 1684 -123 1718 -105
rect 1684 -195 1718 -173
rect 1684 -267 1718 -241
rect 1684 -339 1718 -309
rect 1684 -411 1718 -377
rect 1684 -479 1718 -445
rect 1684 -547 1718 -517
rect 1684 -615 1718 -589
rect 1684 -683 1718 -661
rect 1684 -751 1718 -733
rect 1684 -832 1718 -805
rect 1772 -51 1806 26
rect 1772 -123 1806 -105
rect 1772 -195 1806 -173
rect 1772 -267 1806 -241
rect 1772 -339 1806 -309
rect 1772 -411 1806 -377
rect 1772 -479 1806 -445
rect 1772 -547 1806 -517
rect 1772 -615 1806 -589
rect 1772 -683 1806 -661
rect 1772 -751 1806 -733
rect 1772 -832 1806 -805
rect 1860 -51 1894 26
rect 1860 -123 1894 -105
rect 1860 -195 1894 -173
rect 1860 -267 1894 -241
rect 1860 -339 1894 -309
rect 1860 -411 1894 -377
rect 1860 -479 1894 -445
rect 1860 -547 1894 -517
rect 1860 -615 1894 -589
rect 1860 -683 1894 -661
rect 1860 -751 1894 -733
rect 1860 -832 1894 -805
rect 1948 -51 1982 26
rect 1948 -123 1982 -105
rect 1948 -195 1982 -173
rect 1948 -267 1982 -241
rect 1948 -339 1982 -309
rect 1948 -411 1982 -377
rect 1948 -479 1982 -445
rect 1948 -547 1982 -517
rect 1948 -615 1982 -589
rect 1948 -683 1982 -661
rect 1948 -751 1982 -733
rect 1948 -832 1982 -805
rect 2036 -51 2070 26
rect 2036 -123 2070 -105
rect 2036 -195 2070 -173
rect 2036 -267 2070 -241
rect 2036 -339 2070 -309
rect 2036 -411 2070 -377
rect 2036 -479 2070 -445
rect 2036 -547 2070 -517
rect 2036 -615 2070 -589
rect 2036 -683 2070 -661
rect 2036 -751 2070 -733
rect 2036 -832 2070 -805
rect 2124 -51 2158 26
rect 2124 -123 2158 -105
rect 2124 -195 2158 -173
rect 2124 -267 2158 -241
rect 2124 -339 2158 -309
rect 2124 -411 2158 -377
rect 2124 -479 2158 -445
rect 2124 -547 2158 -517
rect 2124 -615 2158 -589
rect 2124 -683 2158 -661
rect 2124 -751 2158 -733
rect 2124 -832 2158 -805
rect 2212 -51 2246 26
rect 2212 -123 2246 -105
rect 2212 -195 2246 -173
rect 2212 -267 2246 -241
rect 2212 -339 2246 -309
rect 2212 -411 2246 -377
rect 2212 -479 2246 -445
rect 2212 -547 2246 -517
rect 2212 -615 2246 -589
rect 2212 -683 2246 -661
rect 2212 -751 2246 -733
rect 2212 -832 2246 -805
rect 2406 -809 2412 857
rect 2514 -809 2520 857
rect 58 -881 2200 -866
rect 58 -915 91 -881
rect 137 -915 159 -881
rect 209 -915 227 -881
rect 281 -915 295 -881
rect 353 -915 363 -881
rect 425 -915 431 -881
rect 497 -915 499 -881
rect 533 -915 535 -881
rect 601 -915 607 -881
rect 669 -915 679 -881
rect 737 -915 751 -881
rect 805 -915 823 -881
rect 873 -915 895 -881
rect 941 -915 967 -881
rect 1009 -915 1039 -881
rect 1077 -915 1111 -881
rect 1145 -915 1179 -881
rect 1217 -915 1247 -881
rect 1289 -915 1315 -881
rect 1361 -915 1383 -881
rect 1433 -915 1451 -881
rect 1505 -915 1519 -881
rect 1577 -915 1587 -881
rect 1649 -915 1655 -881
rect 1721 -915 1723 -881
rect 1757 -915 1759 -881
rect 1825 -915 1831 -881
rect 1893 -915 1903 -881
rect 1961 -915 1975 -881
rect 2029 -915 2047 -881
rect 2097 -915 2119 -881
rect 2165 -915 2200 -881
rect 58 -926 2200 -915
rect 2406 -1052 2520 -809
rect -229 -1068 2520 -1052
rect -229 -1170 3 -1068
rect 2281 -1170 2520 -1068
rect -229 -1186 2520 -1170
<< viali >>
rect 103 880 125 914
rect 125 880 137 914
rect 175 880 193 914
rect 193 880 209 914
rect 247 880 261 914
rect 261 880 281 914
rect 319 880 329 914
rect 329 880 353 914
rect 391 880 397 914
rect 397 880 425 914
rect 463 880 465 914
rect 465 880 497 914
rect 535 880 567 914
rect 567 880 569 914
rect 607 880 635 914
rect 635 880 641 914
rect 679 880 703 914
rect 703 880 713 914
rect 751 880 771 914
rect 771 880 785 914
rect 823 880 839 914
rect 839 880 857 914
rect 895 880 907 914
rect 907 880 929 914
rect 967 880 975 914
rect 975 880 1001 914
rect 1039 880 1043 914
rect 1043 880 1073 914
rect 1111 880 1145 914
rect 1183 880 1213 914
rect 1213 880 1217 914
rect 1255 880 1281 914
rect 1281 880 1289 914
rect 1327 880 1349 914
rect 1349 880 1361 914
rect 1399 880 1417 914
rect 1417 880 1433 914
rect 1471 880 1485 914
rect 1485 880 1505 914
rect 1543 880 1553 914
rect 1553 880 1577 914
rect 1615 880 1621 914
rect 1621 880 1649 914
rect 1687 880 1689 914
rect 1689 880 1721 914
rect 1759 880 1791 914
rect 1791 880 1793 914
rect 1831 880 1859 914
rect 1859 880 1865 914
rect 1903 880 1927 914
rect 1927 880 1937 914
rect 1975 880 1995 914
rect 1995 880 2009 914
rect 2047 880 2063 914
rect 2063 880 2081 914
rect 2119 880 2131 914
rect 2131 880 2153 914
rect 12 -71 46 -51
rect 12 -85 46 -71
rect 12 -139 46 -123
rect 12 -157 46 -139
rect 12 -207 46 -195
rect 12 -229 46 -207
rect 12 -275 46 -267
rect 12 -301 46 -275
rect 12 -343 46 -339
rect 12 -373 46 -343
rect 12 -445 46 -411
rect 12 -513 46 -483
rect 12 -517 46 -513
rect 12 -581 46 -555
rect 12 -589 46 -581
rect 12 -649 46 -627
rect 12 -661 46 -649
rect 12 -717 46 -699
rect 12 -733 46 -717
rect 12 -785 46 -771
rect 12 -805 46 -785
rect 100 -71 134 -51
rect 100 -85 134 -71
rect 100 -139 134 -123
rect 100 -157 134 -139
rect 100 -207 134 -195
rect 100 -229 134 -207
rect 100 -275 134 -267
rect 100 -301 134 -275
rect 100 -343 134 -339
rect 100 -373 134 -343
rect 100 -445 134 -411
rect 100 -513 134 -483
rect 100 -517 134 -513
rect 100 -581 134 -555
rect 100 -589 134 -581
rect 100 -649 134 -627
rect 100 -661 134 -649
rect 100 -717 134 -699
rect 100 -733 134 -717
rect 100 -785 134 -771
rect 100 -805 134 -785
rect 188 -71 222 -51
rect 188 -85 222 -71
rect 188 -139 222 -123
rect 188 -157 222 -139
rect 188 -207 222 -195
rect 188 -229 222 -207
rect 188 -275 222 -267
rect 188 -301 222 -275
rect 188 -343 222 -339
rect 188 -373 222 -343
rect 188 -445 222 -411
rect 188 -513 222 -483
rect 188 -517 222 -513
rect 188 -581 222 -555
rect 188 -589 222 -581
rect 188 -649 222 -627
rect 188 -661 222 -649
rect 188 -717 222 -699
rect 188 -733 222 -717
rect 188 -785 222 -771
rect 188 -805 222 -785
rect 276 -71 310 -51
rect 276 -85 310 -71
rect 276 -139 310 -123
rect 276 -157 310 -139
rect 276 -207 310 -195
rect 276 -229 310 -207
rect 276 -275 310 -267
rect 276 -301 310 -275
rect 276 -343 310 -339
rect 276 -373 310 -343
rect 276 -445 310 -411
rect 276 -513 310 -483
rect 276 -517 310 -513
rect 276 -581 310 -555
rect 276 -589 310 -581
rect 276 -649 310 -627
rect 276 -661 310 -649
rect 276 -717 310 -699
rect 276 -733 310 -717
rect 276 -785 310 -771
rect 276 -805 310 -785
rect 364 -71 398 -51
rect 364 -85 398 -71
rect 364 -139 398 -123
rect 364 -157 398 -139
rect 364 -207 398 -195
rect 364 -229 398 -207
rect 364 -275 398 -267
rect 364 -301 398 -275
rect 364 -343 398 -339
rect 364 -373 398 -343
rect 364 -445 398 -411
rect 364 -513 398 -483
rect 364 -517 398 -513
rect 364 -581 398 -555
rect 364 -589 398 -581
rect 364 -649 398 -627
rect 364 -661 398 -649
rect 364 -717 398 -699
rect 364 -733 398 -717
rect 364 -785 398 -771
rect 364 -805 398 -785
rect 452 -71 486 -51
rect 452 -85 486 -71
rect 452 -139 486 -123
rect 452 -157 486 -139
rect 452 -207 486 -195
rect 452 -229 486 -207
rect 452 -275 486 -267
rect 452 -301 486 -275
rect 452 -343 486 -339
rect 452 -373 486 -343
rect 452 -445 486 -411
rect 452 -513 486 -483
rect 452 -517 486 -513
rect 452 -581 486 -555
rect 452 -589 486 -581
rect 452 -649 486 -627
rect 452 -661 486 -649
rect 452 -717 486 -699
rect 452 -733 486 -717
rect 452 -785 486 -771
rect 452 -805 486 -785
rect 540 -71 574 -51
rect 540 -85 574 -71
rect 540 -139 574 -123
rect 540 -157 574 -139
rect 540 -207 574 -195
rect 540 -229 574 -207
rect 540 -275 574 -267
rect 540 -301 574 -275
rect 540 -343 574 -339
rect 540 -373 574 -343
rect 540 -445 574 -411
rect 540 -513 574 -483
rect 540 -517 574 -513
rect 540 -581 574 -555
rect 540 -589 574 -581
rect 540 -649 574 -627
rect 540 -661 574 -649
rect 540 -717 574 -699
rect 540 -733 574 -717
rect 540 -785 574 -771
rect 540 -805 574 -785
rect 628 -71 662 -51
rect 628 -85 662 -71
rect 628 -139 662 -123
rect 628 -157 662 -139
rect 628 -207 662 -195
rect 628 -229 662 -207
rect 628 -275 662 -267
rect 628 -301 662 -275
rect 628 -343 662 -339
rect 628 -373 662 -343
rect 628 -445 662 -411
rect 628 -513 662 -483
rect 628 -517 662 -513
rect 628 -581 662 -555
rect 628 -589 662 -581
rect 628 -649 662 -627
rect 628 -661 662 -649
rect 628 -717 662 -699
rect 628 -733 662 -717
rect 628 -785 662 -771
rect 628 -805 662 -785
rect 716 -71 750 -51
rect 716 -85 750 -71
rect 716 -139 750 -123
rect 716 -157 750 -139
rect 716 -207 750 -195
rect 716 -229 750 -207
rect 716 -275 750 -267
rect 716 -301 750 -275
rect 716 -343 750 -339
rect 716 -373 750 -343
rect 716 -445 750 -411
rect 716 -513 750 -483
rect 716 -517 750 -513
rect 716 -581 750 -555
rect 716 -589 750 -581
rect 716 -649 750 -627
rect 716 -661 750 -649
rect 716 -717 750 -699
rect 716 -733 750 -717
rect 716 -785 750 -771
rect 716 -805 750 -785
rect 804 -71 838 -51
rect 804 -85 838 -71
rect 804 -139 838 -123
rect 804 -157 838 -139
rect 804 -207 838 -195
rect 804 -229 838 -207
rect 804 -275 838 -267
rect 804 -301 838 -275
rect 804 -343 838 -339
rect 804 -373 838 -343
rect 804 -445 838 -411
rect 804 -513 838 -483
rect 804 -517 838 -513
rect 804 -581 838 -555
rect 804 -589 838 -581
rect 804 -649 838 -627
rect 804 -661 838 -649
rect 804 -717 838 -699
rect 804 -733 838 -717
rect 804 -785 838 -771
rect 804 -805 838 -785
rect 892 -71 926 -51
rect 892 -85 926 -71
rect 892 -139 926 -123
rect 892 -157 926 -139
rect 892 -207 926 -195
rect 892 -229 926 -207
rect 892 -275 926 -267
rect 892 -301 926 -275
rect 892 -343 926 -339
rect 892 -373 926 -343
rect 892 -445 926 -411
rect 892 -513 926 -483
rect 892 -517 926 -513
rect 892 -581 926 -555
rect 892 -589 926 -581
rect 892 -649 926 -627
rect 892 -661 926 -649
rect 892 -717 926 -699
rect 892 -733 926 -717
rect 892 -785 926 -771
rect 892 -805 926 -785
rect 980 -71 1014 -51
rect 980 -85 1014 -71
rect 980 -139 1014 -123
rect 980 -157 1014 -139
rect 980 -207 1014 -195
rect 980 -229 1014 -207
rect 980 -275 1014 -267
rect 980 -301 1014 -275
rect 980 -343 1014 -339
rect 980 -373 1014 -343
rect 980 -445 1014 -411
rect 980 -513 1014 -483
rect 980 -517 1014 -513
rect 980 -581 1014 -555
rect 980 -589 1014 -581
rect 980 -649 1014 -627
rect 980 -661 1014 -649
rect 980 -717 1014 -699
rect 980 -733 1014 -717
rect 980 -785 1014 -771
rect 980 -805 1014 -785
rect 1068 -71 1102 -51
rect 1068 -85 1102 -71
rect 1068 -139 1102 -123
rect 1068 -157 1102 -139
rect 1068 -207 1102 -195
rect 1068 -229 1102 -207
rect 1068 -275 1102 -267
rect 1068 -301 1102 -275
rect 1068 -343 1102 -339
rect 1068 -373 1102 -343
rect 1068 -445 1102 -411
rect 1068 -513 1102 -483
rect 1068 -517 1102 -513
rect 1068 -581 1102 -555
rect 1068 -589 1102 -581
rect 1068 -649 1102 -627
rect 1068 -661 1102 -649
rect 1068 -717 1102 -699
rect 1068 -733 1102 -717
rect 1068 -785 1102 -771
rect 1068 -805 1102 -785
rect 1156 -71 1190 -51
rect 1156 -85 1190 -71
rect 1156 -139 1190 -123
rect 1156 -157 1190 -139
rect 1156 -207 1190 -195
rect 1156 -229 1190 -207
rect 1156 -275 1190 -267
rect 1156 -301 1190 -275
rect 1156 -343 1190 -339
rect 1156 -373 1190 -343
rect 1156 -445 1190 -411
rect 1156 -513 1190 -483
rect 1156 -517 1190 -513
rect 1156 -581 1190 -555
rect 1156 -589 1190 -581
rect 1156 -649 1190 -627
rect 1156 -661 1190 -649
rect 1156 -717 1190 -699
rect 1156 -733 1190 -717
rect 1156 -785 1190 -771
rect 1156 -805 1190 -785
rect 1244 -71 1278 -51
rect 1244 -85 1278 -71
rect 1244 -139 1278 -123
rect 1244 -157 1278 -139
rect 1244 -207 1278 -195
rect 1244 -229 1278 -207
rect 1244 -275 1278 -267
rect 1244 -301 1278 -275
rect 1244 -343 1278 -339
rect 1244 -373 1278 -343
rect 1244 -445 1278 -411
rect 1244 -513 1278 -483
rect 1244 -517 1278 -513
rect 1244 -581 1278 -555
rect 1244 -589 1278 -581
rect 1244 -649 1278 -627
rect 1244 -661 1278 -649
rect 1244 -717 1278 -699
rect 1244 -733 1278 -717
rect 1244 -785 1278 -771
rect 1244 -805 1278 -785
rect 1332 -71 1366 -51
rect 1332 -85 1366 -71
rect 1332 -139 1366 -123
rect 1332 -157 1366 -139
rect 1332 -207 1366 -195
rect 1332 -229 1366 -207
rect 1332 -275 1366 -267
rect 1332 -301 1366 -275
rect 1332 -343 1366 -339
rect 1332 -373 1366 -343
rect 1332 -445 1366 -411
rect 1332 -513 1366 -483
rect 1332 -517 1366 -513
rect 1332 -581 1366 -555
rect 1332 -589 1366 -581
rect 1332 -649 1366 -627
rect 1332 -661 1366 -649
rect 1332 -717 1366 -699
rect 1332 -733 1366 -717
rect 1332 -785 1366 -771
rect 1332 -805 1366 -785
rect 1420 -71 1454 -51
rect 1420 -85 1454 -71
rect 1420 -139 1454 -123
rect 1420 -157 1454 -139
rect 1420 -207 1454 -195
rect 1420 -229 1454 -207
rect 1420 -275 1454 -267
rect 1420 -301 1454 -275
rect 1420 -343 1454 -339
rect 1420 -373 1454 -343
rect 1420 -445 1454 -411
rect 1420 -513 1454 -483
rect 1420 -517 1454 -513
rect 1420 -581 1454 -555
rect 1420 -589 1454 -581
rect 1420 -649 1454 -627
rect 1420 -661 1454 -649
rect 1420 -717 1454 -699
rect 1420 -733 1454 -717
rect 1420 -785 1454 -771
rect 1420 -805 1454 -785
rect 1508 -71 1542 -51
rect 1508 -85 1542 -71
rect 1508 -139 1542 -123
rect 1508 -157 1542 -139
rect 1508 -207 1542 -195
rect 1508 -229 1542 -207
rect 1508 -275 1542 -267
rect 1508 -301 1542 -275
rect 1508 -343 1542 -339
rect 1508 -373 1542 -343
rect 1508 -445 1542 -411
rect 1508 -513 1542 -483
rect 1508 -517 1542 -513
rect 1508 -581 1542 -555
rect 1508 -589 1542 -581
rect 1508 -649 1542 -627
rect 1508 -661 1542 -649
rect 1508 -717 1542 -699
rect 1508 -733 1542 -717
rect 1508 -785 1542 -771
rect 1508 -805 1542 -785
rect 1596 -71 1630 -51
rect 1596 -85 1630 -71
rect 1596 -139 1630 -123
rect 1596 -157 1630 -139
rect 1596 -207 1630 -195
rect 1596 -229 1630 -207
rect 1596 -275 1630 -267
rect 1596 -301 1630 -275
rect 1596 -343 1630 -339
rect 1596 -373 1630 -343
rect 1596 -445 1630 -411
rect 1596 -513 1630 -483
rect 1596 -517 1630 -513
rect 1596 -581 1630 -555
rect 1596 -589 1630 -581
rect 1596 -649 1630 -627
rect 1596 -661 1630 -649
rect 1596 -717 1630 -699
rect 1596 -733 1630 -717
rect 1596 -785 1630 -771
rect 1596 -805 1630 -785
rect 1684 -71 1718 -51
rect 1684 -85 1718 -71
rect 1684 -139 1718 -123
rect 1684 -157 1718 -139
rect 1684 -207 1718 -195
rect 1684 -229 1718 -207
rect 1684 -275 1718 -267
rect 1684 -301 1718 -275
rect 1684 -343 1718 -339
rect 1684 -373 1718 -343
rect 1684 -445 1718 -411
rect 1684 -513 1718 -483
rect 1684 -517 1718 -513
rect 1684 -581 1718 -555
rect 1684 -589 1718 -581
rect 1684 -649 1718 -627
rect 1684 -661 1718 -649
rect 1684 -717 1718 -699
rect 1684 -733 1718 -717
rect 1684 -785 1718 -771
rect 1684 -805 1718 -785
rect 1772 -71 1806 -51
rect 1772 -85 1806 -71
rect 1772 -139 1806 -123
rect 1772 -157 1806 -139
rect 1772 -207 1806 -195
rect 1772 -229 1806 -207
rect 1772 -275 1806 -267
rect 1772 -301 1806 -275
rect 1772 -343 1806 -339
rect 1772 -373 1806 -343
rect 1772 -445 1806 -411
rect 1772 -513 1806 -483
rect 1772 -517 1806 -513
rect 1772 -581 1806 -555
rect 1772 -589 1806 -581
rect 1772 -649 1806 -627
rect 1772 -661 1806 -649
rect 1772 -717 1806 -699
rect 1772 -733 1806 -717
rect 1772 -785 1806 -771
rect 1772 -805 1806 -785
rect 1860 -71 1894 -51
rect 1860 -85 1894 -71
rect 1860 -139 1894 -123
rect 1860 -157 1894 -139
rect 1860 -207 1894 -195
rect 1860 -229 1894 -207
rect 1860 -275 1894 -267
rect 1860 -301 1894 -275
rect 1860 -343 1894 -339
rect 1860 -373 1894 -343
rect 1860 -445 1894 -411
rect 1860 -513 1894 -483
rect 1860 -517 1894 -513
rect 1860 -581 1894 -555
rect 1860 -589 1894 -581
rect 1860 -649 1894 -627
rect 1860 -661 1894 -649
rect 1860 -717 1894 -699
rect 1860 -733 1894 -717
rect 1860 -785 1894 -771
rect 1860 -805 1894 -785
rect 1948 -71 1982 -51
rect 1948 -85 1982 -71
rect 1948 -139 1982 -123
rect 1948 -157 1982 -139
rect 1948 -207 1982 -195
rect 1948 -229 1982 -207
rect 1948 -275 1982 -267
rect 1948 -301 1982 -275
rect 1948 -343 1982 -339
rect 1948 -373 1982 -343
rect 1948 -445 1982 -411
rect 1948 -513 1982 -483
rect 1948 -517 1982 -513
rect 1948 -581 1982 -555
rect 1948 -589 1982 -581
rect 1948 -649 1982 -627
rect 1948 -661 1982 -649
rect 1948 -717 1982 -699
rect 1948 -733 1982 -717
rect 1948 -785 1982 -771
rect 1948 -805 1982 -785
rect 2036 -71 2070 -51
rect 2036 -85 2070 -71
rect 2036 -139 2070 -123
rect 2036 -157 2070 -139
rect 2036 -207 2070 -195
rect 2036 -229 2070 -207
rect 2036 -275 2070 -267
rect 2036 -301 2070 -275
rect 2036 -343 2070 -339
rect 2036 -373 2070 -343
rect 2036 -445 2070 -411
rect 2036 -513 2070 -483
rect 2036 -517 2070 -513
rect 2036 -581 2070 -555
rect 2036 -589 2070 -581
rect 2036 -649 2070 -627
rect 2036 -661 2070 -649
rect 2036 -717 2070 -699
rect 2036 -733 2070 -717
rect 2036 -785 2070 -771
rect 2036 -805 2070 -785
rect 2124 -71 2158 -51
rect 2124 -85 2158 -71
rect 2124 -139 2158 -123
rect 2124 -157 2158 -139
rect 2124 -207 2158 -195
rect 2124 -229 2158 -207
rect 2124 -275 2158 -267
rect 2124 -301 2158 -275
rect 2124 -343 2158 -339
rect 2124 -373 2158 -343
rect 2124 -445 2158 -411
rect 2124 -513 2158 -483
rect 2124 -517 2158 -513
rect 2124 -581 2158 -555
rect 2124 -589 2158 -581
rect 2124 -649 2158 -627
rect 2124 -661 2158 -649
rect 2124 -717 2158 -699
rect 2124 -733 2158 -717
rect 2124 -785 2158 -771
rect 2124 -805 2158 -785
rect 2212 -71 2246 -51
rect 2212 -85 2246 -71
rect 2212 -139 2246 -123
rect 2212 -157 2246 -139
rect 2212 -207 2246 -195
rect 2212 -229 2246 -207
rect 2212 -275 2246 -267
rect 2212 -301 2246 -275
rect 2212 -343 2246 -339
rect 2212 -373 2246 -343
rect 2212 -445 2246 -411
rect 2212 -513 2246 -483
rect 2212 -517 2246 -513
rect 2212 -581 2246 -555
rect 2212 -589 2246 -581
rect 2212 -649 2246 -627
rect 2212 -661 2246 -649
rect 2212 -717 2246 -699
rect 2212 -733 2246 -717
rect 2212 -785 2246 -771
rect 2212 -805 2246 -785
rect 103 -915 125 -881
rect 125 -915 137 -881
rect 175 -915 193 -881
rect 193 -915 209 -881
rect 247 -915 261 -881
rect 261 -915 281 -881
rect 319 -915 329 -881
rect 329 -915 353 -881
rect 391 -915 397 -881
rect 397 -915 425 -881
rect 463 -915 465 -881
rect 465 -915 497 -881
rect 535 -915 567 -881
rect 567 -915 569 -881
rect 607 -915 635 -881
rect 635 -915 641 -881
rect 679 -915 703 -881
rect 703 -915 713 -881
rect 751 -915 771 -881
rect 771 -915 785 -881
rect 823 -915 839 -881
rect 839 -915 857 -881
rect 895 -915 907 -881
rect 907 -915 929 -881
rect 967 -915 975 -881
rect 975 -915 1001 -881
rect 1039 -915 1043 -881
rect 1043 -915 1073 -881
rect 1111 -915 1145 -881
rect 1183 -915 1213 -881
rect 1213 -915 1217 -881
rect 1255 -915 1281 -881
rect 1281 -915 1289 -881
rect 1327 -915 1349 -881
rect 1349 -915 1361 -881
rect 1399 -915 1417 -881
rect 1417 -915 1433 -881
rect 1471 -915 1485 -881
rect 1485 -915 1505 -881
rect 1543 -915 1553 -881
rect 1553 -915 1577 -881
rect 1615 -915 1621 -881
rect 1621 -915 1649 -881
rect 1687 -915 1689 -881
rect 1689 -915 1721 -881
rect 1759 -915 1791 -881
rect 1791 -915 1793 -881
rect 1831 -915 1859 -881
rect 1859 -915 1865 -881
rect 1903 -915 1927 -881
rect 1927 -915 1937 -881
rect 1975 -915 1995 -881
rect 1995 -915 2009 -881
rect 2047 -915 2063 -881
rect 2063 -915 2081 -881
rect 2119 -915 2131 -881
rect 2131 -915 2153 -881
<< metal1 >>
rect 56 1299 2201 1403
rect 56 991 177 1299
rect 2085 991 2201 1299
rect 56 914 2201 991
rect 56 880 103 914
rect 137 880 175 914
rect 209 880 247 914
rect 281 880 319 914
rect 353 880 391 914
rect 425 880 463 914
rect 497 880 535 914
rect 569 880 607 914
rect 641 880 679 914
rect 713 880 751 914
rect 785 880 823 914
rect 857 880 895 914
rect 929 880 967 914
rect 1001 880 1039 914
rect 1073 880 1111 914
rect 1145 880 1183 914
rect 1217 880 1255 914
rect 1289 880 1327 914
rect 1361 880 1399 914
rect 1433 880 1471 914
rect 1505 880 1543 914
rect 1577 880 1615 914
rect 1649 880 1687 914
rect 1721 880 1759 914
rect 1793 880 1831 914
rect 1865 880 1903 914
rect 1937 880 1975 914
rect 2009 880 2047 914
rect 2081 880 2119 914
rect 2153 880 2201 914
rect 56 864 2201 880
rect 0 800 64 816
rect 0 748 6 800
rect 58 748 64 800
rect 0 736 64 748
rect 0 684 6 736
rect 58 684 64 736
rect 0 667 64 684
rect 176 800 240 816
rect 176 748 182 800
rect 234 748 240 800
rect 176 736 240 748
rect 176 684 182 736
rect 234 684 240 736
rect 176 667 240 684
rect 352 800 416 816
rect 352 748 358 800
rect 410 748 416 800
rect 352 736 416 748
rect 352 684 358 736
rect 410 684 416 736
rect 352 667 416 684
rect 528 800 592 816
rect 528 748 534 800
rect 586 748 592 800
rect 528 736 592 748
rect 528 684 534 736
rect 586 684 592 736
rect 528 667 592 684
rect 704 800 768 816
rect 704 748 710 800
rect 762 748 768 800
rect 704 736 768 748
rect 704 684 710 736
rect 762 684 768 736
rect 704 667 768 684
rect 880 800 944 816
rect 880 748 886 800
rect 938 748 944 800
rect 880 736 944 748
rect 880 684 886 736
rect 938 684 944 736
rect 880 667 944 684
rect 1056 800 1120 816
rect 1056 748 1062 800
rect 1114 748 1120 800
rect 1056 736 1120 748
rect 1056 684 1062 736
rect 1114 684 1120 736
rect 1056 667 1120 684
rect 1232 800 1296 816
rect 1232 748 1238 800
rect 1290 748 1296 800
rect 1232 736 1296 748
rect 1232 684 1238 736
rect 1290 684 1296 736
rect 1232 667 1296 684
rect 1408 800 1472 816
rect 1408 748 1414 800
rect 1466 748 1472 800
rect 1408 736 1472 748
rect 1408 684 1414 736
rect 1466 684 1472 736
rect 1408 667 1472 684
rect 1584 800 1648 816
rect 1584 748 1590 800
rect 1642 748 1648 800
rect 1584 736 1648 748
rect 1584 684 1590 736
rect 1642 684 1648 736
rect 1584 667 1648 684
rect 1760 800 1824 816
rect 1760 748 1766 800
rect 1818 748 1824 800
rect 1760 736 1824 748
rect 1760 684 1766 736
rect 1818 684 1824 736
rect 1760 667 1824 684
rect 1936 800 2000 816
rect 1936 748 1942 800
rect 1994 748 2000 800
rect 1936 736 2000 748
rect 1936 684 1942 736
rect 1994 684 2000 736
rect 1936 667 2000 684
rect 2112 800 2176 816
rect 2112 748 2118 800
rect 2170 748 2176 800
rect 2112 736 2176 748
rect 2112 684 2118 736
rect 2170 684 2176 736
rect 2112 667 2176 684
rect 0 547 64 563
rect 0 495 6 547
rect 58 495 64 547
rect 0 483 64 495
rect 0 431 6 483
rect 58 431 64 483
rect 0 415 64 431
rect 176 547 240 563
rect 176 495 182 547
rect 234 495 240 547
rect 176 483 240 495
rect 176 431 182 483
rect 234 431 240 483
rect 176 415 240 431
rect 352 547 416 563
rect 352 495 358 547
rect 410 495 416 547
rect 352 483 416 495
rect 352 431 358 483
rect 410 431 416 483
rect 352 415 416 431
rect 528 547 592 563
rect 528 495 534 547
rect 586 495 592 547
rect 528 483 592 495
rect 528 431 534 483
rect 586 431 592 483
rect 528 415 592 431
rect 704 547 768 563
rect 704 495 710 547
rect 762 495 768 547
rect 704 483 768 495
rect 704 431 710 483
rect 762 431 768 483
rect 704 415 768 431
rect 880 547 944 563
rect 880 495 886 547
rect 938 495 944 547
rect 880 483 944 495
rect 880 431 886 483
rect 938 431 944 483
rect 880 415 944 431
rect 1056 547 1120 563
rect 1056 495 1062 547
rect 1114 495 1120 547
rect 1056 483 1120 495
rect 1056 431 1062 483
rect 1114 431 1120 483
rect 1056 415 1120 431
rect 1232 547 1296 563
rect 1232 495 1238 547
rect 1290 495 1296 547
rect 1232 483 1296 495
rect 1232 431 1238 483
rect 1290 431 1296 483
rect 1232 415 1296 431
rect 1408 547 1472 563
rect 1408 495 1414 547
rect 1466 495 1472 547
rect 1408 483 1472 495
rect 1408 431 1414 483
rect 1466 431 1472 483
rect 1408 415 1472 431
rect 1584 547 1648 563
rect 1584 495 1590 547
rect 1642 495 1648 547
rect 1584 483 1648 495
rect 1584 431 1590 483
rect 1642 431 1648 483
rect 1584 415 1648 431
rect 1760 547 1824 563
rect 1760 495 1766 547
rect 1818 495 1824 547
rect 1760 483 1824 495
rect 1760 431 1766 483
rect 1818 431 1824 483
rect 1760 415 1824 431
rect 1936 547 2000 563
rect 1936 495 1942 547
rect 1994 495 2000 547
rect 1936 483 2000 495
rect 1936 431 1942 483
rect 1994 431 2000 483
rect 1936 415 2000 431
rect 2112 547 2176 563
rect 2112 495 2118 547
rect 2170 495 2176 547
rect 2112 483 2176 495
rect 2112 431 2118 483
rect 2170 431 2176 483
rect 2112 415 2176 431
rect 12 309 64 315
rect 188 309 240 315
rect 364 309 416 315
rect 540 309 592 315
rect 716 309 768 315
rect 892 309 944 315
rect 1068 309 1120 315
rect 1244 309 1296 315
rect 1420 309 1472 315
rect 1596 309 1648 315
rect 1772 309 1824 315
rect 1948 309 2000 315
rect 2124 309 2176 315
rect 6 299 64 309
rect 58 247 64 299
rect 6 235 64 247
rect 58 183 64 235
rect 6 173 64 183
rect 182 299 240 309
rect 234 247 240 299
rect 182 235 240 247
rect 234 183 240 235
rect 182 173 240 183
rect 358 299 416 309
rect 410 247 416 299
rect 358 235 416 247
rect 410 183 416 235
rect 358 173 416 183
rect 534 299 592 309
rect 586 247 592 299
rect 534 235 592 247
rect 586 183 592 235
rect 534 173 592 183
rect 710 299 768 309
rect 762 247 768 299
rect 710 235 768 247
rect 762 183 768 235
rect 710 173 768 183
rect 886 299 944 309
rect 938 247 944 299
rect 886 235 944 247
rect 938 183 944 235
rect 886 173 944 183
rect 1062 299 1120 309
rect 1114 247 1120 299
rect 1062 235 1120 247
rect 1114 183 1120 235
rect 1062 173 1120 183
rect 1238 299 1296 309
rect 1290 247 1296 299
rect 1238 235 1296 247
rect 1290 183 1296 235
rect 1238 173 1296 183
rect 1414 299 1472 309
rect 1466 247 1472 299
rect 1414 235 1472 247
rect 1466 183 1472 235
rect 1414 173 1472 183
rect 1590 299 1648 309
rect 1642 247 1648 299
rect 1590 235 1648 247
rect 1642 183 1648 235
rect 1590 173 1648 183
rect 1766 299 1824 309
rect 1818 247 1824 299
rect 1766 235 1824 247
rect 1818 183 1824 235
rect 1766 173 1824 183
rect 1942 299 2000 309
rect 1994 247 2000 299
rect 1942 235 2000 247
rect 1994 183 2000 235
rect 1942 173 2000 183
rect 2118 299 2176 309
rect 2170 247 2176 299
rect 2118 235 2176 247
rect 2170 183 2176 235
rect 2118 173 2176 183
rect 12 167 64 173
rect 188 167 240 173
rect 364 167 416 173
rect 540 167 592 173
rect 716 167 768 173
rect 892 167 944 173
rect 1068 167 1120 173
rect 1244 167 1296 173
rect 1420 167 1472 173
rect 1596 167 1648 173
rect 1772 167 1824 173
rect 1948 167 2000 173
rect 2124 167 2176 173
rect 12 -28 46 26
rect 100 -28 134 26
rect 188 -28 222 26
rect 276 -28 310 26
rect 364 -28 398 26
rect 452 -28 486 26
rect 540 -28 574 26
rect 628 -28 662 26
rect 716 -28 750 26
rect 804 -28 838 26
rect 892 -28 926 26
rect 980 -28 1014 26
rect 1068 -28 1102 26
rect 1156 -28 1190 26
rect 1244 -28 1278 26
rect 1332 -28 1366 26
rect 1420 -28 1454 26
rect 1508 -28 1542 26
rect 1596 -28 1630 26
rect 1684 -28 1718 26
rect 1772 -28 1806 26
rect 1860 -28 1894 26
rect 1948 -28 1982 26
rect 2036 -28 2070 26
rect 2124 -28 2158 26
rect 2212 -28 2246 26
rect 6 -51 52 -28
rect 94 -39 140 -28
rect 6 -85 12 -51
rect 46 -85 52 -51
rect 6 -123 52 -85
rect 6 -157 12 -123
rect 46 -157 52 -123
rect 6 -195 52 -157
rect 85 -51 149 -39
rect 85 -55 100 -51
rect 134 -55 149 -51
rect 85 -107 91 -55
rect 143 -107 149 -55
rect 85 -119 149 -107
rect 85 -171 91 -119
rect 143 -171 149 -119
rect 85 -187 149 -171
rect 182 -51 228 -28
rect 270 -39 316 -28
rect 182 -85 188 -51
rect 222 -85 228 -51
rect 182 -123 228 -85
rect 182 -157 188 -123
rect 222 -157 228 -123
rect 6 -229 12 -195
rect 46 -229 52 -195
rect 6 -267 52 -229
rect 6 -301 12 -267
rect 46 -301 52 -267
rect 94 -195 140 -187
rect 94 -229 100 -195
rect 134 -229 140 -195
rect 94 -267 140 -229
rect 94 -289 100 -267
rect 6 -339 52 -301
rect 6 -373 12 -339
rect 46 -373 52 -339
rect 6 -411 52 -373
rect 6 -445 12 -411
rect 46 -445 52 -411
rect 85 -301 100 -289
rect 134 -289 140 -267
rect 182 -195 228 -157
rect 261 -51 325 -39
rect 261 -55 276 -51
rect 310 -55 325 -51
rect 261 -107 267 -55
rect 319 -107 325 -55
rect 261 -119 325 -107
rect 261 -171 267 -119
rect 319 -171 325 -119
rect 261 -187 325 -171
rect 358 -51 404 -28
rect 446 -39 492 -28
rect 358 -85 364 -51
rect 398 -85 404 -51
rect 358 -123 404 -85
rect 358 -157 364 -123
rect 398 -157 404 -123
rect 182 -229 188 -195
rect 222 -229 228 -195
rect 182 -267 228 -229
rect 134 -301 149 -289
rect 85 -305 149 -301
rect 85 -357 91 -305
rect 143 -357 149 -305
rect 85 -369 100 -357
rect 134 -369 149 -357
rect 85 -421 91 -369
rect 143 -421 149 -369
rect 85 -437 100 -421
rect 6 -483 52 -445
rect 6 -517 12 -483
rect 46 -517 52 -483
rect 6 -555 52 -517
rect 94 -445 100 -437
rect 134 -437 149 -421
rect 182 -301 188 -267
rect 222 -301 228 -267
rect 270 -195 316 -187
rect 270 -229 276 -195
rect 310 -229 316 -195
rect 270 -267 316 -229
rect 270 -289 276 -267
rect 182 -339 228 -301
rect 182 -373 188 -339
rect 222 -373 228 -339
rect 182 -411 228 -373
rect 134 -445 140 -437
rect 94 -483 140 -445
rect 94 -517 100 -483
rect 134 -517 140 -483
rect 94 -539 140 -517
rect 182 -445 188 -411
rect 222 -445 228 -411
rect 261 -301 276 -289
rect 310 -289 316 -267
rect 358 -195 404 -157
rect 437 -51 501 -39
rect 437 -55 452 -51
rect 486 -55 501 -51
rect 437 -107 443 -55
rect 495 -107 501 -55
rect 437 -119 501 -107
rect 437 -171 443 -119
rect 495 -171 501 -119
rect 437 -187 501 -171
rect 534 -51 580 -28
rect 622 -39 668 -28
rect 534 -85 540 -51
rect 574 -85 580 -51
rect 534 -123 580 -85
rect 534 -157 540 -123
rect 574 -157 580 -123
rect 358 -229 364 -195
rect 398 -229 404 -195
rect 358 -267 404 -229
rect 310 -301 325 -289
rect 261 -305 325 -301
rect 261 -357 267 -305
rect 319 -357 325 -305
rect 261 -369 276 -357
rect 310 -369 325 -357
rect 261 -421 267 -369
rect 319 -421 325 -369
rect 261 -437 276 -421
rect 182 -483 228 -445
rect 182 -517 188 -483
rect 222 -517 228 -483
rect 6 -589 12 -555
rect 46 -589 52 -555
rect 6 -627 52 -589
rect 6 -661 12 -627
rect 46 -661 52 -627
rect 6 -699 52 -661
rect 85 -555 149 -539
rect 85 -607 91 -555
rect 143 -607 149 -555
rect 85 -619 149 -607
rect 85 -671 91 -619
rect 143 -671 149 -619
rect 85 -687 149 -671
rect 182 -555 228 -517
rect 270 -445 276 -437
rect 310 -437 325 -421
rect 358 -301 364 -267
rect 398 -301 404 -267
rect 446 -195 492 -187
rect 446 -229 452 -195
rect 486 -229 492 -195
rect 446 -267 492 -229
rect 446 -289 452 -267
rect 358 -339 404 -301
rect 358 -373 364 -339
rect 398 -373 404 -339
rect 358 -411 404 -373
rect 310 -445 316 -437
rect 270 -483 316 -445
rect 270 -517 276 -483
rect 310 -517 316 -483
rect 270 -539 316 -517
rect 358 -445 364 -411
rect 398 -445 404 -411
rect 437 -301 452 -289
rect 486 -289 492 -267
rect 534 -195 580 -157
rect 613 -51 677 -39
rect 613 -55 628 -51
rect 662 -55 677 -51
rect 613 -107 619 -55
rect 671 -107 677 -55
rect 613 -119 677 -107
rect 613 -171 619 -119
rect 671 -171 677 -119
rect 613 -187 677 -171
rect 710 -51 756 -28
rect 798 -39 844 -28
rect 710 -85 716 -51
rect 750 -85 756 -51
rect 710 -123 756 -85
rect 710 -157 716 -123
rect 750 -157 756 -123
rect 534 -229 540 -195
rect 574 -229 580 -195
rect 534 -267 580 -229
rect 486 -301 501 -289
rect 437 -305 501 -301
rect 437 -357 443 -305
rect 495 -357 501 -305
rect 437 -369 452 -357
rect 486 -369 501 -357
rect 437 -421 443 -369
rect 495 -421 501 -369
rect 437 -437 452 -421
rect 358 -483 404 -445
rect 358 -517 364 -483
rect 398 -517 404 -483
rect 182 -589 188 -555
rect 222 -589 228 -555
rect 182 -627 228 -589
rect 182 -661 188 -627
rect 222 -661 228 -627
rect 6 -733 12 -699
rect 46 -733 52 -699
rect 6 -771 52 -733
rect 6 -805 12 -771
rect 46 -805 52 -771
rect 6 -828 52 -805
rect 94 -699 140 -687
rect 94 -733 100 -699
rect 134 -733 140 -699
rect 94 -771 140 -733
rect 94 -805 100 -771
rect 134 -805 140 -771
rect 94 -828 140 -805
rect 182 -699 228 -661
rect 261 -555 325 -539
rect 261 -607 267 -555
rect 319 -607 325 -555
rect 261 -619 325 -607
rect 261 -671 267 -619
rect 319 -671 325 -619
rect 261 -687 325 -671
rect 358 -555 404 -517
rect 446 -445 452 -437
rect 486 -437 501 -421
rect 534 -301 540 -267
rect 574 -301 580 -267
rect 622 -195 668 -187
rect 622 -229 628 -195
rect 662 -229 668 -195
rect 622 -267 668 -229
rect 622 -289 628 -267
rect 534 -339 580 -301
rect 534 -373 540 -339
rect 574 -373 580 -339
rect 534 -411 580 -373
rect 486 -445 492 -437
rect 446 -483 492 -445
rect 446 -517 452 -483
rect 486 -517 492 -483
rect 446 -539 492 -517
rect 534 -445 540 -411
rect 574 -445 580 -411
rect 613 -301 628 -289
rect 662 -289 668 -267
rect 710 -195 756 -157
rect 789 -51 853 -39
rect 789 -55 804 -51
rect 838 -55 853 -51
rect 789 -107 795 -55
rect 847 -107 853 -55
rect 789 -119 853 -107
rect 789 -171 795 -119
rect 847 -171 853 -119
rect 789 -187 853 -171
rect 886 -51 932 -28
rect 974 -39 1020 -28
rect 886 -85 892 -51
rect 926 -85 932 -51
rect 886 -123 932 -85
rect 886 -157 892 -123
rect 926 -157 932 -123
rect 710 -229 716 -195
rect 750 -229 756 -195
rect 710 -267 756 -229
rect 662 -301 677 -289
rect 613 -305 677 -301
rect 613 -357 619 -305
rect 671 -357 677 -305
rect 613 -369 628 -357
rect 662 -369 677 -357
rect 613 -421 619 -369
rect 671 -421 677 -369
rect 613 -437 628 -421
rect 534 -483 580 -445
rect 534 -517 540 -483
rect 574 -517 580 -483
rect 358 -589 364 -555
rect 398 -589 404 -555
rect 358 -627 404 -589
rect 358 -661 364 -627
rect 398 -661 404 -627
rect 182 -733 188 -699
rect 222 -733 228 -699
rect 182 -771 228 -733
rect 182 -805 188 -771
rect 222 -805 228 -771
rect 182 -828 228 -805
rect 270 -699 316 -687
rect 270 -733 276 -699
rect 310 -733 316 -699
rect 270 -771 316 -733
rect 270 -805 276 -771
rect 310 -805 316 -771
rect 270 -828 316 -805
rect 358 -699 404 -661
rect 437 -555 501 -539
rect 437 -607 443 -555
rect 495 -607 501 -555
rect 437 -619 501 -607
rect 437 -671 443 -619
rect 495 -671 501 -619
rect 437 -687 501 -671
rect 534 -555 580 -517
rect 622 -445 628 -437
rect 662 -437 677 -421
rect 710 -301 716 -267
rect 750 -301 756 -267
rect 798 -195 844 -187
rect 798 -229 804 -195
rect 838 -229 844 -195
rect 798 -267 844 -229
rect 798 -289 804 -267
rect 710 -339 756 -301
rect 710 -373 716 -339
rect 750 -373 756 -339
rect 710 -411 756 -373
rect 662 -445 668 -437
rect 622 -483 668 -445
rect 622 -517 628 -483
rect 662 -517 668 -483
rect 622 -539 668 -517
rect 710 -445 716 -411
rect 750 -445 756 -411
rect 789 -301 804 -289
rect 838 -289 844 -267
rect 886 -195 932 -157
rect 965 -51 1029 -39
rect 965 -55 980 -51
rect 1014 -55 1029 -51
rect 965 -107 971 -55
rect 1023 -107 1029 -55
rect 965 -119 1029 -107
rect 965 -171 971 -119
rect 1023 -171 1029 -119
rect 965 -187 1029 -171
rect 1062 -51 1108 -28
rect 1150 -39 1196 -28
rect 1062 -85 1068 -51
rect 1102 -85 1108 -51
rect 1062 -123 1108 -85
rect 1062 -157 1068 -123
rect 1102 -157 1108 -123
rect 886 -229 892 -195
rect 926 -229 932 -195
rect 886 -267 932 -229
rect 838 -301 853 -289
rect 789 -305 853 -301
rect 789 -357 795 -305
rect 847 -357 853 -305
rect 789 -369 804 -357
rect 838 -369 853 -357
rect 789 -421 795 -369
rect 847 -421 853 -369
rect 789 -437 804 -421
rect 710 -483 756 -445
rect 710 -517 716 -483
rect 750 -517 756 -483
rect 534 -589 540 -555
rect 574 -589 580 -555
rect 534 -627 580 -589
rect 534 -661 540 -627
rect 574 -661 580 -627
rect 358 -733 364 -699
rect 398 -733 404 -699
rect 358 -771 404 -733
rect 358 -805 364 -771
rect 398 -805 404 -771
rect 358 -828 404 -805
rect 446 -699 492 -687
rect 446 -733 452 -699
rect 486 -733 492 -699
rect 446 -771 492 -733
rect 446 -805 452 -771
rect 486 -805 492 -771
rect 446 -828 492 -805
rect 534 -699 580 -661
rect 613 -555 677 -539
rect 613 -607 619 -555
rect 671 -607 677 -555
rect 613 -619 677 -607
rect 613 -671 619 -619
rect 671 -671 677 -619
rect 613 -687 677 -671
rect 710 -555 756 -517
rect 798 -445 804 -437
rect 838 -437 853 -421
rect 886 -301 892 -267
rect 926 -301 932 -267
rect 974 -195 1020 -187
rect 974 -229 980 -195
rect 1014 -229 1020 -195
rect 974 -267 1020 -229
rect 974 -289 980 -267
rect 886 -339 932 -301
rect 886 -373 892 -339
rect 926 -373 932 -339
rect 886 -411 932 -373
rect 838 -445 844 -437
rect 798 -483 844 -445
rect 798 -517 804 -483
rect 838 -517 844 -483
rect 798 -539 844 -517
rect 886 -445 892 -411
rect 926 -445 932 -411
rect 965 -301 980 -289
rect 1014 -289 1020 -267
rect 1062 -195 1108 -157
rect 1141 -51 1205 -39
rect 1141 -55 1156 -51
rect 1190 -55 1205 -51
rect 1141 -107 1147 -55
rect 1199 -107 1205 -55
rect 1141 -119 1205 -107
rect 1141 -171 1147 -119
rect 1199 -171 1205 -119
rect 1141 -187 1205 -171
rect 1238 -51 1284 -28
rect 1326 -39 1372 -28
rect 1238 -85 1244 -51
rect 1278 -85 1284 -51
rect 1238 -123 1284 -85
rect 1238 -157 1244 -123
rect 1278 -157 1284 -123
rect 1062 -229 1068 -195
rect 1102 -229 1108 -195
rect 1062 -267 1108 -229
rect 1014 -301 1029 -289
rect 965 -305 1029 -301
rect 965 -357 971 -305
rect 1023 -357 1029 -305
rect 965 -369 980 -357
rect 1014 -369 1029 -357
rect 965 -421 971 -369
rect 1023 -421 1029 -369
rect 965 -437 980 -421
rect 886 -483 932 -445
rect 886 -517 892 -483
rect 926 -517 932 -483
rect 710 -589 716 -555
rect 750 -589 756 -555
rect 710 -627 756 -589
rect 710 -661 716 -627
rect 750 -661 756 -627
rect 534 -733 540 -699
rect 574 -733 580 -699
rect 534 -771 580 -733
rect 534 -805 540 -771
rect 574 -805 580 -771
rect 534 -828 580 -805
rect 622 -699 668 -687
rect 622 -733 628 -699
rect 662 -733 668 -699
rect 622 -771 668 -733
rect 622 -805 628 -771
rect 662 -805 668 -771
rect 622 -828 668 -805
rect 710 -699 756 -661
rect 789 -555 853 -539
rect 789 -607 795 -555
rect 847 -607 853 -555
rect 789 -619 853 -607
rect 789 -671 795 -619
rect 847 -671 853 -619
rect 789 -687 853 -671
rect 886 -555 932 -517
rect 974 -445 980 -437
rect 1014 -437 1029 -421
rect 1062 -301 1068 -267
rect 1102 -301 1108 -267
rect 1150 -195 1196 -187
rect 1150 -229 1156 -195
rect 1190 -229 1196 -195
rect 1150 -267 1196 -229
rect 1150 -289 1156 -267
rect 1062 -339 1108 -301
rect 1062 -373 1068 -339
rect 1102 -373 1108 -339
rect 1062 -411 1108 -373
rect 1014 -445 1020 -437
rect 974 -483 1020 -445
rect 974 -517 980 -483
rect 1014 -517 1020 -483
rect 974 -539 1020 -517
rect 1062 -445 1068 -411
rect 1102 -445 1108 -411
rect 1141 -301 1156 -289
rect 1190 -289 1196 -267
rect 1238 -195 1284 -157
rect 1317 -51 1381 -39
rect 1317 -55 1332 -51
rect 1366 -55 1381 -51
rect 1317 -107 1323 -55
rect 1375 -107 1381 -55
rect 1317 -119 1381 -107
rect 1317 -171 1323 -119
rect 1375 -171 1381 -119
rect 1317 -187 1381 -171
rect 1414 -51 1460 -28
rect 1502 -39 1548 -28
rect 1414 -85 1420 -51
rect 1454 -85 1460 -51
rect 1414 -123 1460 -85
rect 1414 -157 1420 -123
rect 1454 -157 1460 -123
rect 1238 -229 1244 -195
rect 1278 -229 1284 -195
rect 1238 -267 1284 -229
rect 1190 -301 1205 -289
rect 1141 -305 1205 -301
rect 1141 -357 1147 -305
rect 1199 -357 1205 -305
rect 1141 -369 1156 -357
rect 1190 -369 1205 -357
rect 1141 -421 1147 -369
rect 1199 -421 1205 -369
rect 1141 -437 1156 -421
rect 1062 -483 1108 -445
rect 1062 -517 1068 -483
rect 1102 -517 1108 -483
rect 886 -589 892 -555
rect 926 -589 932 -555
rect 886 -627 932 -589
rect 886 -661 892 -627
rect 926 -661 932 -627
rect 710 -733 716 -699
rect 750 -733 756 -699
rect 710 -771 756 -733
rect 710 -805 716 -771
rect 750 -805 756 -771
rect 710 -828 756 -805
rect 798 -699 844 -687
rect 798 -733 804 -699
rect 838 -733 844 -699
rect 798 -771 844 -733
rect 798 -805 804 -771
rect 838 -805 844 -771
rect 798 -828 844 -805
rect 886 -699 932 -661
rect 965 -555 1029 -539
rect 965 -607 971 -555
rect 1023 -607 1029 -555
rect 965 -619 1029 -607
rect 965 -671 971 -619
rect 1023 -671 1029 -619
rect 965 -687 1029 -671
rect 1062 -555 1108 -517
rect 1150 -445 1156 -437
rect 1190 -437 1205 -421
rect 1238 -301 1244 -267
rect 1278 -301 1284 -267
rect 1326 -195 1372 -187
rect 1326 -229 1332 -195
rect 1366 -229 1372 -195
rect 1326 -267 1372 -229
rect 1326 -289 1332 -267
rect 1238 -339 1284 -301
rect 1238 -373 1244 -339
rect 1278 -373 1284 -339
rect 1238 -411 1284 -373
rect 1190 -445 1196 -437
rect 1150 -483 1196 -445
rect 1150 -517 1156 -483
rect 1190 -517 1196 -483
rect 1150 -539 1196 -517
rect 1238 -445 1244 -411
rect 1278 -445 1284 -411
rect 1317 -301 1332 -289
rect 1366 -289 1372 -267
rect 1414 -195 1460 -157
rect 1493 -51 1557 -39
rect 1493 -55 1508 -51
rect 1542 -55 1557 -51
rect 1493 -107 1499 -55
rect 1551 -107 1557 -55
rect 1493 -119 1557 -107
rect 1493 -171 1499 -119
rect 1551 -171 1557 -119
rect 1493 -187 1557 -171
rect 1590 -51 1636 -28
rect 1678 -39 1724 -28
rect 1590 -85 1596 -51
rect 1630 -85 1636 -51
rect 1590 -123 1636 -85
rect 1590 -157 1596 -123
rect 1630 -157 1636 -123
rect 1414 -229 1420 -195
rect 1454 -229 1460 -195
rect 1414 -267 1460 -229
rect 1366 -301 1381 -289
rect 1317 -305 1381 -301
rect 1317 -357 1323 -305
rect 1375 -357 1381 -305
rect 1317 -369 1332 -357
rect 1366 -369 1381 -357
rect 1317 -421 1323 -369
rect 1375 -421 1381 -369
rect 1317 -437 1332 -421
rect 1238 -483 1284 -445
rect 1238 -517 1244 -483
rect 1278 -517 1284 -483
rect 1062 -589 1068 -555
rect 1102 -589 1108 -555
rect 1062 -627 1108 -589
rect 1062 -661 1068 -627
rect 1102 -661 1108 -627
rect 886 -733 892 -699
rect 926 -733 932 -699
rect 886 -771 932 -733
rect 886 -805 892 -771
rect 926 -805 932 -771
rect 886 -828 932 -805
rect 974 -699 1020 -687
rect 974 -733 980 -699
rect 1014 -733 1020 -699
rect 974 -771 1020 -733
rect 974 -805 980 -771
rect 1014 -805 1020 -771
rect 974 -828 1020 -805
rect 1062 -699 1108 -661
rect 1141 -555 1205 -539
rect 1141 -607 1147 -555
rect 1199 -607 1205 -555
rect 1141 -619 1205 -607
rect 1141 -671 1147 -619
rect 1199 -671 1205 -619
rect 1141 -687 1205 -671
rect 1238 -555 1284 -517
rect 1326 -445 1332 -437
rect 1366 -437 1381 -421
rect 1414 -301 1420 -267
rect 1454 -301 1460 -267
rect 1502 -195 1548 -187
rect 1502 -229 1508 -195
rect 1542 -229 1548 -195
rect 1502 -267 1548 -229
rect 1502 -289 1508 -267
rect 1414 -339 1460 -301
rect 1414 -373 1420 -339
rect 1454 -373 1460 -339
rect 1414 -411 1460 -373
rect 1366 -445 1372 -437
rect 1326 -483 1372 -445
rect 1326 -517 1332 -483
rect 1366 -517 1372 -483
rect 1326 -539 1372 -517
rect 1414 -445 1420 -411
rect 1454 -445 1460 -411
rect 1493 -301 1508 -289
rect 1542 -289 1548 -267
rect 1590 -195 1636 -157
rect 1669 -51 1733 -39
rect 1669 -55 1684 -51
rect 1718 -55 1733 -51
rect 1669 -107 1675 -55
rect 1727 -107 1733 -55
rect 1669 -119 1733 -107
rect 1669 -171 1675 -119
rect 1727 -171 1733 -119
rect 1669 -187 1733 -171
rect 1766 -51 1812 -28
rect 1854 -39 1900 -28
rect 1766 -85 1772 -51
rect 1806 -85 1812 -51
rect 1766 -123 1812 -85
rect 1766 -157 1772 -123
rect 1806 -157 1812 -123
rect 1590 -229 1596 -195
rect 1630 -229 1636 -195
rect 1590 -267 1636 -229
rect 1542 -301 1557 -289
rect 1493 -305 1557 -301
rect 1493 -357 1499 -305
rect 1551 -357 1557 -305
rect 1493 -369 1508 -357
rect 1542 -369 1557 -357
rect 1493 -421 1499 -369
rect 1551 -421 1557 -369
rect 1493 -437 1508 -421
rect 1414 -483 1460 -445
rect 1414 -517 1420 -483
rect 1454 -517 1460 -483
rect 1238 -589 1244 -555
rect 1278 -589 1284 -555
rect 1238 -627 1284 -589
rect 1238 -661 1244 -627
rect 1278 -661 1284 -627
rect 1062 -733 1068 -699
rect 1102 -733 1108 -699
rect 1062 -771 1108 -733
rect 1062 -805 1068 -771
rect 1102 -805 1108 -771
rect 1062 -828 1108 -805
rect 1150 -699 1196 -687
rect 1150 -733 1156 -699
rect 1190 -733 1196 -699
rect 1150 -771 1196 -733
rect 1150 -805 1156 -771
rect 1190 -805 1196 -771
rect 1150 -828 1196 -805
rect 1238 -699 1284 -661
rect 1317 -555 1381 -539
rect 1317 -607 1323 -555
rect 1375 -607 1381 -555
rect 1317 -619 1381 -607
rect 1317 -671 1323 -619
rect 1375 -671 1381 -619
rect 1317 -687 1381 -671
rect 1414 -555 1460 -517
rect 1502 -445 1508 -437
rect 1542 -437 1557 -421
rect 1590 -301 1596 -267
rect 1630 -301 1636 -267
rect 1678 -195 1724 -187
rect 1678 -229 1684 -195
rect 1718 -229 1724 -195
rect 1678 -267 1724 -229
rect 1678 -289 1684 -267
rect 1590 -339 1636 -301
rect 1590 -373 1596 -339
rect 1630 -373 1636 -339
rect 1590 -411 1636 -373
rect 1542 -445 1548 -437
rect 1502 -483 1548 -445
rect 1502 -517 1508 -483
rect 1542 -517 1548 -483
rect 1502 -539 1548 -517
rect 1590 -445 1596 -411
rect 1630 -445 1636 -411
rect 1669 -301 1684 -289
rect 1718 -289 1724 -267
rect 1766 -195 1812 -157
rect 1845 -51 1909 -39
rect 1845 -55 1860 -51
rect 1894 -55 1909 -51
rect 1845 -107 1851 -55
rect 1903 -107 1909 -55
rect 1845 -119 1909 -107
rect 1845 -171 1851 -119
rect 1903 -171 1909 -119
rect 1845 -187 1909 -171
rect 1942 -51 1988 -28
rect 2030 -39 2076 -28
rect 1942 -85 1948 -51
rect 1982 -85 1988 -51
rect 1942 -123 1988 -85
rect 1942 -157 1948 -123
rect 1982 -157 1988 -123
rect 1766 -229 1772 -195
rect 1806 -229 1812 -195
rect 1766 -267 1812 -229
rect 1718 -301 1733 -289
rect 1669 -305 1733 -301
rect 1669 -357 1675 -305
rect 1727 -357 1733 -305
rect 1669 -369 1684 -357
rect 1718 -369 1733 -357
rect 1669 -421 1675 -369
rect 1727 -421 1733 -369
rect 1669 -437 1684 -421
rect 1590 -483 1636 -445
rect 1590 -517 1596 -483
rect 1630 -517 1636 -483
rect 1414 -589 1420 -555
rect 1454 -589 1460 -555
rect 1414 -627 1460 -589
rect 1414 -661 1420 -627
rect 1454 -661 1460 -627
rect 1238 -733 1244 -699
rect 1278 -733 1284 -699
rect 1238 -771 1284 -733
rect 1238 -805 1244 -771
rect 1278 -805 1284 -771
rect 1238 -828 1284 -805
rect 1326 -699 1372 -687
rect 1326 -733 1332 -699
rect 1366 -733 1372 -699
rect 1326 -771 1372 -733
rect 1326 -805 1332 -771
rect 1366 -805 1372 -771
rect 1326 -828 1372 -805
rect 1414 -699 1460 -661
rect 1493 -555 1557 -539
rect 1493 -607 1499 -555
rect 1551 -607 1557 -555
rect 1493 -619 1557 -607
rect 1493 -671 1499 -619
rect 1551 -671 1557 -619
rect 1493 -687 1557 -671
rect 1590 -555 1636 -517
rect 1678 -445 1684 -437
rect 1718 -437 1733 -421
rect 1766 -301 1772 -267
rect 1806 -301 1812 -267
rect 1854 -195 1900 -187
rect 1854 -229 1860 -195
rect 1894 -229 1900 -195
rect 1854 -267 1900 -229
rect 1854 -289 1860 -267
rect 1766 -339 1812 -301
rect 1766 -373 1772 -339
rect 1806 -373 1812 -339
rect 1766 -411 1812 -373
rect 1718 -445 1724 -437
rect 1678 -483 1724 -445
rect 1678 -517 1684 -483
rect 1718 -517 1724 -483
rect 1678 -539 1724 -517
rect 1766 -445 1772 -411
rect 1806 -445 1812 -411
rect 1845 -301 1860 -289
rect 1894 -289 1900 -267
rect 1942 -195 1988 -157
rect 2021 -51 2085 -39
rect 2021 -55 2036 -51
rect 2070 -55 2085 -51
rect 2021 -107 2027 -55
rect 2079 -107 2085 -55
rect 2021 -119 2085 -107
rect 2021 -171 2027 -119
rect 2079 -171 2085 -119
rect 2021 -187 2085 -171
rect 2118 -51 2164 -28
rect 2206 -39 2252 -28
rect 2118 -85 2124 -51
rect 2158 -85 2164 -51
rect 2118 -123 2164 -85
rect 2118 -157 2124 -123
rect 2158 -157 2164 -123
rect 1942 -229 1948 -195
rect 1982 -229 1988 -195
rect 1942 -267 1988 -229
rect 1894 -301 1909 -289
rect 1845 -305 1909 -301
rect 1845 -357 1851 -305
rect 1903 -357 1909 -305
rect 1845 -369 1860 -357
rect 1894 -369 1909 -357
rect 1845 -421 1851 -369
rect 1903 -421 1909 -369
rect 1845 -437 1860 -421
rect 1766 -483 1812 -445
rect 1766 -517 1772 -483
rect 1806 -517 1812 -483
rect 1590 -589 1596 -555
rect 1630 -589 1636 -555
rect 1590 -627 1636 -589
rect 1590 -661 1596 -627
rect 1630 -661 1636 -627
rect 1414 -733 1420 -699
rect 1454 -733 1460 -699
rect 1414 -771 1460 -733
rect 1414 -805 1420 -771
rect 1454 -805 1460 -771
rect 1414 -828 1460 -805
rect 1502 -699 1548 -687
rect 1502 -733 1508 -699
rect 1542 -733 1548 -699
rect 1502 -771 1548 -733
rect 1502 -805 1508 -771
rect 1542 -805 1548 -771
rect 1502 -828 1548 -805
rect 1590 -699 1636 -661
rect 1669 -555 1733 -539
rect 1669 -607 1675 -555
rect 1727 -607 1733 -555
rect 1669 -619 1733 -607
rect 1669 -671 1675 -619
rect 1727 -671 1733 -619
rect 1669 -687 1733 -671
rect 1766 -555 1812 -517
rect 1854 -445 1860 -437
rect 1894 -437 1909 -421
rect 1942 -301 1948 -267
rect 1982 -301 1988 -267
rect 2030 -195 2076 -187
rect 2030 -229 2036 -195
rect 2070 -229 2076 -195
rect 2030 -267 2076 -229
rect 2030 -289 2036 -267
rect 1942 -339 1988 -301
rect 1942 -373 1948 -339
rect 1982 -373 1988 -339
rect 1942 -411 1988 -373
rect 1894 -445 1900 -437
rect 1854 -483 1900 -445
rect 1854 -517 1860 -483
rect 1894 -517 1900 -483
rect 1854 -539 1900 -517
rect 1942 -445 1948 -411
rect 1982 -445 1988 -411
rect 2021 -301 2036 -289
rect 2070 -289 2076 -267
rect 2118 -195 2164 -157
rect 2197 -51 2261 -39
rect 2197 -55 2212 -51
rect 2246 -55 2261 -51
rect 2197 -107 2203 -55
rect 2255 -107 2261 -55
rect 2197 -119 2261 -107
rect 2197 -171 2203 -119
rect 2255 -171 2261 -119
rect 2197 -187 2261 -171
rect 2118 -229 2124 -195
rect 2158 -229 2164 -195
rect 2118 -267 2164 -229
rect 2070 -301 2085 -289
rect 2021 -305 2085 -301
rect 2021 -357 2027 -305
rect 2079 -357 2085 -305
rect 2021 -369 2036 -357
rect 2070 -369 2085 -357
rect 2021 -421 2027 -369
rect 2079 -421 2085 -369
rect 2021 -437 2036 -421
rect 1942 -483 1988 -445
rect 1942 -517 1948 -483
rect 1982 -517 1988 -483
rect 1766 -589 1772 -555
rect 1806 -589 1812 -555
rect 1766 -627 1812 -589
rect 1766 -661 1772 -627
rect 1806 -661 1812 -627
rect 1590 -733 1596 -699
rect 1630 -733 1636 -699
rect 1590 -771 1636 -733
rect 1590 -805 1596 -771
rect 1630 -805 1636 -771
rect 1590 -828 1636 -805
rect 1678 -699 1724 -687
rect 1678 -733 1684 -699
rect 1718 -733 1724 -699
rect 1678 -771 1724 -733
rect 1678 -805 1684 -771
rect 1718 -805 1724 -771
rect 1678 -828 1724 -805
rect 1766 -699 1812 -661
rect 1845 -555 1909 -539
rect 1845 -607 1851 -555
rect 1903 -607 1909 -555
rect 1845 -619 1909 -607
rect 1845 -671 1851 -619
rect 1903 -671 1909 -619
rect 1845 -687 1909 -671
rect 1942 -555 1988 -517
rect 2030 -445 2036 -437
rect 2070 -437 2085 -421
rect 2118 -301 2124 -267
rect 2158 -301 2164 -267
rect 2206 -195 2252 -187
rect 2206 -229 2212 -195
rect 2246 -229 2252 -195
rect 2206 -267 2252 -229
rect 2206 -289 2212 -267
rect 2118 -339 2164 -301
rect 2118 -373 2124 -339
rect 2158 -373 2164 -339
rect 2118 -411 2164 -373
rect 2070 -445 2076 -437
rect 2030 -483 2076 -445
rect 2030 -517 2036 -483
rect 2070 -517 2076 -483
rect 2030 -539 2076 -517
rect 2118 -445 2124 -411
rect 2158 -445 2164 -411
rect 2197 -301 2212 -289
rect 2246 -289 2252 -267
rect 2246 -301 2261 -289
rect 2197 -305 2261 -301
rect 2197 -357 2203 -305
rect 2255 -357 2261 -305
rect 2197 -369 2212 -357
rect 2246 -369 2261 -357
rect 2197 -421 2203 -369
rect 2255 -421 2261 -369
rect 2197 -437 2212 -421
rect 2118 -483 2164 -445
rect 2118 -517 2124 -483
rect 2158 -517 2164 -483
rect 1942 -589 1948 -555
rect 1982 -589 1988 -555
rect 1942 -627 1988 -589
rect 1942 -661 1948 -627
rect 1982 -661 1988 -627
rect 1766 -733 1772 -699
rect 1806 -733 1812 -699
rect 1766 -771 1812 -733
rect 1766 -805 1772 -771
rect 1806 -805 1812 -771
rect 1766 -828 1812 -805
rect 1854 -699 1900 -687
rect 1854 -733 1860 -699
rect 1894 -733 1900 -699
rect 1854 -771 1900 -733
rect 1854 -805 1860 -771
rect 1894 -805 1900 -771
rect 1854 -828 1900 -805
rect 1942 -699 1988 -661
rect 2021 -555 2085 -539
rect 2021 -607 2027 -555
rect 2079 -607 2085 -555
rect 2021 -619 2085 -607
rect 2021 -671 2027 -619
rect 2079 -671 2085 -619
rect 2021 -687 2085 -671
rect 2118 -555 2164 -517
rect 2206 -445 2212 -437
rect 2246 -437 2261 -421
rect 2246 -445 2252 -437
rect 2206 -483 2252 -445
rect 2206 -517 2212 -483
rect 2246 -517 2252 -483
rect 2206 -539 2252 -517
rect 2118 -589 2124 -555
rect 2158 -589 2164 -555
rect 2118 -627 2164 -589
rect 2118 -661 2124 -627
rect 2158 -661 2164 -627
rect 1942 -733 1948 -699
rect 1982 -733 1988 -699
rect 1942 -771 1988 -733
rect 1942 -805 1948 -771
rect 1982 -805 1988 -771
rect 1942 -828 1988 -805
rect 2030 -699 2076 -687
rect 2030 -733 2036 -699
rect 2070 -733 2076 -699
rect 2030 -771 2076 -733
rect 2030 -805 2036 -771
rect 2070 -805 2076 -771
rect 2030 -828 2076 -805
rect 2118 -699 2164 -661
rect 2197 -555 2261 -539
rect 2197 -607 2203 -555
rect 2255 -607 2261 -555
rect 2197 -619 2261 -607
rect 2197 -671 2203 -619
rect 2255 -671 2261 -619
rect 2197 -687 2261 -671
rect 2118 -733 2124 -699
rect 2158 -733 2164 -699
rect 2118 -771 2164 -733
rect 2118 -805 2124 -771
rect 2158 -805 2164 -771
rect 2118 -828 2164 -805
rect 2206 -699 2252 -687
rect 2206 -733 2212 -699
rect 2246 -733 2252 -699
rect 2206 -771 2252 -733
rect 2206 -805 2212 -771
rect 2246 -805 2252 -771
rect 2206 -828 2252 -805
rect 57 -881 3371 -865
rect 57 -915 103 -881
rect 137 -915 175 -881
rect 209 -915 247 -881
rect 281 -915 319 -881
rect 353 -915 391 -881
rect 425 -915 463 -881
rect 497 -915 535 -881
rect 569 -915 607 -881
rect 641 -915 679 -881
rect 713 -915 751 -881
rect 785 -915 823 -881
rect 857 -915 895 -881
rect 929 -915 967 -881
rect 1001 -915 1039 -881
rect 1073 -915 1111 -881
rect 1145 -915 1183 -881
rect 1217 -915 1255 -881
rect 1289 -915 1327 -881
rect 1361 -915 1399 -881
rect 1433 -915 1471 -881
rect 1505 -915 1543 -881
rect 1577 -915 1615 -881
rect 1649 -915 1687 -881
rect 1721 -915 1759 -881
rect 1793 -915 1831 -881
rect 1865 -915 1903 -881
rect 1937 -915 1975 -881
rect 2009 -915 2047 -881
rect 2081 -915 2119 -881
rect 2153 -915 3371 -881
rect 57 -1025 3371 -915
<< via1 >>
rect 177 991 2085 1299
rect 6 748 58 800
rect 6 684 58 736
rect 182 748 234 800
rect 182 684 234 736
rect 358 748 410 800
rect 358 684 410 736
rect 534 748 586 800
rect 534 684 586 736
rect 710 748 762 800
rect 710 684 762 736
rect 886 748 938 800
rect 886 684 938 736
rect 1062 748 1114 800
rect 1062 684 1114 736
rect 1238 748 1290 800
rect 1238 684 1290 736
rect 1414 748 1466 800
rect 1414 684 1466 736
rect 1590 748 1642 800
rect 1590 684 1642 736
rect 1766 748 1818 800
rect 1766 684 1818 736
rect 1942 748 1994 800
rect 1942 684 1994 736
rect 2118 748 2170 800
rect 2118 684 2170 736
rect 6 495 58 547
rect 6 431 58 483
rect 182 495 234 547
rect 182 431 234 483
rect 358 495 410 547
rect 358 431 410 483
rect 534 495 586 547
rect 534 431 586 483
rect 710 495 762 547
rect 710 431 762 483
rect 886 495 938 547
rect 886 431 938 483
rect 1062 495 1114 547
rect 1062 431 1114 483
rect 1238 495 1290 547
rect 1238 431 1290 483
rect 1414 495 1466 547
rect 1414 431 1466 483
rect 1590 495 1642 547
rect 1590 431 1642 483
rect 1766 495 1818 547
rect 1766 431 1818 483
rect 1942 495 1994 547
rect 1942 431 1994 483
rect 2118 495 2170 547
rect 2118 431 2170 483
rect 6 247 58 299
rect 6 183 58 235
rect 182 247 234 299
rect 182 183 234 235
rect 358 247 410 299
rect 358 183 410 235
rect 534 247 586 299
rect 534 183 586 235
rect 710 247 762 299
rect 710 183 762 235
rect 886 247 938 299
rect 886 183 938 235
rect 1062 247 1114 299
rect 1062 183 1114 235
rect 1238 247 1290 299
rect 1238 183 1290 235
rect 1414 247 1466 299
rect 1414 183 1466 235
rect 1590 247 1642 299
rect 1590 183 1642 235
rect 1766 247 1818 299
rect 1766 183 1818 235
rect 1942 247 1994 299
rect 1942 183 1994 235
rect 2118 247 2170 299
rect 2118 183 2170 235
rect 91 -85 100 -55
rect 100 -85 134 -55
rect 134 -85 143 -55
rect 91 -107 143 -85
rect 91 -123 143 -119
rect 91 -157 100 -123
rect 100 -157 134 -123
rect 134 -157 143 -123
rect 91 -171 143 -157
rect 267 -85 276 -55
rect 276 -85 310 -55
rect 310 -85 319 -55
rect 267 -107 319 -85
rect 267 -123 319 -119
rect 267 -157 276 -123
rect 276 -157 310 -123
rect 310 -157 319 -123
rect 267 -171 319 -157
rect 91 -339 143 -305
rect 91 -357 100 -339
rect 100 -357 134 -339
rect 134 -357 143 -339
rect 91 -373 100 -369
rect 100 -373 134 -369
rect 134 -373 143 -369
rect 91 -411 143 -373
rect 91 -421 100 -411
rect 100 -421 134 -411
rect 134 -421 143 -411
rect 443 -85 452 -55
rect 452 -85 486 -55
rect 486 -85 495 -55
rect 443 -107 495 -85
rect 443 -123 495 -119
rect 443 -157 452 -123
rect 452 -157 486 -123
rect 486 -157 495 -123
rect 443 -171 495 -157
rect 267 -339 319 -305
rect 267 -357 276 -339
rect 276 -357 310 -339
rect 310 -357 319 -339
rect 267 -373 276 -369
rect 276 -373 310 -369
rect 310 -373 319 -369
rect 267 -411 319 -373
rect 267 -421 276 -411
rect 276 -421 310 -411
rect 310 -421 319 -411
rect 91 -589 100 -555
rect 100 -589 134 -555
rect 134 -589 143 -555
rect 91 -607 143 -589
rect 91 -627 143 -619
rect 91 -661 100 -627
rect 100 -661 134 -627
rect 134 -661 143 -627
rect 91 -671 143 -661
rect 619 -85 628 -55
rect 628 -85 662 -55
rect 662 -85 671 -55
rect 619 -107 671 -85
rect 619 -123 671 -119
rect 619 -157 628 -123
rect 628 -157 662 -123
rect 662 -157 671 -123
rect 619 -171 671 -157
rect 443 -339 495 -305
rect 443 -357 452 -339
rect 452 -357 486 -339
rect 486 -357 495 -339
rect 443 -373 452 -369
rect 452 -373 486 -369
rect 486 -373 495 -369
rect 443 -411 495 -373
rect 443 -421 452 -411
rect 452 -421 486 -411
rect 486 -421 495 -411
rect 267 -589 276 -555
rect 276 -589 310 -555
rect 310 -589 319 -555
rect 267 -607 319 -589
rect 267 -627 319 -619
rect 267 -661 276 -627
rect 276 -661 310 -627
rect 310 -661 319 -627
rect 267 -671 319 -661
rect 795 -85 804 -55
rect 804 -85 838 -55
rect 838 -85 847 -55
rect 795 -107 847 -85
rect 795 -123 847 -119
rect 795 -157 804 -123
rect 804 -157 838 -123
rect 838 -157 847 -123
rect 795 -171 847 -157
rect 619 -339 671 -305
rect 619 -357 628 -339
rect 628 -357 662 -339
rect 662 -357 671 -339
rect 619 -373 628 -369
rect 628 -373 662 -369
rect 662 -373 671 -369
rect 619 -411 671 -373
rect 619 -421 628 -411
rect 628 -421 662 -411
rect 662 -421 671 -411
rect 443 -589 452 -555
rect 452 -589 486 -555
rect 486 -589 495 -555
rect 443 -607 495 -589
rect 443 -627 495 -619
rect 443 -661 452 -627
rect 452 -661 486 -627
rect 486 -661 495 -627
rect 443 -671 495 -661
rect 971 -85 980 -55
rect 980 -85 1014 -55
rect 1014 -85 1023 -55
rect 971 -107 1023 -85
rect 971 -123 1023 -119
rect 971 -157 980 -123
rect 980 -157 1014 -123
rect 1014 -157 1023 -123
rect 971 -171 1023 -157
rect 795 -339 847 -305
rect 795 -357 804 -339
rect 804 -357 838 -339
rect 838 -357 847 -339
rect 795 -373 804 -369
rect 804 -373 838 -369
rect 838 -373 847 -369
rect 795 -411 847 -373
rect 795 -421 804 -411
rect 804 -421 838 -411
rect 838 -421 847 -411
rect 619 -589 628 -555
rect 628 -589 662 -555
rect 662 -589 671 -555
rect 619 -607 671 -589
rect 619 -627 671 -619
rect 619 -661 628 -627
rect 628 -661 662 -627
rect 662 -661 671 -627
rect 619 -671 671 -661
rect 1147 -85 1156 -55
rect 1156 -85 1190 -55
rect 1190 -85 1199 -55
rect 1147 -107 1199 -85
rect 1147 -123 1199 -119
rect 1147 -157 1156 -123
rect 1156 -157 1190 -123
rect 1190 -157 1199 -123
rect 1147 -171 1199 -157
rect 971 -339 1023 -305
rect 971 -357 980 -339
rect 980 -357 1014 -339
rect 1014 -357 1023 -339
rect 971 -373 980 -369
rect 980 -373 1014 -369
rect 1014 -373 1023 -369
rect 971 -411 1023 -373
rect 971 -421 980 -411
rect 980 -421 1014 -411
rect 1014 -421 1023 -411
rect 795 -589 804 -555
rect 804 -589 838 -555
rect 838 -589 847 -555
rect 795 -607 847 -589
rect 795 -627 847 -619
rect 795 -661 804 -627
rect 804 -661 838 -627
rect 838 -661 847 -627
rect 795 -671 847 -661
rect 1323 -85 1332 -55
rect 1332 -85 1366 -55
rect 1366 -85 1375 -55
rect 1323 -107 1375 -85
rect 1323 -123 1375 -119
rect 1323 -157 1332 -123
rect 1332 -157 1366 -123
rect 1366 -157 1375 -123
rect 1323 -171 1375 -157
rect 1147 -339 1199 -305
rect 1147 -357 1156 -339
rect 1156 -357 1190 -339
rect 1190 -357 1199 -339
rect 1147 -373 1156 -369
rect 1156 -373 1190 -369
rect 1190 -373 1199 -369
rect 1147 -411 1199 -373
rect 1147 -421 1156 -411
rect 1156 -421 1190 -411
rect 1190 -421 1199 -411
rect 971 -589 980 -555
rect 980 -589 1014 -555
rect 1014 -589 1023 -555
rect 971 -607 1023 -589
rect 971 -627 1023 -619
rect 971 -661 980 -627
rect 980 -661 1014 -627
rect 1014 -661 1023 -627
rect 971 -671 1023 -661
rect 1499 -85 1508 -55
rect 1508 -85 1542 -55
rect 1542 -85 1551 -55
rect 1499 -107 1551 -85
rect 1499 -123 1551 -119
rect 1499 -157 1508 -123
rect 1508 -157 1542 -123
rect 1542 -157 1551 -123
rect 1499 -171 1551 -157
rect 1323 -339 1375 -305
rect 1323 -357 1332 -339
rect 1332 -357 1366 -339
rect 1366 -357 1375 -339
rect 1323 -373 1332 -369
rect 1332 -373 1366 -369
rect 1366 -373 1375 -369
rect 1323 -411 1375 -373
rect 1323 -421 1332 -411
rect 1332 -421 1366 -411
rect 1366 -421 1375 -411
rect 1147 -589 1156 -555
rect 1156 -589 1190 -555
rect 1190 -589 1199 -555
rect 1147 -607 1199 -589
rect 1147 -627 1199 -619
rect 1147 -661 1156 -627
rect 1156 -661 1190 -627
rect 1190 -661 1199 -627
rect 1147 -671 1199 -661
rect 1675 -85 1684 -55
rect 1684 -85 1718 -55
rect 1718 -85 1727 -55
rect 1675 -107 1727 -85
rect 1675 -123 1727 -119
rect 1675 -157 1684 -123
rect 1684 -157 1718 -123
rect 1718 -157 1727 -123
rect 1675 -171 1727 -157
rect 1499 -339 1551 -305
rect 1499 -357 1508 -339
rect 1508 -357 1542 -339
rect 1542 -357 1551 -339
rect 1499 -373 1508 -369
rect 1508 -373 1542 -369
rect 1542 -373 1551 -369
rect 1499 -411 1551 -373
rect 1499 -421 1508 -411
rect 1508 -421 1542 -411
rect 1542 -421 1551 -411
rect 1323 -589 1332 -555
rect 1332 -589 1366 -555
rect 1366 -589 1375 -555
rect 1323 -607 1375 -589
rect 1323 -627 1375 -619
rect 1323 -661 1332 -627
rect 1332 -661 1366 -627
rect 1366 -661 1375 -627
rect 1323 -671 1375 -661
rect 1851 -85 1860 -55
rect 1860 -85 1894 -55
rect 1894 -85 1903 -55
rect 1851 -107 1903 -85
rect 1851 -123 1903 -119
rect 1851 -157 1860 -123
rect 1860 -157 1894 -123
rect 1894 -157 1903 -123
rect 1851 -171 1903 -157
rect 1675 -339 1727 -305
rect 1675 -357 1684 -339
rect 1684 -357 1718 -339
rect 1718 -357 1727 -339
rect 1675 -373 1684 -369
rect 1684 -373 1718 -369
rect 1718 -373 1727 -369
rect 1675 -411 1727 -373
rect 1675 -421 1684 -411
rect 1684 -421 1718 -411
rect 1718 -421 1727 -411
rect 1499 -589 1508 -555
rect 1508 -589 1542 -555
rect 1542 -589 1551 -555
rect 1499 -607 1551 -589
rect 1499 -627 1551 -619
rect 1499 -661 1508 -627
rect 1508 -661 1542 -627
rect 1542 -661 1551 -627
rect 1499 -671 1551 -661
rect 2027 -85 2036 -55
rect 2036 -85 2070 -55
rect 2070 -85 2079 -55
rect 2027 -107 2079 -85
rect 2027 -123 2079 -119
rect 2027 -157 2036 -123
rect 2036 -157 2070 -123
rect 2070 -157 2079 -123
rect 2027 -171 2079 -157
rect 1851 -339 1903 -305
rect 1851 -357 1860 -339
rect 1860 -357 1894 -339
rect 1894 -357 1903 -339
rect 1851 -373 1860 -369
rect 1860 -373 1894 -369
rect 1894 -373 1903 -369
rect 1851 -411 1903 -373
rect 1851 -421 1860 -411
rect 1860 -421 1894 -411
rect 1894 -421 1903 -411
rect 1675 -589 1684 -555
rect 1684 -589 1718 -555
rect 1718 -589 1727 -555
rect 1675 -607 1727 -589
rect 1675 -627 1727 -619
rect 1675 -661 1684 -627
rect 1684 -661 1718 -627
rect 1718 -661 1727 -627
rect 1675 -671 1727 -661
rect 2203 -85 2212 -55
rect 2212 -85 2246 -55
rect 2246 -85 2255 -55
rect 2203 -107 2255 -85
rect 2203 -123 2255 -119
rect 2203 -157 2212 -123
rect 2212 -157 2246 -123
rect 2246 -157 2255 -123
rect 2203 -171 2255 -157
rect 2027 -339 2079 -305
rect 2027 -357 2036 -339
rect 2036 -357 2070 -339
rect 2070 -357 2079 -339
rect 2027 -373 2036 -369
rect 2036 -373 2070 -369
rect 2070 -373 2079 -369
rect 2027 -411 2079 -373
rect 2027 -421 2036 -411
rect 2036 -421 2070 -411
rect 2070 -421 2079 -411
rect 1851 -589 1860 -555
rect 1860 -589 1894 -555
rect 1894 -589 1903 -555
rect 1851 -607 1903 -589
rect 1851 -627 1903 -619
rect 1851 -661 1860 -627
rect 1860 -661 1894 -627
rect 1894 -661 1903 -627
rect 1851 -671 1903 -661
rect 2203 -339 2255 -305
rect 2203 -357 2212 -339
rect 2212 -357 2246 -339
rect 2246 -357 2255 -339
rect 2203 -373 2212 -369
rect 2212 -373 2246 -369
rect 2246 -373 2255 -369
rect 2203 -411 2255 -373
rect 2203 -421 2212 -411
rect 2212 -421 2246 -411
rect 2246 -421 2255 -411
rect 2027 -589 2036 -555
rect 2036 -589 2070 -555
rect 2070 -589 2079 -555
rect 2027 -607 2079 -589
rect 2027 -627 2079 -619
rect 2027 -661 2036 -627
rect 2036 -661 2070 -627
rect 2070 -661 2079 -627
rect 2027 -671 2079 -661
rect 2203 -589 2212 -555
rect 2212 -589 2246 -555
rect 2246 -589 2255 -555
rect 2203 -607 2255 -589
rect 2203 -627 2255 -619
rect 2203 -661 2212 -627
rect 2212 -661 2246 -627
rect 2246 -661 2255 -627
rect 2203 -671 2255 -661
<< metal2 >>
rect 56 1299 2201 1403
rect 56 991 177 1299
rect 2085 991 2201 1299
rect 56 864 2201 991
rect 0 800 2246 814
rect 0 748 6 800
rect 58 748 182 800
rect 234 748 358 800
rect 410 748 534 800
rect 586 748 710 800
rect 762 748 886 800
rect 938 748 1062 800
rect 1114 748 1238 800
rect 1290 748 1414 800
rect 1466 748 1590 800
rect 1642 748 1766 800
rect 1818 748 1942 800
rect 1994 748 2118 800
rect 2170 748 2246 800
rect 0 736 2246 748
rect 0 684 6 736
rect 58 684 182 736
rect 234 684 358 736
rect 410 684 534 736
rect 586 684 710 736
rect 762 684 886 736
rect 938 684 1062 736
rect 1114 684 1238 736
rect 1290 684 1414 736
rect 1466 684 1590 736
rect 1642 684 1766 736
rect 1818 684 1942 736
rect 1994 684 2118 736
rect 2170 684 2246 736
rect 0 674 2246 684
rect 12 667 2246 674
rect 0 547 2867 627
rect 0 495 6 547
rect 58 495 182 547
rect 234 495 358 547
rect 410 495 534 547
rect 586 495 710 547
rect 762 495 886 547
rect 938 495 1062 547
rect 1114 495 1238 547
rect 1290 495 1414 547
rect 1466 495 1590 547
rect 1642 495 1766 547
rect 1818 495 1942 547
rect 1994 495 2118 547
rect 2170 495 2867 547
rect 0 483 2867 495
rect 0 431 6 483
rect 58 431 182 483
rect 234 431 358 483
rect 410 431 534 483
rect 586 431 710 483
rect 762 431 886 483
rect 938 431 1062 483
rect 1114 431 1238 483
rect 1290 431 1414 483
rect 1466 431 1590 483
rect 1642 431 1766 483
rect 1818 431 1942 483
rect 1994 431 2118 483
rect 2170 431 2867 483
rect 0 299 2867 431
rect 0 247 6 299
rect 58 247 182 299
rect 234 247 358 299
rect 410 247 534 299
rect 586 247 710 299
rect 762 247 886 299
rect 938 247 1062 299
rect 1114 247 1238 299
rect 1290 247 1414 299
rect 1466 247 1590 299
rect 1642 247 1766 299
rect 1818 247 1942 299
rect 1994 247 2118 299
rect 2170 247 2867 299
rect 0 235 2867 247
rect 0 183 6 235
rect 58 183 182 235
rect 234 183 358 235
rect 410 183 534 235
rect 586 183 710 235
rect 762 183 886 235
rect 938 183 1062 235
rect 1114 183 1238 235
rect 1290 183 1414 235
rect 1466 183 1590 235
rect 1642 183 1766 235
rect 1818 183 1942 235
rect 1994 183 2118 235
rect 2170 183 2867 235
rect 0 172 2867 183
rect 12 167 2246 172
rect -641 -55 2261 -39
rect -641 -107 91 -55
rect 143 -107 267 -55
rect 319 -107 443 -55
rect 495 -107 619 -55
rect 671 -107 795 -55
rect 847 -107 971 -55
rect 1023 -107 1147 -55
rect 1199 -107 1323 -55
rect 1375 -107 1499 -55
rect 1551 -107 1675 -55
rect 1727 -107 1851 -55
rect 1903 -107 2027 -55
rect 2079 -107 2203 -55
rect 2255 -107 2261 -55
rect -641 -119 2261 -107
rect -641 -171 91 -119
rect 143 -171 267 -119
rect 319 -171 443 -119
rect 495 -171 619 -119
rect 671 -171 795 -119
rect 847 -171 971 -119
rect 1023 -171 1147 -119
rect 1199 -171 1323 -119
rect 1375 -171 1499 -119
rect 1551 -171 1675 -119
rect 1727 -171 1851 -119
rect 1903 -171 2027 -119
rect 2079 -171 2203 -119
rect 2255 -171 2261 -119
rect -641 -305 2261 -171
rect -641 -357 91 -305
rect 143 -357 267 -305
rect 319 -357 443 -305
rect 495 -357 619 -305
rect 671 -357 795 -305
rect 847 -357 971 -305
rect 1023 -357 1147 -305
rect 1199 -357 1323 -305
rect 1375 -357 1499 -305
rect 1551 -357 1675 -305
rect 1727 -357 1851 -305
rect 1903 -357 2027 -305
rect 2079 -357 2203 -305
rect 2255 -357 2261 -305
rect -641 -369 2261 -357
rect -641 -421 91 -369
rect 143 -421 267 -369
rect 319 -421 443 -369
rect 495 -421 619 -369
rect 671 -421 795 -369
rect 847 -421 971 -369
rect 1023 -421 1147 -369
rect 1199 -421 1323 -369
rect 1375 -421 1499 -369
rect 1551 -421 1675 -369
rect 1727 -421 1851 -369
rect 1903 -421 2027 -369
rect 2079 -421 2203 -369
rect 2255 -421 2261 -369
rect -641 -555 2261 -421
rect -641 -607 91 -555
rect 143 -607 267 -555
rect 319 -607 443 -555
rect 495 -607 619 -555
rect 671 -607 795 -555
rect 847 -607 971 -555
rect 1023 -607 1147 -555
rect 1199 -607 1323 -555
rect 1375 -607 1499 -555
rect 1551 -607 1675 -555
rect 1727 -607 1851 -555
rect 1903 -607 2027 -555
rect 2079 -607 2203 -555
rect 2255 -607 2261 -555
rect -641 -619 2261 -607
rect -641 -671 91 -619
rect 143 -671 267 -619
rect 319 -671 443 -619
rect 495 -671 619 -619
rect 671 -671 795 -619
rect 847 -671 971 -619
rect 1023 -671 1147 -619
rect 1199 -671 1323 -619
rect 1375 -671 1499 -619
rect 1551 -671 1675 -619
rect 1727 -671 1851 -619
rect 1903 -671 2027 -619
rect 2079 -671 2203 -619
rect 2255 -671 2261 -619
rect -641 -687 2261 -671
<< via2 >>
rect 183 997 2079 1293
<< metal3 >>
rect 56 1297 2201 1403
rect 56 993 179 1297
rect 2083 993 2201 1297
rect 56 864 2201 993
<< via3 >>
rect 179 1293 2083 1297
rect 179 997 183 1293
rect 183 997 2079 1293
rect 2079 997 2083 1293
rect 179 993 2083 997
<< metal4 >>
rect 56 1297 2201 1403
rect 56 993 179 1297
rect 2083 993 2201 1297
rect 56 864 2201 993
<< via4 >>
rect 213 1027 449 1263
rect 533 1027 769 1263
rect 853 1027 1089 1263
rect 1173 1027 1409 1263
rect 1493 1027 1729 1263
rect 1813 1027 2049 1263
<< metal5 >>
rect 57 1263 2201 2330
rect 57 1027 213 1263
rect 449 1027 533 1263
rect 769 1027 853 1263
rect 1089 1027 1173 1263
rect 1409 1027 1493 1263
rect 1729 1027 1813 1263
rect 2049 1027 2201 1263
rect 57 863 2201 1027
use sky130_fd_pr__res_xhigh_po_0p35_9FS993  sky130_fd_pr__res_xhigh_po_0p35_9FS993_0
timestamp 1636132012
transform 0 1 4870 -1 0 -947
box -191 -2088 191 2088
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_24
timestamp 1636132012
transform 1 0 73 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_23
timestamp 1636132012
transform 1 0 161 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_22
timestamp 1636132012
transform 1 0 249 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_21
timestamp 1636132012
transform 1 0 337 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_20
timestamp 1636132012
transform 1 0 425 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_19
timestamp 1636132012
transform 1 0 513 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_18
timestamp 1636132012
transform 1 0 601 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_17
timestamp 1636132012
transform 1 0 689 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_16
timestamp 1636132012
transform 1 0 777 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_15
timestamp 1636132012
transform 1 0 865 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_14
timestamp 1636132012
transform 1 0 953 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_13
timestamp 1636132012
transform 1 0 1129 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_12
timestamp 1636132012
transform 1 0 1041 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_11
timestamp 1636132012
transform 1 0 1217 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_10
timestamp 1636132012
transform 1 0 1305 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_9
timestamp 1636132012
transform 1 0 1481 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_8
timestamp 1636132012
transform 1 0 1393 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_7
timestamp 1636132012
transform 1 0 1657 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_6
timestamp 1636132012
transform 1 0 1569 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_5
timestamp 1636132012
transform 1 0 1745 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_4
timestamp 1636132012
transform 1 0 1833 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_3
timestamp 1636132012
transform 1 0 2009 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_2
timestamp 1636132012
transform 1 0 1921 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_1
timestamp 1636132012
transform 1 0 2097 0 1 426
box -99 -426 99 426
use sky130_fd_pr__nfet_01v8_lvt_BG9PLE  sky130_fd_pr__nfet_01v8_lvt_BG9PLE_0
timestamp 1636132012
transform 1 0 2185 0 1 426
box -99 -426 99 426
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1636132012
transform 1 0 3050 0 1 5035
box -3351 -3101 3373 3101
<< end >>
