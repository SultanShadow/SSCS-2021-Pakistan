magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< pwell >>
rect 2689 2588 2814 2589
rect -1711 2431 2814 2588
rect -1711 2282 -1586 2431
rect -5952 2196 -1586 2282
rect -5952 1986 -5866 2196
rect -1862 2132 -1586 2196
rect -1862 1986 392 2132
rect -5952 1773 392 1986
rect -5957 1687 392 1773
rect -5957 1477 -5871 1687
rect -1867 1477 392 1687
rect -5957 1234 392 1477
rect -5996 1148 392 1234
rect -5996 938 -5910 1148
rect -1906 938 392 1148
rect -5996 880 392 938
rect -5996 852 -1586 880
rect -1711 463 -1586 852
rect 2689 463 2814 2431
rect -1711 306 2814 463
<< nmoslvt >>
rect -1394 906 -1364 2106
rect -1306 906 -1276 2106
rect -1218 906 -1188 2106
rect -1130 906 -1100 2106
rect -1042 906 -1012 2106
rect -954 906 -924 2106
rect -866 906 -836 2106
rect -778 906 -748 2106
rect -690 906 -660 2106
rect -602 906 -572 2106
rect -514 906 -484 2106
rect -426 906 -396 2106
rect -338 906 -308 2106
rect -250 906 -220 2106
rect -162 906 -132 2106
rect -74 906 -44 2106
rect 14 906 44 2106
rect 102 906 132 2106
rect 190 906 220 2106
rect 278 906 308 2106
<< ndiff >>
rect -1452 2067 -1394 2106
rect -1452 2033 -1440 2067
rect -1406 2033 -1394 2067
rect -1452 1999 -1394 2033
rect -1452 1965 -1440 1999
rect -1406 1965 -1394 1999
rect -1452 1931 -1394 1965
rect -1452 1897 -1440 1931
rect -1406 1897 -1394 1931
rect -1452 1863 -1394 1897
rect -1452 1829 -1440 1863
rect -1406 1829 -1394 1863
rect -1452 1795 -1394 1829
rect -1452 1761 -1440 1795
rect -1406 1761 -1394 1795
rect -1452 1727 -1394 1761
rect -1452 1693 -1440 1727
rect -1406 1693 -1394 1727
rect -1452 1659 -1394 1693
rect -1452 1625 -1440 1659
rect -1406 1625 -1394 1659
rect -1452 1591 -1394 1625
rect -1452 1557 -1440 1591
rect -1406 1557 -1394 1591
rect -1452 1523 -1394 1557
rect -1452 1489 -1440 1523
rect -1406 1489 -1394 1523
rect -1452 1455 -1394 1489
rect -1452 1421 -1440 1455
rect -1406 1421 -1394 1455
rect -1452 1387 -1394 1421
rect -1452 1353 -1440 1387
rect -1406 1353 -1394 1387
rect -1452 1319 -1394 1353
rect -1452 1285 -1440 1319
rect -1406 1285 -1394 1319
rect -1452 1251 -1394 1285
rect -1452 1217 -1440 1251
rect -1406 1217 -1394 1251
rect -1452 1183 -1394 1217
rect -1452 1149 -1440 1183
rect -1406 1149 -1394 1183
rect -1452 1115 -1394 1149
rect -1452 1081 -1440 1115
rect -1406 1081 -1394 1115
rect -1452 1047 -1394 1081
rect -1452 1013 -1440 1047
rect -1406 1013 -1394 1047
rect -1452 979 -1394 1013
rect -1452 945 -1440 979
rect -1406 945 -1394 979
rect -1452 906 -1394 945
rect -1364 2067 -1306 2106
rect -1364 2033 -1352 2067
rect -1318 2033 -1306 2067
rect -1364 1999 -1306 2033
rect -1364 1965 -1352 1999
rect -1318 1965 -1306 1999
rect -1364 1931 -1306 1965
rect -1364 1897 -1352 1931
rect -1318 1897 -1306 1931
rect -1364 1863 -1306 1897
rect -1364 1829 -1352 1863
rect -1318 1829 -1306 1863
rect -1364 1795 -1306 1829
rect -1364 1761 -1352 1795
rect -1318 1761 -1306 1795
rect -1364 1727 -1306 1761
rect -1364 1693 -1352 1727
rect -1318 1693 -1306 1727
rect -1364 1659 -1306 1693
rect -1364 1625 -1352 1659
rect -1318 1625 -1306 1659
rect -1364 1591 -1306 1625
rect -1364 1557 -1352 1591
rect -1318 1557 -1306 1591
rect -1364 1523 -1306 1557
rect -1364 1489 -1352 1523
rect -1318 1489 -1306 1523
rect -1364 1455 -1306 1489
rect -1364 1421 -1352 1455
rect -1318 1421 -1306 1455
rect -1364 1387 -1306 1421
rect -1364 1353 -1352 1387
rect -1318 1353 -1306 1387
rect -1364 1319 -1306 1353
rect -1364 1285 -1352 1319
rect -1318 1285 -1306 1319
rect -1364 1251 -1306 1285
rect -1364 1217 -1352 1251
rect -1318 1217 -1306 1251
rect -1364 1183 -1306 1217
rect -1364 1149 -1352 1183
rect -1318 1149 -1306 1183
rect -1364 1115 -1306 1149
rect -1364 1081 -1352 1115
rect -1318 1081 -1306 1115
rect -1364 1047 -1306 1081
rect -1364 1013 -1352 1047
rect -1318 1013 -1306 1047
rect -1364 979 -1306 1013
rect -1364 945 -1352 979
rect -1318 945 -1306 979
rect -1364 906 -1306 945
rect -1276 2067 -1218 2106
rect -1276 2033 -1264 2067
rect -1230 2033 -1218 2067
rect -1276 1999 -1218 2033
rect -1276 1965 -1264 1999
rect -1230 1965 -1218 1999
rect -1276 1931 -1218 1965
rect -1276 1897 -1264 1931
rect -1230 1897 -1218 1931
rect -1276 1863 -1218 1897
rect -1276 1829 -1264 1863
rect -1230 1829 -1218 1863
rect -1276 1795 -1218 1829
rect -1276 1761 -1264 1795
rect -1230 1761 -1218 1795
rect -1276 1727 -1218 1761
rect -1276 1693 -1264 1727
rect -1230 1693 -1218 1727
rect -1276 1659 -1218 1693
rect -1276 1625 -1264 1659
rect -1230 1625 -1218 1659
rect -1276 1591 -1218 1625
rect -1276 1557 -1264 1591
rect -1230 1557 -1218 1591
rect -1276 1523 -1218 1557
rect -1276 1489 -1264 1523
rect -1230 1489 -1218 1523
rect -1276 1455 -1218 1489
rect -1276 1421 -1264 1455
rect -1230 1421 -1218 1455
rect -1276 1387 -1218 1421
rect -1276 1353 -1264 1387
rect -1230 1353 -1218 1387
rect -1276 1319 -1218 1353
rect -1276 1285 -1264 1319
rect -1230 1285 -1218 1319
rect -1276 1251 -1218 1285
rect -1276 1217 -1264 1251
rect -1230 1217 -1218 1251
rect -1276 1183 -1218 1217
rect -1276 1149 -1264 1183
rect -1230 1149 -1218 1183
rect -1276 1115 -1218 1149
rect -1276 1081 -1264 1115
rect -1230 1081 -1218 1115
rect -1276 1047 -1218 1081
rect -1276 1013 -1264 1047
rect -1230 1013 -1218 1047
rect -1276 979 -1218 1013
rect -1276 945 -1264 979
rect -1230 945 -1218 979
rect -1276 906 -1218 945
rect -1188 2067 -1130 2106
rect -1188 2033 -1176 2067
rect -1142 2033 -1130 2067
rect -1188 1999 -1130 2033
rect -1188 1965 -1176 1999
rect -1142 1965 -1130 1999
rect -1188 1931 -1130 1965
rect -1188 1897 -1176 1931
rect -1142 1897 -1130 1931
rect -1188 1863 -1130 1897
rect -1188 1829 -1176 1863
rect -1142 1829 -1130 1863
rect -1188 1795 -1130 1829
rect -1188 1761 -1176 1795
rect -1142 1761 -1130 1795
rect -1188 1727 -1130 1761
rect -1188 1693 -1176 1727
rect -1142 1693 -1130 1727
rect -1188 1659 -1130 1693
rect -1188 1625 -1176 1659
rect -1142 1625 -1130 1659
rect -1188 1591 -1130 1625
rect -1188 1557 -1176 1591
rect -1142 1557 -1130 1591
rect -1188 1523 -1130 1557
rect -1188 1489 -1176 1523
rect -1142 1489 -1130 1523
rect -1188 1455 -1130 1489
rect -1188 1421 -1176 1455
rect -1142 1421 -1130 1455
rect -1188 1387 -1130 1421
rect -1188 1353 -1176 1387
rect -1142 1353 -1130 1387
rect -1188 1319 -1130 1353
rect -1188 1285 -1176 1319
rect -1142 1285 -1130 1319
rect -1188 1251 -1130 1285
rect -1188 1217 -1176 1251
rect -1142 1217 -1130 1251
rect -1188 1183 -1130 1217
rect -1188 1149 -1176 1183
rect -1142 1149 -1130 1183
rect -1188 1115 -1130 1149
rect -1188 1081 -1176 1115
rect -1142 1081 -1130 1115
rect -1188 1047 -1130 1081
rect -1188 1013 -1176 1047
rect -1142 1013 -1130 1047
rect -1188 979 -1130 1013
rect -1188 945 -1176 979
rect -1142 945 -1130 979
rect -1188 906 -1130 945
rect -1100 2067 -1042 2106
rect -1100 2033 -1088 2067
rect -1054 2033 -1042 2067
rect -1100 1999 -1042 2033
rect -1100 1965 -1088 1999
rect -1054 1965 -1042 1999
rect -1100 1931 -1042 1965
rect -1100 1897 -1088 1931
rect -1054 1897 -1042 1931
rect -1100 1863 -1042 1897
rect -1100 1829 -1088 1863
rect -1054 1829 -1042 1863
rect -1100 1795 -1042 1829
rect -1100 1761 -1088 1795
rect -1054 1761 -1042 1795
rect -1100 1727 -1042 1761
rect -1100 1693 -1088 1727
rect -1054 1693 -1042 1727
rect -1100 1659 -1042 1693
rect -1100 1625 -1088 1659
rect -1054 1625 -1042 1659
rect -1100 1591 -1042 1625
rect -1100 1557 -1088 1591
rect -1054 1557 -1042 1591
rect -1100 1523 -1042 1557
rect -1100 1489 -1088 1523
rect -1054 1489 -1042 1523
rect -1100 1455 -1042 1489
rect -1100 1421 -1088 1455
rect -1054 1421 -1042 1455
rect -1100 1387 -1042 1421
rect -1100 1353 -1088 1387
rect -1054 1353 -1042 1387
rect -1100 1319 -1042 1353
rect -1100 1285 -1088 1319
rect -1054 1285 -1042 1319
rect -1100 1251 -1042 1285
rect -1100 1217 -1088 1251
rect -1054 1217 -1042 1251
rect -1100 1183 -1042 1217
rect -1100 1149 -1088 1183
rect -1054 1149 -1042 1183
rect -1100 1115 -1042 1149
rect -1100 1081 -1088 1115
rect -1054 1081 -1042 1115
rect -1100 1047 -1042 1081
rect -1100 1013 -1088 1047
rect -1054 1013 -1042 1047
rect -1100 979 -1042 1013
rect -1100 945 -1088 979
rect -1054 945 -1042 979
rect -1100 906 -1042 945
rect -1012 2067 -954 2106
rect -1012 2033 -1000 2067
rect -966 2033 -954 2067
rect -1012 1999 -954 2033
rect -1012 1965 -1000 1999
rect -966 1965 -954 1999
rect -1012 1931 -954 1965
rect -1012 1897 -1000 1931
rect -966 1897 -954 1931
rect -1012 1863 -954 1897
rect -1012 1829 -1000 1863
rect -966 1829 -954 1863
rect -1012 1795 -954 1829
rect -1012 1761 -1000 1795
rect -966 1761 -954 1795
rect -1012 1727 -954 1761
rect -1012 1693 -1000 1727
rect -966 1693 -954 1727
rect -1012 1659 -954 1693
rect -1012 1625 -1000 1659
rect -966 1625 -954 1659
rect -1012 1591 -954 1625
rect -1012 1557 -1000 1591
rect -966 1557 -954 1591
rect -1012 1523 -954 1557
rect -1012 1489 -1000 1523
rect -966 1489 -954 1523
rect -1012 1455 -954 1489
rect -1012 1421 -1000 1455
rect -966 1421 -954 1455
rect -1012 1387 -954 1421
rect -1012 1353 -1000 1387
rect -966 1353 -954 1387
rect -1012 1319 -954 1353
rect -1012 1285 -1000 1319
rect -966 1285 -954 1319
rect -1012 1251 -954 1285
rect -1012 1217 -1000 1251
rect -966 1217 -954 1251
rect -1012 1183 -954 1217
rect -1012 1149 -1000 1183
rect -966 1149 -954 1183
rect -1012 1115 -954 1149
rect -1012 1081 -1000 1115
rect -966 1081 -954 1115
rect -1012 1047 -954 1081
rect -1012 1013 -1000 1047
rect -966 1013 -954 1047
rect -1012 979 -954 1013
rect -1012 945 -1000 979
rect -966 945 -954 979
rect -1012 906 -954 945
rect -924 2067 -866 2106
rect -924 2033 -912 2067
rect -878 2033 -866 2067
rect -924 1999 -866 2033
rect -924 1965 -912 1999
rect -878 1965 -866 1999
rect -924 1931 -866 1965
rect -924 1897 -912 1931
rect -878 1897 -866 1931
rect -924 1863 -866 1897
rect -924 1829 -912 1863
rect -878 1829 -866 1863
rect -924 1795 -866 1829
rect -924 1761 -912 1795
rect -878 1761 -866 1795
rect -924 1727 -866 1761
rect -924 1693 -912 1727
rect -878 1693 -866 1727
rect -924 1659 -866 1693
rect -924 1625 -912 1659
rect -878 1625 -866 1659
rect -924 1591 -866 1625
rect -924 1557 -912 1591
rect -878 1557 -866 1591
rect -924 1523 -866 1557
rect -924 1489 -912 1523
rect -878 1489 -866 1523
rect -924 1455 -866 1489
rect -924 1421 -912 1455
rect -878 1421 -866 1455
rect -924 1387 -866 1421
rect -924 1353 -912 1387
rect -878 1353 -866 1387
rect -924 1319 -866 1353
rect -924 1285 -912 1319
rect -878 1285 -866 1319
rect -924 1251 -866 1285
rect -924 1217 -912 1251
rect -878 1217 -866 1251
rect -924 1183 -866 1217
rect -924 1149 -912 1183
rect -878 1149 -866 1183
rect -924 1115 -866 1149
rect -924 1081 -912 1115
rect -878 1081 -866 1115
rect -924 1047 -866 1081
rect -924 1013 -912 1047
rect -878 1013 -866 1047
rect -924 979 -866 1013
rect -924 945 -912 979
rect -878 945 -866 979
rect -924 906 -866 945
rect -836 2067 -778 2106
rect -836 2033 -824 2067
rect -790 2033 -778 2067
rect -836 1999 -778 2033
rect -836 1965 -824 1999
rect -790 1965 -778 1999
rect -836 1931 -778 1965
rect -836 1897 -824 1931
rect -790 1897 -778 1931
rect -836 1863 -778 1897
rect -836 1829 -824 1863
rect -790 1829 -778 1863
rect -836 1795 -778 1829
rect -836 1761 -824 1795
rect -790 1761 -778 1795
rect -836 1727 -778 1761
rect -836 1693 -824 1727
rect -790 1693 -778 1727
rect -836 1659 -778 1693
rect -836 1625 -824 1659
rect -790 1625 -778 1659
rect -836 1591 -778 1625
rect -836 1557 -824 1591
rect -790 1557 -778 1591
rect -836 1523 -778 1557
rect -836 1489 -824 1523
rect -790 1489 -778 1523
rect -836 1455 -778 1489
rect -836 1421 -824 1455
rect -790 1421 -778 1455
rect -836 1387 -778 1421
rect -836 1353 -824 1387
rect -790 1353 -778 1387
rect -836 1319 -778 1353
rect -836 1285 -824 1319
rect -790 1285 -778 1319
rect -836 1251 -778 1285
rect -836 1217 -824 1251
rect -790 1217 -778 1251
rect -836 1183 -778 1217
rect -836 1149 -824 1183
rect -790 1149 -778 1183
rect -836 1115 -778 1149
rect -836 1081 -824 1115
rect -790 1081 -778 1115
rect -836 1047 -778 1081
rect -836 1013 -824 1047
rect -790 1013 -778 1047
rect -836 979 -778 1013
rect -836 945 -824 979
rect -790 945 -778 979
rect -836 906 -778 945
rect -748 2067 -690 2106
rect -748 2033 -736 2067
rect -702 2033 -690 2067
rect -748 1999 -690 2033
rect -748 1965 -736 1999
rect -702 1965 -690 1999
rect -748 1931 -690 1965
rect -748 1897 -736 1931
rect -702 1897 -690 1931
rect -748 1863 -690 1897
rect -748 1829 -736 1863
rect -702 1829 -690 1863
rect -748 1795 -690 1829
rect -748 1761 -736 1795
rect -702 1761 -690 1795
rect -748 1727 -690 1761
rect -748 1693 -736 1727
rect -702 1693 -690 1727
rect -748 1659 -690 1693
rect -748 1625 -736 1659
rect -702 1625 -690 1659
rect -748 1591 -690 1625
rect -748 1557 -736 1591
rect -702 1557 -690 1591
rect -748 1523 -690 1557
rect -748 1489 -736 1523
rect -702 1489 -690 1523
rect -748 1455 -690 1489
rect -748 1421 -736 1455
rect -702 1421 -690 1455
rect -748 1387 -690 1421
rect -748 1353 -736 1387
rect -702 1353 -690 1387
rect -748 1319 -690 1353
rect -748 1285 -736 1319
rect -702 1285 -690 1319
rect -748 1251 -690 1285
rect -748 1217 -736 1251
rect -702 1217 -690 1251
rect -748 1183 -690 1217
rect -748 1149 -736 1183
rect -702 1149 -690 1183
rect -748 1115 -690 1149
rect -748 1081 -736 1115
rect -702 1081 -690 1115
rect -748 1047 -690 1081
rect -748 1013 -736 1047
rect -702 1013 -690 1047
rect -748 979 -690 1013
rect -748 945 -736 979
rect -702 945 -690 979
rect -748 906 -690 945
rect -660 2067 -602 2106
rect -660 2033 -648 2067
rect -614 2033 -602 2067
rect -660 1999 -602 2033
rect -660 1965 -648 1999
rect -614 1965 -602 1999
rect -660 1931 -602 1965
rect -660 1897 -648 1931
rect -614 1897 -602 1931
rect -660 1863 -602 1897
rect -660 1829 -648 1863
rect -614 1829 -602 1863
rect -660 1795 -602 1829
rect -660 1761 -648 1795
rect -614 1761 -602 1795
rect -660 1727 -602 1761
rect -660 1693 -648 1727
rect -614 1693 -602 1727
rect -660 1659 -602 1693
rect -660 1625 -648 1659
rect -614 1625 -602 1659
rect -660 1591 -602 1625
rect -660 1557 -648 1591
rect -614 1557 -602 1591
rect -660 1523 -602 1557
rect -660 1489 -648 1523
rect -614 1489 -602 1523
rect -660 1455 -602 1489
rect -660 1421 -648 1455
rect -614 1421 -602 1455
rect -660 1387 -602 1421
rect -660 1353 -648 1387
rect -614 1353 -602 1387
rect -660 1319 -602 1353
rect -660 1285 -648 1319
rect -614 1285 -602 1319
rect -660 1251 -602 1285
rect -660 1217 -648 1251
rect -614 1217 -602 1251
rect -660 1183 -602 1217
rect -660 1149 -648 1183
rect -614 1149 -602 1183
rect -660 1115 -602 1149
rect -660 1081 -648 1115
rect -614 1081 -602 1115
rect -660 1047 -602 1081
rect -660 1013 -648 1047
rect -614 1013 -602 1047
rect -660 979 -602 1013
rect -660 945 -648 979
rect -614 945 -602 979
rect -660 906 -602 945
rect -572 2067 -514 2106
rect -572 2033 -560 2067
rect -526 2033 -514 2067
rect -572 1999 -514 2033
rect -572 1965 -560 1999
rect -526 1965 -514 1999
rect -572 1931 -514 1965
rect -572 1897 -560 1931
rect -526 1897 -514 1931
rect -572 1863 -514 1897
rect -572 1829 -560 1863
rect -526 1829 -514 1863
rect -572 1795 -514 1829
rect -572 1761 -560 1795
rect -526 1761 -514 1795
rect -572 1727 -514 1761
rect -572 1693 -560 1727
rect -526 1693 -514 1727
rect -572 1659 -514 1693
rect -572 1625 -560 1659
rect -526 1625 -514 1659
rect -572 1591 -514 1625
rect -572 1557 -560 1591
rect -526 1557 -514 1591
rect -572 1523 -514 1557
rect -572 1489 -560 1523
rect -526 1489 -514 1523
rect -572 1455 -514 1489
rect -572 1421 -560 1455
rect -526 1421 -514 1455
rect -572 1387 -514 1421
rect -572 1353 -560 1387
rect -526 1353 -514 1387
rect -572 1319 -514 1353
rect -572 1285 -560 1319
rect -526 1285 -514 1319
rect -572 1251 -514 1285
rect -572 1217 -560 1251
rect -526 1217 -514 1251
rect -572 1183 -514 1217
rect -572 1149 -560 1183
rect -526 1149 -514 1183
rect -572 1115 -514 1149
rect -572 1081 -560 1115
rect -526 1081 -514 1115
rect -572 1047 -514 1081
rect -572 1013 -560 1047
rect -526 1013 -514 1047
rect -572 979 -514 1013
rect -572 945 -560 979
rect -526 945 -514 979
rect -572 906 -514 945
rect -484 2067 -426 2106
rect -484 2033 -472 2067
rect -438 2033 -426 2067
rect -484 1999 -426 2033
rect -484 1965 -472 1999
rect -438 1965 -426 1999
rect -484 1931 -426 1965
rect -484 1897 -472 1931
rect -438 1897 -426 1931
rect -484 1863 -426 1897
rect -484 1829 -472 1863
rect -438 1829 -426 1863
rect -484 1795 -426 1829
rect -484 1761 -472 1795
rect -438 1761 -426 1795
rect -484 1727 -426 1761
rect -484 1693 -472 1727
rect -438 1693 -426 1727
rect -484 1659 -426 1693
rect -484 1625 -472 1659
rect -438 1625 -426 1659
rect -484 1591 -426 1625
rect -484 1557 -472 1591
rect -438 1557 -426 1591
rect -484 1523 -426 1557
rect -484 1489 -472 1523
rect -438 1489 -426 1523
rect -484 1455 -426 1489
rect -484 1421 -472 1455
rect -438 1421 -426 1455
rect -484 1387 -426 1421
rect -484 1353 -472 1387
rect -438 1353 -426 1387
rect -484 1319 -426 1353
rect -484 1285 -472 1319
rect -438 1285 -426 1319
rect -484 1251 -426 1285
rect -484 1217 -472 1251
rect -438 1217 -426 1251
rect -484 1183 -426 1217
rect -484 1149 -472 1183
rect -438 1149 -426 1183
rect -484 1115 -426 1149
rect -484 1081 -472 1115
rect -438 1081 -426 1115
rect -484 1047 -426 1081
rect -484 1013 -472 1047
rect -438 1013 -426 1047
rect -484 979 -426 1013
rect -484 945 -472 979
rect -438 945 -426 979
rect -484 906 -426 945
rect -396 2067 -338 2106
rect -396 2033 -384 2067
rect -350 2033 -338 2067
rect -396 1999 -338 2033
rect -396 1965 -384 1999
rect -350 1965 -338 1999
rect -396 1931 -338 1965
rect -396 1897 -384 1931
rect -350 1897 -338 1931
rect -396 1863 -338 1897
rect -396 1829 -384 1863
rect -350 1829 -338 1863
rect -396 1795 -338 1829
rect -396 1761 -384 1795
rect -350 1761 -338 1795
rect -396 1727 -338 1761
rect -396 1693 -384 1727
rect -350 1693 -338 1727
rect -396 1659 -338 1693
rect -396 1625 -384 1659
rect -350 1625 -338 1659
rect -396 1591 -338 1625
rect -396 1557 -384 1591
rect -350 1557 -338 1591
rect -396 1523 -338 1557
rect -396 1489 -384 1523
rect -350 1489 -338 1523
rect -396 1455 -338 1489
rect -396 1421 -384 1455
rect -350 1421 -338 1455
rect -396 1387 -338 1421
rect -396 1353 -384 1387
rect -350 1353 -338 1387
rect -396 1319 -338 1353
rect -396 1285 -384 1319
rect -350 1285 -338 1319
rect -396 1251 -338 1285
rect -396 1217 -384 1251
rect -350 1217 -338 1251
rect -396 1183 -338 1217
rect -396 1149 -384 1183
rect -350 1149 -338 1183
rect -396 1115 -338 1149
rect -396 1081 -384 1115
rect -350 1081 -338 1115
rect -396 1047 -338 1081
rect -396 1013 -384 1047
rect -350 1013 -338 1047
rect -396 979 -338 1013
rect -396 945 -384 979
rect -350 945 -338 979
rect -396 906 -338 945
rect -308 2067 -250 2106
rect -308 2033 -296 2067
rect -262 2033 -250 2067
rect -308 1999 -250 2033
rect -308 1965 -296 1999
rect -262 1965 -250 1999
rect -308 1931 -250 1965
rect -308 1897 -296 1931
rect -262 1897 -250 1931
rect -308 1863 -250 1897
rect -308 1829 -296 1863
rect -262 1829 -250 1863
rect -308 1795 -250 1829
rect -308 1761 -296 1795
rect -262 1761 -250 1795
rect -308 1727 -250 1761
rect -308 1693 -296 1727
rect -262 1693 -250 1727
rect -308 1659 -250 1693
rect -308 1625 -296 1659
rect -262 1625 -250 1659
rect -308 1591 -250 1625
rect -308 1557 -296 1591
rect -262 1557 -250 1591
rect -308 1523 -250 1557
rect -308 1489 -296 1523
rect -262 1489 -250 1523
rect -308 1455 -250 1489
rect -308 1421 -296 1455
rect -262 1421 -250 1455
rect -308 1387 -250 1421
rect -308 1353 -296 1387
rect -262 1353 -250 1387
rect -308 1319 -250 1353
rect -308 1285 -296 1319
rect -262 1285 -250 1319
rect -308 1251 -250 1285
rect -308 1217 -296 1251
rect -262 1217 -250 1251
rect -308 1183 -250 1217
rect -308 1149 -296 1183
rect -262 1149 -250 1183
rect -308 1115 -250 1149
rect -308 1081 -296 1115
rect -262 1081 -250 1115
rect -308 1047 -250 1081
rect -308 1013 -296 1047
rect -262 1013 -250 1047
rect -308 979 -250 1013
rect -308 945 -296 979
rect -262 945 -250 979
rect -308 906 -250 945
rect -220 2067 -162 2106
rect -220 2033 -208 2067
rect -174 2033 -162 2067
rect -220 1999 -162 2033
rect -220 1965 -208 1999
rect -174 1965 -162 1999
rect -220 1931 -162 1965
rect -220 1897 -208 1931
rect -174 1897 -162 1931
rect -220 1863 -162 1897
rect -220 1829 -208 1863
rect -174 1829 -162 1863
rect -220 1795 -162 1829
rect -220 1761 -208 1795
rect -174 1761 -162 1795
rect -220 1727 -162 1761
rect -220 1693 -208 1727
rect -174 1693 -162 1727
rect -220 1659 -162 1693
rect -220 1625 -208 1659
rect -174 1625 -162 1659
rect -220 1591 -162 1625
rect -220 1557 -208 1591
rect -174 1557 -162 1591
rect -220 1523 -162 1557
rect -220 1489 -208 1523
rect -174 1489 -162 1523
rect -220 1455 -162 1489
rect -220 1421 -208 1455
rect -174 1421 -162 1455
rect -220 1387 -162 1421
rect -220 1353 -208 1387
rect -174 1353 -162 1387
rect -220 1319 -162 1353
rect -220 1285 -208 1319
rect -174 1285 -162 1319
rect -220 1251 -162 1285
rect -220 1217 -208 1251
rect -174 1217 -162 1251
rect -220 1183 -162 1217
rect -220 1149 -208 1183
rect -174 1149 -162 1183
rect -220 1115 -162 1149
rect -220 1081 -208 1115
rect -174 1081 -162 1115
rect -220 1047 -162 1081
rect -220 1013 -208 1047
rect -174 1013 -162 1047
rect -220 979 -162 1013
rect -220 945 -208 979
rect -174 945 -162 979
rect -220 906 -162 945
rect -132 2067 -74 2106
rect -132 2033 -120 2067
rect -86 2033 -74 2067
rect -132 1999 -74 2033
rect -132 1965 -120 1999
rect -86 1965 -74 1999
rect -132 1931 -74 1965
rect -132 1897 -120 1931
rect -86 1897 -74 1931
rect -132 1863 -74 1897
rect -132 1829 -120 1863
rect -86 1829 -74 1863
rect -132 1795 -74 1829
rect -132 1761 -120 1795
rect -86 1761 -74 1795
rect -132 1727 -74 1761
rect -132 1693 -120 1727
rect -86 1693 -74 1727
rect -132 1659 -74 1693
rect -132 1625 -120 1659
rect -86 1625 -74 1659
rect -132 1591 -74 1625
rect -132 1557 -120 1591
rect -86 1557 -74 1591
rect -132 1523 -74 1557
rect -132 1489 -120 1523
rect -86 1489 -74 1523
rect -132 1455 -74 1489
rect -132 1421 -120 1455
rect -86 1421 -74 1455
rect -132 1387 -74 1421
rect -132 1353 -120 1387
rect -86 1353 -74 1387
rect -132 1319 -74 1353
rect -132 1285 -120 1319
rect -86 1285 -74 1319
rect -132 1251 -74 1285
rect -132 1217 -120 1251
rect -86 1217 -74 1251
rect -132 1183 -74 1217
rect -132 1149 -120 1183
rect -86 1149 -74 1183
rect -132 1115 -74 1149
rect -132 1081 -120 1115
rect -86 1081 -74 1115
rect -132 1047 -74 1081
rect -132 1013 -120 1047
rect -86 1013 -74 1047
rect -132 979 -74 1013
rect -132 945 -120 979
rect -86 945 -74 979
rect -132 906 -74 945
rect -44 2067 14 2106
rect -44 2033 -32 2067
rect 2 2033 14 2067
rect -44 1999 14 2033
rect -44 1965 -32 1999
rect 2 1965 14 1999
rect -44 1931 14 1965
rect -44 1897 -32 1931
rect 2 1897 14 1931
rect -44 1863 14 1897
rect -44 1829 -32 1863
rect 2 1829 14 1863
rect -44 1795 14 1829
rect -44 1761 -32 1795
rect 2 1761 14 1795
rect -44 1727 14 1761
rect -44 1693 -32 1727
rect 2 1693 14 1727
rect -44 1659 14 1693
rect -44 1625 -32 1659
rect 2 1625 14 1659
rect -44 1591 14 1625
rect -44 1557 -32 1591
rect 2 1557 14 1591
rect -44 1523 14 1557
rect -44 1489 -32 1523
rect 2 1489 14 1523
rect -44 1455 14 1489
rect -44 1421 -32 1455
rect 2 1421 14 1455
rect -44 1387 14 1421
rect -44 1353 -32 1387
rect 2 1353 14 1387
rect -44 1319 14 1353
rect -44 1285 -32 1319
rect 2 1285 14 1319
rect -44 1251 14 1285
rect -44 1217 -32 1251
rect 2 1217 14 1251
rect -44 1183 14 1217
rect -44 1149 -32 1183
rect 2 1149 14 1183
rect -44 1115 14 1149
rect -44 1081 -32 1115
rect 2 1081 14 1115
rect -44 1047 14 1081
rect -44 1013 -32 1047
rect 2 1013 14 1047
rect -44 979 14 1013
rect -44 945 -32 979
rect 2 945 14 979
rect -44 906 14 945
rect 44 2067 102 2106
rect 44 2033 56 2067
rect 90 2033 102 2067
rect 44 1999 102 2033
rect 44 1965 56 1999
rect 90 1965 102 1999
rect 44 1931 102 1965
rect 44 1897 56 1931
rect 90 1897 102 1931
rect 44 1863 102 1897
rect 44 1829 56 1863
rect 90 1829 102 1863
rect 44 1795 102 1829
rect 44 1761 56 1795
rect 90 1761 102 1795
rect 44 1727 102 1761
rect 44 1693 56 1727
rect 90 1693 102 1727
rect 44 1659 102 1693
rect 44 1625 56 1659
rect 90 1625 102 1659
rect 44 1591 102 1625
rect 44 1557 56 1591
rect 90 1557 102 1591
rect 44 1523 102 1557
rect 44 1489 56 1523
rect 90 1489 102 1523
rect 44 1455 102 1489
rect 44 1421 56 1455
rect 90 1421 102 1455
rect 44 1387 102 1421
rect 44 1353 56 1387
rect 90 1353 102 1387
rect 44 1319 102 1353
rect 44 1285 56 1319
rect 90 1285 102 1319
rect 44 1251 102 1285
rect 44 1217 56 1251
rect 90 1217 102 1251
rect 44 1183 102 1217
rect 44 1149 56 1183
rect 90 1149 102 1183
rect 44 1115 102 1149
rect 44 1081 56 1115
rect 90 1081 102 1115
rect 44 1047 102 1081
rect 44 1013 56 1047
rect 90 1013 102 1047
rect 44 979 102 1013
rect 44 945 56 979
rect 90 945 102 979
rect 44 906 102 945
rect 132 2067 190 2106
rect 132 2033 144 2067
rect 178 2033 190 2067
rect 132 1999 190 2033
rect 132 1965 144 1999
rect 178 1965 190 1999
rect 132 1931 190 1965
rect 132 1897 144 1931
rect 178 1897 190 1931
rect 132 1863 190 1897
rect 132 1829 144 1863
rect 178 1829 190 1863
rect 132 1795 190 1829
rect 132 1761 144 1795
rect 178 1761 190 1795
rect 132 1727 190 1761
rect 132 1693 144 1727
rect 178 1693 190 1727
rect 132 1659 190 1693
rect 132 1625 144 1659
rect 178 1625 190 1659
rect 132 1591 190 1625
rect 132 1557 144 1591
rect 178 1557 190 1591
rect 132 1523 190 1557
rect 132 1489 144 1523
rect 178 1489 190 1523
rect 132 1455 190 1489
rect 132 1421 144 1455
rect 178 1421 190 1455
rect 132 1387 190 1421
rect 132 1353 144 1387
rect 178 1353 190 1387
rect 132 1319 190 1353
rect 132 1285 144 1319
rect 178 1285 190 1319
rect 132 1251 190 1285
rect 132 1217 144 1251
rect 178 1217 190 1251
rect 132 1183 190 1217
rect 132 1149 144 1183
rect 178 1149 190 1183
rect 132 1115 190 1149
rect 132 1081 144 1115
rect 178 1081 190 1115
rect 132 1047 190 1081
rect 132 1013 144 1047
rect 178 1013 190 1047
rect 132 979 190 1013
rect 132 945 144 979
rect 178 945 190 979
rect 132 906 190 945
rect 220 2067 278 2106
rect 220 2033 232 2067
rect 266 2033 278 2067
rect 220 1999 278 2033
rect 220 1965 232 1999
rect 266 1965 278 1999
rect 220 1931 278 1965
rect 220 1897 232 1931
rect 266 1897 278 1931
rect 220 1863 278 1897
rect 220 1829 232 1863
rect 266 1829 278 1863
rect 220 1795 278 1829
rect 220 1761 232 1795
rect 266 1761 278 1795
rect 220 1727 278 1761
rect 220 1693 232 1727
rect 266 1693 278 1727
rect 220 1659 278 1693
rect 220 1625 232 1659
rect 266 1625 278 1659
rect 220 1591 278 1625
rect 220 1557 232 1591
rect 266 1557 278 1591
rect 220 1523 278 1557
rect 220 1489 232 1523
rect 266 1489 278 1523
rect 220 1455 278 1489
rect 220 1421 232 1455
rect 266 1421 278 1455
rect 220 1387 278 1421
rect 220 1353 232 1387
rect 266 1353 278 1387
rect 220 1319 278 1353
rect 220 1285 232 1319
rect 266 1285 278 1319
rect 220 1251 278 1285
rect 220 1217 232 1251
rect 266 1217 278 1251
rect 220 1183 278 1217
rect 220 1149 232 1183
rect 266 1149 278 1183
rect 220 1115 278 1149
rect 220 1081 232 1115
rect 266 1081 278 1115
rect 220 1047 278 1081
rect 220 1013 232 1047
rect 266 1013 278 1047
rect 220 979 278 1013
rect 220 945 232 979
rect 266 945 278 979
rect 220 906 278 945
rect 308 2067 366 2106
rect 308 2033 320 2067
rect 354 2033 366 2067
rect 308 1999 366 2033
rect 308 1965 320 1999
rect 354 1965 366 1999
rect 308 1931 366 1965
rect 308 1897 320 1931
rect 354 1897 366 1931
rect 308 1863 366 1897
rect 308 1829 320 1863
rect 354 1829 366 1863
rect 308 1795 366 1829
rect 308 1761 320 1795
rect 354 1761 366 1795
rect 308 1727 366 1761
rect 308 1693 320 1727
rect 354 1693 366 1727
rect 308 1659 366 1693
rect 308 1625 320 1659
rect 354 1625 366 1659
rect 308 1591 366 1625
rect 308 1557 320 1591
rect 354 1557 366 1591
rect 308 1523 366 1557
rect 308 1489 320 1523
rect 354 1489 366 1523
rect 308 1455 366 1489
rect 308 1421 320 1455
rect 354 1421 366 1455
rect 308 1387 366 1421
rect 308 1353 320 1387
rect 354 1353 366 1387
rect 308 1319 366 1353
rect 308 1285 320 1319
rect 354 1285 366 1319
rect 308 1251 366 1285
rect 308 1217 320 1251
rect 354 1217 366 1251
rect 308 1183 366 1217
rect 308 1149 320 1183
rect 354 1149 366 1183
rect 308 1115 366 1149
rect 308 1081 320 1115
rect 354 1081 366 1115
rect 308 1047 366 1081
rect 308 1013 320 1047
rect 354 1013 366 1047
rect 308 979 366 1013
rect 308 945 320 979
rect 354 945 366 979
rect 308 906 366 945
<< ndiffc >>
rect -1440 2033 -1406 2067
rect -1440 1965 -1406 1999
rect -1440 1897 -1406 1931
rect -1440 1829 -1406 1863
rect -1440 1761 -1406 1795
rect -1440 1693 -1406 1727
rect -1440 1625 -1406 1659
rect -1440 1557 -1406 1591
rect -1440 1489 -1406 1523
rect -1440 1421 -1406 1455
rect -1440 1353 -1406 1387
rect -1440 1285 -1406 1319
rect -1440 1217 -1406 1251
rect -1440 1149 -1406 1183
rect -1440 1081 -1406 1115
rect -1440 1013 -1406 1047
rect -1440 945 -1406 979
rect -1352 2033 -1318 2067
rect -1352 1965 -1318 1999
rect -1352 1897 -1318 1931
rect -1352 1829 -1318 1863
rect -1352 1761 -1318 1795
rect -1352 1693 -1318 1727
rect -1352 1625 -1318 1659
rect -1352 1557 -1318 1591
rect -1352 1489 -1318 1523
rect -1352 1421 -1318 1455
rect -1352 1353 -1318 1387
rect -1352 1285 -1318 1319
rect -1352 1217 -1318 1251
rect -1352 1149 -1318 1183
rect -1352 1081 -1318 1115
rect -1352 1013 -1318 1047
rect -1352 945 -1318 979
rect -1264 2033 -1230 2067
rect -1264 1965 -1230 1999
rect -1264 1897 -1230 1931
rect -1264 1829 -1230 1863
rect -1264 1761 -1230 1795
rect -1264 1693 -1230 1727
rect -1264 1625 -1230 1659
rect -1264 1557 -1230 1591
rect -1264 1489 -1230 1523
rect -1264 1421 -1230 1455
rect -1264 1353 -1230 1387
rect -1264 1285 -1230 1319
rect -1264 1217 -1230 1251
rect -1264 1149 -1230 1183
rect -1264 1081 -1230 1115
rect -1264 1013 -1230 1047
rect -1264 945 -1230 979
rect -1176 2033 -1142 2067
rect -1176 1965 -1142 1999
rect -1176 1897 -1142 1931
rect -1176 1829 -1142 1863
rect -1176 1761 -1142 1795
rect -1176 1693 -1142 1727
rect -1176 1625 -1142 1659
rect -1176 1557 -1142 1591
rect -1176 1489 -1142 1523
rect -1176 1421 -1142 1455
rect -1176 1353 -1142 1387
rect -1176 1285 -1142 1319
rect -1176 1217 -1142 1251
rect -1176 1149 -1142 1183
rect -1176 1081 -1142 1115
rect -1176 1013 -1142 1047
rect -1176 945 -1142 979
rect -1088 2033 -1054 2067
rect -1088 1965 -1054 1999
rect -1088 1897 -1054 1931
rect -1088 1829 -1054 1863
rect -1088 1761 -1054 1795
rect -1088 1693 -1054 1727
rect -1088 1625 -1054 1659
rect -1088 1557 -1054 1591
rect -1088 1489 -1054 1523
rect -1088 1421 -1054 1455
rect -1088 1353 -1054 1387
rect -1088 1285 -1054 1319
rect -1088 1217 -1054 1251
rect -1088 1149 -1054 1183
rect -1088 1081 -1054 1115
rect -1088 1013 -1054 1047
rect -1088 945 -1054 979
rect -1000 2033 -966 2067
rect -1000 1965 -966 1999
rect -1000 1897 -966 1931
rect -1000 1829 -966 1863
rect -1000 1761 -966 1795
rect -1000 1693 -966 1727
rect -1000 1625 -966 1659
rect -1000 1557 -966 1591
rect -1000 1489 -966 1523
rect -1000 1421 -966 1455
rect -1000 1353 -966 1387
rect -1000 1285 -966 1319
rect -1000 1217 -966 1251
rect -1000 1149 -966 1183
rect -1000 1081 -966 1115
rect -1000 1013 -966 1047
rect -1000 945 -966 979
rect -912 2033 -878 2067
rect -912 1965 -878 1999
rect -912 1897 -878 1931
rect -912 1829 -878 1863
rect -912 1761 -878 1795
rect -912 1693 -878 1727
rect -912 1625 -878 1659
rect -912 1557 -878 1591
rect -912 1489 -878 1523
rect -912 1421 -878 1455
rect -912 1353 -878 1387
rect -912 1285 -878 1319
rect -912 1217 -878 1251
rect -912 1149 -878 1183
rect -912 1081 -878 1115
rect -912 1013 -878 1047
rect -912 945 -878 979
rect -824 2033 -790 2067
rect -824 1965 -790 1999
rect -824 1897 -790 1931
rect -824 1829 -790 1863
rect -824 1761 -790 1795
rect -824 1693 -790 1727
rect -824 1625 -790 1659
rect -824 1557 -790 1591
rect -824 1489 -790 1523
rect -824 1421 -790 1455
rect -824 1353 -790 1387
rect -824 1285 -790 1319
rect -824 1217 -790 1251
rect -824 1149 -790 1183
rect -824 1081 -790 1115
rect -824 1013 -790 1047
rect -824 945 -790 979
rect -736 2033 -702 2067
rect -736 1965 -702 1999
rect -736 1897 -702 1931
rect -736 1829 -702 1863
rect -736 1761 -702 1795
rect -736 1693 -702 1727
rect -736 1625 -702 1659
rect -736 1557 -702 1591
rect -736 1489 -702 1523
rect -736 1421 -702 1455
rect -736 1353 -702 1387
rect -736 1285 -702 1319
rect -736 1217 -702 1251
rect -736 1149 -702 1183
rect -736 1081 -702 1115
rect -736 1013 -702 1047
rect -736 945 -702 979
rect -648 2033 -614 2067
rect -648 1965 -614 1999
rect -648 1897 -614 1931
rect -648 1829 -614 1863
rect -648 1761 -614 1795
rect -648 1693 -614 1727
rect -648 1625 -614 1659
rect -648 1557 -614 1591
rect -648 1489 -614 1523
rect -648 1421 -614 1455
rect -648 1353 -614 1387
rect -648 1285 -614 1319
rect -648 1217 -614 1251
rect -648 1149 -614 1183
rect -648 1081 -614 1115
rect -648 1013 -614 1047
rect -648 945 -614 979
rect -560 2033 -526 2067
rect -560 1965 -526 1999
rect -560 1897 -526 1931
rect -560 1829 -526 1863
rect -560 1761 -526 1795
rect -560 1693 -526 1727
rect -560 1625 -526 1659
rect -560 1557 -526 1591
rect -560 1489 -526 1523
rect -560 1421 -526 1455
rect -560 1353 -526 1387
rect -560 1285 -526 1319
rect -560 1217 -526 1251
rect -560 1149 -526 1183
rect -560 1081 -526 1115
rect -560 1013 -526 1047
rect -560 945 -526 979
rect -472 2033 -438 2067
rect -472 1965 -438 1999
rect -472 1897 -438 1931
rect -472 1829 -438 1863
rect -472 1761 -438 1795
rect -472 1693 -438 1727
rect -472 1625 -438 1659
rect -472 1557 -438 1591
rect -472 1489 -438 1523
rect -472 1421 -438 1455
rect -472 1353 -438 1387
rect -472 1285 -438 1319
rect -472 1217 -438 1251
rect -472 1149 -438 1183
rect -472 1081 -438 1115
rect -472 1013 -438 1047
rect -472 945 -438 979
rect -384 2033 -350 2067
rect -384 1965 -350 1999
rect -384 1897 -350 1931
rect -384 1829 -350 1863
rect -384 1761 -350 1795
rect -384 1693 -350 1727
rect -384 1625 -350 1659
rect -384 1557 -350 1591
rect -384 1489 -350 1523
rect -384 1421 -350 1455
rect -384 1353 -350 1387
rect -384 1285 -350 1319
rect -384 1217 -350 1251
rect -384 1149 -350 1183
rect -384 1081 -350 1115
rect -384 1013 -350 1047
rect -384 945 -350 979
rect -296 2033 -262 2067
rect -296 1965 -262 1999
rect -296 1897 -262 1931
rect -296 1829 -262 1863
rect -296 1761 -262 1795
rect -296 1693 -262 1727
rect -296 1625 -262 1659
rect -296 1557 -262 1591
rect -296 1489 -262 1523
rect -296 1421 -262 1455
rect -296 1353 -262 1387
rect -296 1285 -262 1319
rect -296 1217 -262 1251
rect -296 1149 -262 1183
rect -296 1081 -262 1115
rect -296 1013 -262 1047
rect -296 945 -262 979
rect -208 2033 -174 2067
rect -208 1965 -174 1999
rect -208 1897 -174 1931
rect -208 1829 -174 1863
rect -208 1761 -174 1795
rect -208 1693 -174 1727
rect -208 1625 -174 1659
rect -208 1557 -174 1591
rect -208 1489 -174 1523
rect -208 1421 -174 1455
rect -208 1353 -174 1387
rect -208 1285 -174 1319
rect -208 1217 -174 1251
rect -208 1149 -174 1183
rect -208 1081 -174 1115
rect -208 1013 -174 1047
rect -208 945 -174 979
rect -120 2033 -86 2067
rect -120 1965 -86 1999
rect -120 1897 -86 1931
rect -120 1829 -86 1863
rect -120 1761 -86 1795
rect -120 1693 -86 1727
rect -120 1625 -86 1659
rect -120 1557 -86 1591
rect -120 1489 -86 1523
rect -120 1421 -86 1455
rect -120 1353 -86 1387
rect -120 1285 -86 1319
rect -120 1217 -86 1251
rect -120 1149 -86 1183
rect -120 1081 -86 1115
rect -120 1013 -86 1047
rect -120 945 -86 979
rect -32 2033 2 2067
rect -32 1965 2 1999
rect -32 1897 2 1931
rect -32 1829 2 1863
rect -32 1761 2 1795
rect -32 1693 2 1727
rect -32 1625 2 1659
rect -32 1557 2 1591
rect -32 1489 2 1523
rect -32 1421 2 1455
rect -32 1353 2 1387
rect -32 1285 2 1319
rect -32 1217 2 1251
rect -32 1149 2 1183
rect -32 1081 2 1115
rect -32 1013 2 1047
rect -32 945 2 979
rect 56 2033 90 2067
rect 56 1965 90 1999
rect 56 1897 90 1931
rect 56 1829 90 1863
rect 56 1761 90 1795
rect 56 1693 90 1727
rect 56 1625 90 1659
rect 56 1557 90 1591
rect 56 1489 90 1523
rect 56 1421 90 1455
rect 56 1353 90 1387
rect 56 1285 90 1319
rect 56 1217 90 1251
rect 56 1149 90 1183
rect 56 1081 90 1115
rect 56 1013 90 1047
rect 56 945 90 979
rect 144 2033 178 2067
rect 144 1965 178 1999
rect 144 1897 178 1931
rect 144 1829 178 1863
rect 144 1761 178 1795
rect 144 1693 178 1727
rect 144 1625 178 1659
rect 144 1557 178 1591
rect 144 1489 178 1523
rect 144 1421 178 1455
rect 144 1353 178 1387
rect 144 1285 178 1319
rect 144 1217 178 1251
rect 144 1149 178 1183
rect 144 1081 178 1115
rect 144 1013 178 1047
rect 144 945 178 979
rect 232 2033 266 2067
rect 232 1965 266 1999
rect 232 1897 266 1931
rect 232 1829 266 1863
rect 232 1761 266 1795
rect 232 1693 266 1727
rect 232 1625 266 1659
rect 232 1557 266 1591
rect 232 1489 266 1523
rect 232 1421 266 1455
rect 232 1353 266 1387
rect 232 1285 266 1319
rect 232 1217 266 1251
rect 232 1149 266 1183
rect 232 1081 266 1115
rect 232 1013 266 1047
rect 232 945 266 979
rect 320 2033 354 2067
rect 320 1965 354 1999
rect 320 1897 354 1931
rect 320 1829 354 1863
rect 320 1761 354 1795
rect 320 1693 354 1727
rect 320 1625 354 1659
rect 320 1557 354 1591
rect 320 1489 354 1523
rect 320 1421 354 1455
rect 320 1353 354 1387
rect 320 1285 354 1319
rect 320 1217 354 1251
rect 320 1149 354 1183
rect 320 1081 354 1115
rect 320 1013 354 1047
rect 320 945 354 979
<< psubdiff >>
rect 2715 2562 2788 2563
rect -1685 2560 2788 2562
rect -1685 2458 -1420 2560
rect 2490 2458 2788 2560
rect -1685 2457 2788 2458
rect -5926 2222 -5819 2256
rect -5785 2222 -5751 2256
rect -5717 2222 -5683 2256
rect -5649 2222 -5615 2256
rect -5581 2222 -5547 2256
rect -5513 2222 -5479 2256
rect -5445 2222 -5411 2256
rect -5377 2222 -5343 2256
rect -5309 2222 -5275 2256
rect -5241 2222 -5207 2256
rect -5173 2222 -5139 2256
rect -5105 2222 -5071 2256
rect -5037 2222 -5003 2256
rect -4969 2222 -4935 2256
rect -4901 2222 -4867 2256
rect -4833 2222 -4799 2256
rect -4765 2222 -4731 2256
rect -4697 2222 -4663 2256
rect -4629 2222 -4595 2256
rect -4561 2222 -4527 2256
rect -4493 2222 -4459 2256
rect -4425 2222 -4391 2256
rect -4357 2222 -4323 2256
rect -4289 2222 -4255 2256
rect -4221 2222 -4187 2256
rect -4153 2222 -4119 2256
rect -4085 2222 -4051 2256
rect -4017 2222 -3983 2256
rect -3949 2222 -3915 2256
rect -3881 2222 -3847 2256
rect -3813 2222 -3779 2256
rect -3745 2222 -3711 2256
rect -3677 2222 -3643 2256
rect -3609 2222 -3575 2256
rect -3541 2222 -3507 2256
rect -3473 2222 -3439 2256
rect -3405 2222 -3371 2256
rect -3337 2222 -3303 2256
rect -3269 2222 -3235 2256
rect -3201 2222 -3167 2256
rect -3133 2222 -3099 2256
rect -3065 2222 -3031 2256
rect -2997 2222 -2963 2256
rect -2929 2222 -2895 2256
rect -2861 2222 -2827 2256
rect -2793 2222 -2759 2256
rect -2725 2222 -2691 2256
rect -2657 2222 -2623 2256
rect -2589 2222 -2555 2256
rect -2521 2222 -2487 2256
rect -2453 2222 -2419 2256
rect -2385 2222 -2351 2256
rect -2317 2222 -2283 2256
rect -2249 2222 -2215 2256
rect -2181 2222 -2147 2256
rect -2113 2222 -2079 2256
rect -2045 2222 -2011 2256
rect -1977 2222 -1943 2256
rect -1909 2222 -1802 2256
rect -5926 2142 -5892 2222
rect -1836 2142 -1802 2222
rect -5926 2074 -5892 2108
rect -1836 2074 -1802 2108
rect -5926 1960 -5892 2040
rect -1836 1960 -1802 2040
rect -5926 1926 -5819 1960
rect -5785 1926 -5751 1960
rect -5717 1926 -5683 1960
rect -5649 1926 -5615 1960
rect -5581 1926 -5547 1960
rect -5513 1926 -5479 1960
rect -5445 1926 -5411 1960
rect -5377 1926 -5343 1960
rect -5309 1926 -5275 1960
rect -5241 1926 -5207 1960
rect -5173 1926 -5139 1960
rect -5105 1926 -5071 1960
rect -5037 1926 -5003 1960
rect -4969 1926 -4935 1960
rect -4901 1926 -4867 1960
rect -4833 1926 -4799 1960
rect -4765 1926 -4731 1960
rect -4697 1926 -4663 1960
rect -4629 1926 -4595 1960
rect -4561 1926 -4527 1960
rect -4493 1926 -4459 1960
rect -4425 1926 -4391 1960
rect -4357 1926 -4323 1960
rect -4289 1926 -4255 1960
rect -4221 1926 -4187 1960
rect -4153 1926 -4119 1960
rect -4085 1926 -4051 1960
rect -4017 1926 -3983 1960
rect -3949 1926 -3915 1960
rect -3881 1926 -3847 1960
rect -3813 1926 -3779 1960
rect -3745 1926 -3711 1960
rect -3677 1926 -3643 1960
rect -3609 1926 -3575 1960
rect -3541 1926 -3507 1960
rect -3473 1926 -3439 1960
rect -3405 1926 -3371 1960
rect -3337 1926 -3303 1960
rect -3269 1926 -3235 1960
rect -3201 1926 -3167 1960
rect -3133 1926 -3099 1960
rect -3065 1926 -3031 1960
rect -2997 1926 -2963 1960
rect -2929 1926 -2895 1960
rect -2861 1926 -2827 1960
rect -2793 1926 -2759 1960
rect -2725 1926 -2691 1960
rect -2657 1926 -2623 1960
rect -2589 1926 -2555 1960
rect -2521 1926 -2487 1960
rect -2453 1926 -2419 1960
rect -2385 1926 -2351 1960
rect -2317 1926 -2283 1960
rect -2249 1926 -2215 1960
rect -2181 1926 -2147 1960
rect -2113 1926 -2079 1960
rect -2045 1926 -2011 1960
rect -1977 1926 -1943 1960
rect -1909 1926 -1802 1960
rect -1685 2118 -1612 2457
rect -1685 2084 -1666 2118
rect -1632 2084 -1612 2118
rect -1685 2050 -1612 2084
rect -1685 2016 -1666 2050
rect -1632 2016 -1612 2050
rect -1685 1982 -1612 2016
rect -1685 1948 -1666 1982
rect -1632 1948 -1612 1982
rect -1685 1914 -1612 1948
rect -1685 1880 -1666 1914
rect -1632 1880 -1612 1914
rect -1685 1846 -1612 1880
rect -1685 1812 -1666 1846
rect -1632 1812 -1612 1846
rect -1685 1778 -1612 1812
rect -5931 1713 -5824 1747
rect -5790 1713 -5756 1747
rect -5722 1713 -5688 1747
rect -5654 1713 -5620 1747
rect -5586 1713 -5552 1747
rect -5518 1713 -5484 1747
rect -5450 1713 -5416 1747
rect -5382 1713 -5348 1747
rect -5314 1713 -5280 1747
rect -5246 1713 -5212 1747
rect -5178 1713 -5144 1747
rect -5110 1713 -5076 1747
rect -5042 1713 -5008 1747
rect -4974 1713 -4940 1747
rect -4906 1713 -4872 1747
rect -4838 1713 -4804 1747
rect -4770 1713 -4736 1747
rect -4702 1713 -4668 1747
rect -4634 1713 -4600 1747
rect -4566 1713 -4532 1747
rect -4498 1713 -4464 1747
rect -4430 1713 -4396 1747
rect -4362 1713 -4328 1747
rect -4294 1713 -4260 1747
rect -4226 1713 -4192 1747
rect -4158 1713 -4124 1747
rect -4090 1713 -4056 1747
rect -4022 1713 -3988 1747
rect -3954 1713 -3920 1747
rect -3886 1713 -3852 1747
rect -3818 1713 -3784 1747
rect -3750 1713 -3716 1747
rect -3682 1713 -3648 1747
rect -3614 1713 -3580 1747
rect -3546 1713 -3512 1747
rect -3478 1713 -3444 1747
rect -3410 1713 -3376 1747
rect -3342 1713 -3308 1747
rect -3274 1713 -3240 1747
rect -3206 1713 -3172 1747
rect -3138 1713 -3104 1747
rect -3070 1713 -3036 1747
rect -3002 1713 -2968 1747
rect -2934 1713 -2900 1747
rect -2866 1713 -2832 1747
rect -2798 1713 -2764 1747
rect -2730 1713 -2696 1747
rect -2662 1713 -2628 1747
rect -2594 1713 -2560 1747
rect -2526 1713 -2492 1747
rect -2458 1713 -2424 1747
rect -2390 1713 -2356 1747
rect -2322 1713 -2288 1747
rect -2254 1713 -2220 1747
rect -2186 1713 -2152 1747
rect -2118 1713 -2084 1747
rect -2050 1713 -2016 1747
rect -1982 1713 -1948 1747
rect -1914 1713 -1807 1747
rect -5931 1633 -5897 1713
rect -1841 1633 -1807 1713
rect -5931 1565 -5897 1599
rect -1841 1565 -1807 1599
rect -5931 1451 -5897 1531
rect -1841 1451 -1807 1531
rect -5931 1417 -5824 1451
rect -5790 1417 -5756 1451
rect -5722 1417 -5688 1451
rect -5654 1417 -5620 1451
rect -5586 1417 -5552 1451
rect -5518 1417 -5484 1451
rect -5450 1417 -5416 1451
rect -5382 1417 -5348 1451
rect -5314 1417 -5280 1451
rect -5246 1417 -5212 1451
rect -5178 1417 -5144 1451
rect -5110 1417 -5076 1451
rect -5042 1417 -5008 1451
rect -4974 1417 -4940 1451
rect -4906 1417 -4872 1451
rect -4838 1417 -4804 1451
rect -4770 1417 -4736 1451
rect -4702 1417 -4668 1451
rect -4634 1417 -4600 1451
rect -4566 1417 -4532 1451
rect -4498 1417 -4464 1451
rect -4430 1417 -4396 1451
rect -4362 1417 -4328 1451
rect -4294 1417 -4260 1451
rect -4226 1417 -4192 1451
rect -4158 1417 -4124 1451
rect -4090 1417 -4056 1451
rect -4022 1417 -3988 1451
rect -3954 1417 -3920 1451
rect -3886 1417 -3852 1451
rect -3818 1417 -3784 1451
rect -3750 1417 -3716 1451
rect -3682 1417 -3648 1451
rect -3614 1417 -3580 1451
rect -3546 1417 -3512 1451
rect -3478 1417 -3444 1451
rect -3410 1417 -3376 1451
rect -3342 1417 -3308 1451
rect -3274 1417 -3240 1451
rect -3206 1417 -3172 1451
rect -3138 1417 -3104 1451
rect -3070 1417 -3036 1451
rect -3002 1417 -2968 1451
rect -2934 1417 -2900 1451
rect -2866 1417 -2832 1451
rect -2798 1417 -2764 1451
rect -2730 1417 -2696 1451
rect -2662 1417 -2628 1451
rect -2594 1417 -2560 1451
rect -2526 1417 -2492 1451
rect -2458 1417 -2424 1451
rect -2390 1417 -2356 1451
rect -2322 1417 -2288 1451
rect -2254 1417 -2220 1451
rect -2186 1417 -2152 1451
rect -2118 1417 -2084 1451
rect -2050 1417 -2016 1451
rect -1982 1417 -1948 1451
rect -1914 1417 -1807 1451
rect -1685 1744 -1666 1778
rect -1632 1744 -1612 1778
rect -1685 1710 -1612 1744
rect -1685 1676 -1666 1710
rect -1632 1676 -1612 1710
rect -1685 1642 -1612 1676
rect -1685 1608 -1666 1642
rect -1632 1608 -1612 1642
rect -1685 1574 -1612 1608
rect -1685 1540 -1666 1574
rect -1632 1540 -1612 1574
rect -1685 1506 -1612 1540
rect -1685 1472 -1666 1506
rect -1632 1472 -1612 1506
rect -1685 1438 -1612 1472
rect -1685 1404 -1666 1438
rect -1632 1404 -1612 1438
rect -1685 1370 -1612 1404
rect -1685 1336 -1666 1370
rect -1632 1336 -1612 1370
rect -1685 1302 -1612 1336
rect -1685 1268 -1666 1302
rect -1632 1268 -1612 1302
rect -1685 1234 -1612 1268
rect -5970 1174 -5863 1208
rect -5829 1174 -5795 1208
rect -5761 1174 -5727 1208
rect -5693 1174 -5659 1208
rect -5625 1174 -5591 1208
rect -5557 1174 -5523 1208
rect -5489 1174 -5455 1208
rect -5421 1174 -5387 1208
rect -5353 1174 -5319 1208
rect -5285 1174 -5251 1208
rect -5217 1174 -5183 1208
rect -5149 1174 -5115 1208
rect -5081 1174 -5047 1208
rect -5013 1174 -4979 1208
rect -4945 1174 -4911 1208
rect -4877 1174 -4843 1208
rect -4809 1174 -4775 1208
rect -4741 1174 -4707 1208
rect -4673 1174 -4639 1208
rect -4605 1174 -4571 1208
rect -4537 1174 -4503 1208
rect -4469 1174 -4435 1208
rect -4401 1174 -4367 1208
rect -4333 1174 -4299 1208
rect -4265 1174 -4231 1208
rect -4197 1174 -4163 1208
rect -4129 1174 -4095 1208
rect -4061 1174 -4027 1208
rect -3993 1174 -3959 1208
rect -3925 1174 -3891 1208
rect -3857 1174 -3823 1208
rect -3789 1174 -3755 1208
rect -3721 1174 -3687 1208
rect -3653 1174 -3619 1208
rect -3585 1174 -3551 1208
rect -3517 1174 -3483 1208
rect -3449 1174 -3415 1208
rect -3381 1174 -3347 1208
rect -3313 1174 -3279 1208
rect -3245 1174 -3211 1208
rect -3177 1174 -3143 1208
rect -3109 1174 -3075 1208
rect -3041 1174 -3007 1208
rect -2973 1174 -2939 1208
rect -2905 1174 -2871 1208
rect -2837 1174 -2803 1208
rect -2769 1174 -2735 1208
rect -2701 1174 -2667 1208
rect -2633 1174 -2599 1208
rect -2565 1174 -2531 1208
rect -2497 1174 -2463 1208
rect -2429 1174 -2395 1208
rect -2361 1174 -2327 1208
rect -2293 1174 -2259 1208
rect -2225 1174 -2191 1208
rect -2157 1174 -2123 1208
rect -2089 1174 -2055 1208
rect -2021 1174 -1987 1208
rect -1953 1174 -1846 1208
rect -5970 1094 -5936 1174
rect -1880 1094 -1846 1174
rect -5970 1026 -5936 1060
rect -1880 1026 -1846 1060
rect -5970 912 -5936 992
rect -1880 912 -1846 992
rect -5970 878 -5863 912
rect -5829 878 -5795 912
rect -5761 878 -5727 912
rect -5693 878 -5659 912
rect -5625 878 -5591 912
rect -5557 878 -5523 912
rect -5489 878 -5455 912
rect -5421 878 -5387 912
rect -5353 878 -5319 912
rect -5285 878 -5251 912
rect -5217 878 -5183 912
rect -5149 878 -5115 912
rect -5081 878 -5047 912
rect -5013 878 -4979 912
rect -4945 878 -4911 912
rect -4877 878 -4843 912
rect -4809 878 -4775 912
rect -4741 878 -4707 912
rect -4673 878 -4639 912
rect -4605 878 -4571 912
rect -4537 878 -4503 912
rect -4469 878 -4435 912
rect -4401 878 -4367 912
rect -4333 878 -4299 912
rect -4265 878 -4231 912
rect -4197 878 -4163 912
rect -4129 878 -4095 912
rect -4061 878 -4027 912
rect -3993 878 -3959 912
rect -3925 878 -3891 912
rect -3857 878 -3823 912
rect -3789 878 -3755 912
rect -3721 878 -3687 912
rect -3653 878 -3619 912
rect -3585 878 -3551 912
rect -3517 878 -3483 912
rect -3449 878 -3415 912
rect -3381 878 -3347 912
rect -3313 878 -3279 912
rect -3245 878 -3211 912
rect -3177 878 -3143 912
rect -3109 878 -3075 912
rect -3041 878 -3007 912
rect -2973 878 -2939 912
rect -2905 878 -2871 912
rect -2837 878 -2803 912
rect -2769 878 -2735 912
rect -2701 878 -2667 912
rect -2633 878 -2599 912
rect -2565 878 -2531 912
rect -2497 878 -2463 912
rect -2429 878 -2395 912
rect -2361 878 -2327 912
rect -2293 878 -2259 912
rect -2225 878 -2191 912
rect -2157 878 -2123 912
rect -2089 878 -2055 912
rect -2021 878 -1987 912
rect -1953 878 -1846 912
rect -1685 1200 -1666 1234
rect -1632 1200 -1612 1234
rect -1685 1166 -1612 1200
rect -1685 1132 -1666 1166
rect -1632 1132 -1612 1166
rect -1685 1098 -1612 1132
rect -1685 1064 -1666 1098
rect -1632 1064 -1612 1098
rect -1685 1030 -1612 1064
rect -1685 996 -1666 1030
rect -1632 996 -1612 1030
rect -1685 962 -1612 996
rect -1685 928 -1666 962
rect -1632 928 -1612 962
rect -1685 437 -1612 928
rect 2715 1973 2788 2457
rect 2715 1939 2734 1973
rect 2768 1939 2788 1973
rect 2715 1905 2788 1939
rect 2715 1871 2734 1905
rect 2768 1871 2788 1905
rect 2715 1837 2788 1871
rect 2715 1803 2734 1837
rect 2768 1803 2788 1837
rect 2715 1769 2788 1803
rect 2715 1735 2734 1769
rect 2768 1735 2788 1769
rect 2715 1701 2788 1735
rect 2715 1667 2734 1701
rect 2768 1667 2788 1701
rect 2715 1633 2788 1667
rect 2715 1599 2734 1633
rect 2768 1599 2788 1633
rect 2715 1565 2788 1599
rect 2715 1531 2734 1565
rect 2768 1531 2788 1565
rect 2715 1497 2788 1531
rect 2715 1463 2734 1497
rect 2768 1463 2788 1497
rect 2715 1429 2788 1463
rect 2715 1395 2734 1429
rect 2768 1395 2788 1429
rect 2715 1361 2788 1395
rect 2715 1327 2734 1361
rect 2768 1327 2788 1361
rect 2715 1293 2788 1327
rect 2715 1259 2734 1293
rect 2768 1259 2788 1293
rect 2715 1225 2788 1259
rect 2715 1191 2734 1225
rect 2768 1191 2788 1225
rect 2715 1157 2788 1191
rect 2715 1123 2734 1157
rect 2768 1123 2788 1157
rect 2715 1089 2788 1123
rect 2715 1055 2734 1089
rect 2768 1055 2788 1089
rect 2715 1021 2788 1055
rect 2715 987 2734 1021
rect 2768 987 2788 1021
rect 2715 953 2788 987
rect 2715 919 2734 953
rect 2768 919 2788 953
rect 2715 885 2788 919
rect 2715 851 2734 885
rect 2768 851 2788 885
rect 2715 817 2788 851
rect 2715 783 2734 817
rect 2768 783 2788 817
rect 2715 437 2788 783
rect -1685 435 2788 437
rect -1685 333 -1454 435
rect 2524 333 2788 435
rect -1685 332 2788 333
<< psubdiffcont >>
rect -1420 2458 2490 2560
rect -5819 2222 -5785 2256
rect -5751 2222 -5717 2256
rect -5683 2222 -5649 2256
rect -5615 2222 -5581 2256
rect -5547 2222 -5513 2256
rect -5479 2222 -5445 2256
rect -5411 2222 -5377 2256
rect -5343 2222 -5309 2256
rect -5275 2222 -5241 2256
rect -5207 2222 -5173 2256
rect -5139 2222 -5105 2256
rect -5071 2222 -5037 2256
rect -5003 2222 -4969 2256
rect -4935 2222 -4901 2256
rect -4867 2222 -4833 2256
rect -4799 2222 -4765 2256
rect -4731 2222 -4697 2256
rect -4663 2222 -4629 2256
rect -4595 2222 -4561 2256
rect -4527 2222 -4493 2256
rect -4459 2222 -4425 2256
rect -4391 2222 -4357 2256
rect -4323 2222 -4289 2256
rect -4255 2222 -4221 2256
rect -4187 2222 -4153 2256
rect -4119 2222 -4085 2256
rect -4051 2222 -4017 2256
rect -3983 2222 -3949 2256
rect -3915 2222 -3881 2256
rect -3847 2222 -3813 2256
rect -3779 2222 -3745 2256
rect -3711 2222 -3677 2256
rect -3643 2222 -3609 2256
rect -3575 2222 -3541 2256
rect -3507 2222 -3473 2256
rect -3439 2222 -3405 2256
rect -3371 2222 -3337 2256
rect -3303 2222 -3269 2256
rect -3235 2222 -3201 2256
rect -3167 2222 -3133 2256
rect -3099 2222 -3065 2256
rect -3031 2222 -2997 2256
rect -2963 2222 -2929 2256
rect -2895 2222 -2861 2256
rect -2827 2222 -2793 2256
rect -2759 2222 -2725 2256
rect -2691 2222 -2657 2256
rect -2623 2222 -2589 2256
rect -2555 2222 -2521 2256
rect -2487 2222 -2453 2256
rect -2419 2222 -2385 2256
rect -2351 2222 -2317 2256
rect -2283 2222 -2249 2256
rect -2215 2222 -2181 2256
rect -2147 2222 -2113 2256
rect -2079 2222 -2045 2256
rect -2011 2222 -1977 2256
rect -1943 2222 -1909 2256
rect -5926 2108 -5892 2142
rect -5926 2040 -5892 2074
rect -1836 2108 -1802 2142
rect -1836 2040 -1802 2074
rect -5819 1926 -5785 1960
rect -5751 1926 -5717 1960
rect -5683 1926 -5649 1960
rect -5615 1926 -5581 1960
rect -5547 1926 -5513 1960
rect -5479 1926 -5445 1960
rect -5411 1926 -5377 1960
rect -5343 1926 -5309 1960
rect -5275 1926 -5241 1960
rect -5207 1926 -5173 1960
rect -5139 1926 -5105 1960
rect -5071 1926 -5037 1960
rect -5003 1926 -4969 1960
rect -4935 1926 -4901 1960
rect -4867 1926 -4833 1960
rect -4799 1926 -4765 1960
rect -4731 1926 -4697 1960
rect -4663 1926 -4629 1960
rect -4595 1926 -4561 1960
rect -4527 1926 -4493 1960
rect -4459 1926 -4425 1960
rect -4391 1926 -4357 1960
rect -4323 1926 -4289 1960
rect -4255 1926 -4221 1960
rect -4187 1926 -4153 1960
rect -4119 1926 -4085 1960
rect -4051 1926 -4017 1960
rect -3983 1926 -3949 1960
rect -3915 1926 -3881 1960
rect -3847 1926 -3813 1960
rect -3779 1926 -3745 1960
rect -3711 1926 -3677 1960
rect -3643 1926 -3609 1960
rect -3575 1926 -3541 1960
rect -3507 1926 -3473 1960
rect -3439 1926 -3405 1960
rect -3371 1926 -3337 1960
rect -3303 1926 -3269 1960
rect -3235 1926 -3201 1960
rect -3167 1926 -3133 1960
rect -3099 1926 -3065 1960
rect -3031 1926 -2997 1960
rect -2963 1926 -2929 1960
rect -2895 1926 -2861 1960
rect -2827 1926 -2793 1960
rect -2759 1926 -2725 1960
rect -2691 1926 -2657 1960
rect -2623 1926 -2589 1960
rect -2555 1926 -2521 1960
rect -2487 1926 -2453 1960
rect -2419 1926 -2385 1960
rect -2351 1926 -2317 1960
rect -2283 1926 -2249 1960
rect -2215 1926 -2181 1960
rect -2147 1926 -2113 1960
rect -2079 1926 -2045 1960
rect -2011 1926 -1977 1960
rect -1943 1926 -1909 1960
rect -1666 2084 -1632 2118
rect -1666 2016 -1632 2050
rect -1666 1948 -1632 1982
rect -1666 1880 -1632 1914
rect -1666 1812 -1632 1846
rect -5824 1713 -5790 1747
rect -5756 1713 -5722 1747
rect -5688 1713 -5654 1747
rect -5620 1713 -5586 1747
rect -5552 1713 -5518 1747
rect -5484 1713 -5450 1747
rect -5416 1713 -5382 1747
rect -5348 1713 -5314 1747
rect -5280 1713 -5246 1747
rect -5212 1713 -5178 1747
rect -5144 1713 -5110 1747
rect -5076 1713 -5042 1747
rect -5008 1713 -4974 1747
rect -4940 1713 -4906 1747
rect -4872 1713 -4838 1747
rect -4804 1713 -4770 1747
rect -4736 1713 -4702 1747
rect -4668 1713 -4634 1747
rect -4600 1713 -4566 1747
rect -4532 1713 -4498 1747
rect -4464 1713 -4430 1747
rect -4396 1713 -4362 1747
rect -4328 1713 -4294 1747
rect -4260 1713 -4226 1747
rect -4192 1713 -4158 1747
rect -4124 1713 -4090 1747
rect -4056 1713 -4022 1747
rect -3988 1713 -3954 1747
rect -3920 1713 -3886 1747
rect -3852 1713 -3818 1747
rect -3784 1713 -3750 1747
rect -3716 1713 -3682 1747
rect -3648 1713 -3614 1747
rect -3580 1713 -3546 1747
rect -3512 1713 -3478 1747
rect -3444 1713 -3410 1747
rect -3376 1713 -3342 1747
rect -3308 1713 -3274 1747
rect -3240 1713 -3206 1747
rect -3172 1713 -3138 1747
rect -3104 1713 -3070 1747
rect -3036 1713 -3002 1747
rect -2968 1713 -2934 1747
rect -2900 1713 -2866 1747
rect -2832 1713 -2798 1747
rect -2764 1713 -2730 1747
rect -2696 1713 -2662 1747
rect -2628 1713 -2594 1747
rect -2560 1713 -2526 1747
rect -2492 1713 -2458 1747
rect -2424 1713 -2390 1747
rect -2356 1713 -2322 1747
rect -2288 1713 -2254 1747
rect -2220 1713 -2186 1747
rect -2152 1713 -2118 1747
rect -2084 1713 -2050 1747
rect -2016 1713 -1982 1747
rect -1948 1713 -1914 1747
rect -5931 1599 -5897 1633
rect -5931 1531 -5897 1565
rect -1841 1599 -1807 1633
rect -1841 1531 -1807 1565
rect -5824 1417 -5790 1451
rect -5756 1417 -5722 1451
rect -5688 1417 -5654 1451
rect -5620 1417 -5586 1451
rect -5552 1417 -5518 1451
rect -5484 1417 -5450 1451
rect -5416 1417 -5382 1451
rect -5348 1417 -5314 1451
rect -5280 1417 -5246 1451
rect -5212 1417 -5178 1451
rect -5144 1417 -5110 1451
rect -5076 1417 -5042 1451
rect -5008 1417 -4974 1451
rect -4940 1417 -4906 1451
rect -4872 1417 -4838 1451
rect -4804 1417 -4770 1451
rect -4736 1417 -4702 1451
rect -4668 1417 -4634 1451
rect -4600 1417 -4566 1451
rect -4532 1417 -4498 1451
rect -4464 1417 -4430 1451
rect -4396 1417 -4362 1451
rect -4328 1417 -4294 1451
rect -4260 1417 -4226 1451
rect -4192 1417 -4158 1451
rect -4124 1417 -4090 1451
rect -4056 1417 -4022 1451
rect -3988 1417 -3954 1451
rect -3920 1417 -3886 1451
rect -3852 1417 -3818 1451
rect -3784 1417 -3750 1451
rect -3716 1417 -3682 1451
rect -3648 1417 -3614 1451
rect -3580 1417 -3546 1451
rect -3512 1417 -3478 1451
rect -3444 1417 -3410 1451
rect -3376 1417 -3342 1451
rect -3308 1417 -3274 1451
rect -3240 1417 -3206 1451
rect -3172 1417 -3138 1451
rect -3104 1417 -3070 1451
rect -3036 1417 -3002 1451
rect -2968 1417 -2934 1451
rect -2900 1417 -2866 1451
rect -2832 1417 -2798 1451
rect -2764 1417 -2730 1451
rect -2696 1417 -2662 1451
rect -2628 1417 -2594 1451
rect -2560 1417 -2526 1451
rect -2492 1417 -2458 1451
rect -2424 1417 -2390 1451
rect -2356 1417 -2322 1451
rect -2288 1417 -2254 1451
rect -2220 1417 -2186 1451
rect -2152 1417 -2118 1451
rect -2084 1417 -2050 1451
rect -2016 1417 -1982 1451
rect -1948 1417 -1914 1451
rect -1666 1744 -1632 1778
rect -1666 1676 -1632 1710
rect -1666 1608 -1632 1642
rect -1666 1540 -1632 1574
rect -1666 1472 -1632 1506
rect -1666 1404 -1632 1438
rect -1666 1336 -1632 1370
rect -1666 1268 -1632 1302
rect -5863 1174 -5829 1208
rect -5795 1174 -5761 1208
rect -5727 1174 -5693 1208
rect -5659 1174 -5625 1208
rect -5591 1174 -5557 1208
rect -5523 1174 -5489 1208
rect -5455 1174 -5421 1208
rect -5387 1174 -5353 1208
rect -5319 1174 -5285 1208
rect -5251 1174 -5217 1208
rect -5183 1174 -5149 1208
rect -5115 1174 -5081 1208
rect -5047 1174 -5013 1208
rect -4979 1174 -4945 1208
rect -4911 1174 -4877 1208
rect -4843 1174 -4809 1208
rect -4775 1174 -4741 1208
rect -4707 1174 -4673 1208
rect -4639 1174 -4605 1208
rect -4571 1174 -4537 1208
rect -4503 1174 -4469 1208
rect -4435 1174 -4401 1208
rect -4367 1174 -4333 1208
rect -4299 1174 -4265 1208
rect -4231 1174 -4197 1208
rect -4163 1174 -4129 1208
rect -4095 1174 -4061 1208
rect -4027 1174 -3993 1208
rect -3959 1174 -3925 1208
rect -3891 1174 -3857 1208
rect -3823 1174 -3789 1208
rect -3755 1174 -3721 1208
rect -3687 1174 -3653 1208
rect -3619 1174 -3585 1208
rect -3551 1174 -3517 1208
rect -3483 1174 -3449 1208
rect -3415 1174 -3381 1208
rect -3347 1174 -3313 1208
rect -3279 1174 -3245 1208
rect -3211 1174 -3177 1208
rect -3143 1174 -3109 1208
rect -3075 1174 -3041 1208
rect -3007 1174 -2973 1208
rect -2939 1174 -2905 1208
rect -2871 1174 -2837 1208
rect -2803 1174 -2769 1208
rect -2735 1174 -2701 1208
rect -2667 1174 -2633 1208
rect -2599 1174 -2565 1208
rect -2531 1174 -2497 1208
rect -2463 1174 -2429 1208
rect -2395 1174 -2361 1208
rect -2327 1174 -2293 1208
rect -2259 1174 -2225 1208
rect -2191 1174 -2157 1208
rect -2123 1174 -2089 1208
rect -2055 1174 -2021 1208
rect -1987 1174 -1953 1208
rect -5970 1060 -5936 1094
rect -5970 992 -5936 1026
rect -1880 1060 -1846 1094
rect -1880 992 -1846 1026
rect -5863 878 -5829 912
rect -5795 878 -5761 912
rect -5727 878 -5693 912
rect -5659 878 -5625 912
rect -5591 878 -5557 912
rect -5523 878 -5489 912
rect -5455 878 -5421 912
rect -5387 878 -5353 912
rect -5319 878 -5285 912
rect -5251 878 -5217 912
rect -5183 878 -5149 912
rect -5115 878 -5081 912
rect -5047 878 -5013 912
rect -4979 878 -4945 912
rect -4911 878 -4877 912
rect -4843 878 -4809 912
rect -4775 878 -4741 912
rect -4707 878 -4673 912
rect -4639 878 -4605 912
rect -4571 878 -4537 912
rect -4503 878 -4469 912
rect -4435 878 -4401 912
rect -4367 878 -4333 912
rect -4299 878 -4265 912
rect -4231 878 -4197 912
rect -4163 878 -4129 912
rect -4095 878 -4061 912
rect -4027 878 -3993 912
rect -3959 878 -3925 912
rect -3891 878 -3857 912
rect -3823 878 -3789 912
rect -3755 878 -3721 912
rect -3687 878 -3653 912
rect -3619 878 -3585 912
rect -3551 878 -3517 912
rect -3483 878 -3449 912
rect -3415 878 -3381 912
rect -3347 878 -3313 912
rect -3279 878 -3245 912
rect -3211 878 -3177 912
rect -3143 878 -3109 912
rect -3075 878 -3041 912
rect -3007 878 -2973 912
rect -2939 878 -2905 912
rect -2871 878 -2837 912
rect -2803 878 -2769 912
rect -2735 878 -2701 912
rect -2667 878 -2633 912
rect -2599 878 -2565 912
rect -2531 878 -2497 912
rect -2463 878 -2429 912
rect -2395 878 -2361 912
rect -2327 878 -2293 912
rect -2259 878 -2225 912
rect -2191 878 -2157 912
rect -2123 878 -2089 912
rect -2055 878 -2021 912
rect -1987 878 -1953 912
rect -1666 1200 -1632 1234
rect -1666 1132 -1632 1166
rect -1666 1064 -1632 1098
rect -1666 996 -1632 1030
rect -1666 928 -1632 962
rect 2734 1939 2768 1973
rect 2734 1871 2768 1905
rect 2734 1803 2768 1837
rect 2734 1735 2768 1769
rect 2734 1667 2768 1701
rect 2734 1599 2768 1633
rect 2734 1531 2768 1565
rect 2734 1463 2768 1497
rect 2734 1395 2768 1429
rect 2734 1327 2768 1361
rect 2734 1259 2768 1293
rect 2734 1191 2768 1225
rect 2734 1123 2768 1157
rect 2734 1055 2768 1089
rect 2734 987 2768 1021
rect 2734 919 2768 953
rect 2734 851 2768 885
rect 2734 783 2768 817
rect -1454 333 2524 435
<< poly >>
rect -1394 2242 308 2260
rect -1394 2208 -1342 2242
rect -1308 2208 -1274 2242
rect -1240 2208 -1206 2242
rect -1172 2208 -1138 2242
rect -1104 2208 -1070 2242
rect -1036 2208 -1002 2242
rect -968 2208 -934 2242
rect -900 2208 -866 2242
rect -832 2208 -798 2242
rect -764 2208 -730 2242
rect -696 2208 -662 2242
rect -628 2208 -594 2242
rect -560 2208 -526 2242
rect -492 2208 -458 2242
rect -424 2208 -390 2242
rect -356 2208 -322 2242
rect -288 2208 -254 2242
rect -220 2208 -186 2242
rect -152 2208 -118 2242
rect -84 2208 -50 2242
rect -16 2208 18 2242
rect 52 2208 86 2242
rect 120 2208 154 2242
rect 188 2208 222 2242
rect 256 2208 308 2242
rect -1394 2190 308 2208
rect -1394 2106 -1364 2190
rect -1306 2106 -1276 2132
rect -1218 2106 -1188 2132
rect -1130 2106 -1100 2190
rect -1042 2106 -1012 2190
rect -954 2106 -924 2132
rect -866 2106 -836 2132
rect -778 2106 -748 2190
rect -690 2106 -660 2190
rect -602 2106 -572 2132
rect -514 2106 -484 2132
rect -426 2106 -396 2190
rect -338 2106 -308 2190
rect -250 2106 -220 2132
rect -162 2106 -132 2132
rect -74 2106 -44 2190
rect 14 2106 44 2190
rect 102 2106 132 2132
rect 190 2106 220 2132
rect 278 2106 308 2190
rect 782 2242 2484 2260
rect 782 2208 834 2242
rect 868 2208 902 2242
rect 936 2208 970 2242
rect 1004 2208 1038 2242
rect 1072 2208 1106 2242
rect 1140 2208 1174 2242
rect 1208 2208 1242 2242
rect 1276 2208 1310 2242
rect 1344 2208 1378 2242
rect 1412 2208 1446 2242
rect 1480 2208 1514 2242
rect 1548 2208 1582 2242
rect 1616 2208 1650 2242
rect 1684 2208 1718 2242
rect 1752 2208 1786 2242
rect 1820 2208 1854 2242
rect 1888 2208 1922 2242
rect 1956 2208 1990 2242
rect 2024 2208 2058 2242
rect 2092 2208 2126 2242
rect 2160 2208 2194 2242
rect 2228 2208 2262 2242
rect 2296 2208 2330 2242
rect 2364 2208 2398 2242
rect 2432 2208 2484 2242
rect 782 2190 2484 2208
rect 782 2130 812 2190
rect 1046 2106 1076 2190
rect 1134 2106 1164 2190
rect 1398 2106 1428 2190
rect 1486 2106 1516 2190
rect 1750 2106 1780 2190
rect 1838 2106 1868 2190
rect 2102 2106 2132 2190
rect 2190 2106 2220 2190
rect 2454 2106 2484 2190
rect -1394 880 -1364 906
rect -1306 796 -1276 906
rect -1218 796 -1188 906
rect -1130 880 -1100 906
rect -1042 880 -1012 906
rect -954 796 -924 906
rect -866 796 -836 906
rect -778 880 -748 906
rect -690 880 -660 906
rect -602 796 -572 906
rect -514 796 -484 906
rect -426 880 -396 906
rect -338 880 -308 906
rect -250 796 -220 906
rect -162 796 -132 906
rect -74 880 -44 906
rect 14 880 44 906
rect 102 796 132 906
rect 190 796 220 906
rect 278 880 308 906
rect -1306 778 220 796
rect -1306 744 -1267 778
rect -1233 744 -1199 778
rect -1165 744 -1131 778
rect -1097 744 -1063 778
rect -1029 744 -995 778
rect -961 744 -927 778
rect -893 744 -859 778
rect -825 744 -791 778
rect -757 744 -723 778
rect -689 744 -655 778
rect -621 744 -587 778
rect -553 744 -519 778
rect -485 744 -451 778
rect -417 744 -383 778
rect -349 744 -315 778
rect -281 744 -247 778
rect -213 744 -179 778
rect -145 744 -111 778
rect -77 744 -43 778
rect -9 744 25 778
rect 59 744 93 778
rect 127 744 161 778
rect 195 744 220 778
rect -1306 726 220 744
rect 870 796 900 880
rect 958 796 988 880
rect 1222 796 1252 880
rect 1310 796 1340 880
rect 1574 796 1604 880
rect 1662 796 1692 880
rect 1926 796 1956 880
rect 2014 796 2044 880
rect 2278 796 2308 880
rect 2366 796 2396 906
rect 870 778 2396 796
rect 870 744 895 778
rect 929 744 963 778
rect 997 744 1031 778
rect 1065 744 1099 778
rect 1133 744 1167 778
rect 1201 744 1235 778
rect 1269 744 1303 778
rect 1337 744 1371 778
rect 1405 744 1439 778
rect 1473 744 1507 778
rect 1541 744 1575 778
rect 1609 744 1643 778
rect 1677 744 1711 778
rect 1745 744 1779 778
rect 1813 744 1847 778
rect 1881 744 1915 778
rect 1949 744 1983 778
rect 2017 744 2051 778
rect 2085 744 2119 778
rect 2153 744 2187 778
rect 2221 744 2255 778
rect 2289 744 2323 778
rect 2357 744 2396 778
rect 870 726 2396 744
<< polycont >>
rect -1342 2208 -1308 2242
rect -1274 2208 -1240 2242
rect -1206 2208 -1172 2242
rect -1138 2208 -1104 2242
rect -1070 2208 -1036 2242
rect -1002 2208 -968 2242
rect -934 2208 -900 2242
rect -866 2208 -832 2242
rect -798 2208 -764 2242
rect -730 2208 -696 2242
rect -662 2208 -628 2242
rect -594 2208 -560 2242
rect -526 2208 -492 2242
rect -458 2208 -424 2242
rect -390 2208 -356 2242
rect -322 2208 -288 2242
rect -254 2208 -220 2242
rect -186 2208 -152 2242
rect -118 2208 -84 2242
rect -50 2208 -16 2242
rect 18 2208 52 2242
rect 86 2208 120 2242
rect 154 2208 188 2242
rect 222 2208 256 2242
rect 834 2208 868 2242
rect 902 2208 936 2242
rect 970 2208 1004 2242
rect 1038 2208 1072 2242
rect 1106 2208 1140 2242
rect 1174 2208 1208 2242
rect 1242 2208 1276 2242
rect 1310 2208 1344 2242
rect 1378 2208 1412 2242
rect 1446 2208 1480 2242
rect 1514 2208 1548 2242
rect 1582 2208 1616 2242
rect 1650 2208 1684 2242
rect 1718 2208 1752 2242
rect 1786 2208 1820 2242
rect 1854 2208 1888 2242
rect 1922 2208 1956 2242
rect 1990 2208 2024 2242
rect 2058 2208 2092 2242
rect 2126 2208 2160 2242
rect 2194 2208 2228 2242
rect 2262 2208 2296 2242
rect 2330 2208 2364 2242
rect 2398 2208 2432 2242
rect -1267 744 -1233 778
rect -1199 744 -1165 778
rect -1131 744 -1097 778
rect -1063 744 -1029 778
rect -995 744 -961 778
rect -927 744 -893 778
rect -859 744 -825 778
rect -791 744 -757 778
rect -723 744 -689 778
rect -655 744 -621 778
rect -587 744 -553 778
rect -519 744 -485 778
rect -451 744 -417 778
rect -383 744 -349 778
rect -315 744 -281 778
rect -247 744 -213 778
rect -179 744 -145 778
rect -111 744 -77 778
rect -43 744 -9 778
rect 25 744 59 778
rect 93 744 127 778
rect 161 744 195 778
rect 895 744 929 778
rect 963 744 997 778
rect 1031 744 1065 778
rect 1099 744 1133 778
rect 1167 744 1201 778
rect 1235 744 1269 778
rect 1303 744 1337 778
rect 1371 744 1405 778
rect 1439 744 1473 778
rect 1507 744 1541 778
rect 1575 744 1609 778
rect 1643 744 1677 778
rect 1711 744 1745 778
rect 1779 744 1813 778
rect 1847 744 1881 778
rect 1915 744 1949 778
rect 1983 744 2017 778
rect 2051 744 2085 778
rect 2119 744 2153 778
rect 2187 744 2221 778
rect 2255 744 2289 778
rect 2323 744 2357 778
<< xpolycontact >>
rect -5796 2056 -5364 2126
rect -2364 2056 -1932 2126
rect -5801 1547 -5369 1617
rect -2369 1547 -1937 1617
rect -5840 1008 -5408 1078
rect -2408 1008 -1976 1078
<< xpolyres >>
rect -5364 2056 -2364 2126
rect -5369 1547 -2369 1617
rect -5408 1008 -2408 1078
<< locali >>
rect -1685 2560 2788 2562
rect -1685 2458 -1420 2560
rect 2490 2458 2788 2560
rect -1685 2457 2788 2458
rect -1685 2305 -1612 2457
rect -1885 2256 -1612 2305
rect 2715 2293 2788 2457
rect -5926 2222 -5819 2256
rect -5785 2222 -5751 2256
rect -5717 2222 -5683 2256
rect -5649 2222 -5615 2256
rect -5581 2222 -5547 2256
rect -5513 2222 -5479 2256
rect -5445 2222 -5411 2256
rect -5377 2222 -5343 2256
rect -5309 2222 -5275 2256
rect -5241 2222 -5207 2256
rect -5173 2222 -5139 2256
rect -5105 2222 -5071 2256
rect -5037 2222 -5003 2256
rect -4969 2222 -4935 2256
rect -4901 2222 -4867 2256
rect -4833 2222 -4799 2256
rect -4765 2222 -4731 2256
rect -4697 2222 -4663 2256
rect -4629 2222 -4595 2256
rect -4561 2222 -4527 2256
rect -4493 2222 -4459 2256
rect -4425 2222 -4391 2256
rect -4357 2222 -4323 2256
rect -4289 2222 -4255 2256
rect -4221 2222 -4187 2256
rect -4153 2222 -4119 2256
rect -4085 2222 -4051 2256
rect -4017 2222 -3983 2256
rect -3949 2222 -3915 2256
rect -3881 2222 -3847 2256
rect -3813 2222 -3779 2256
rect -3745 2222 -3711 2256
rect -3677 2222 -3643 2256
rect -3609 2222 -3575 2256
rect -3541 2222 -3507 2256
rect -3473 2222 -3439 2256
rect -3405 2222 -3371 2256
rect -3337 2222 -3303 2256
rect -3269 2222 -3235 2256
rect -3201 2222 -3167 2256
rect -3133 2222 -3099 2256
rect -3065 2222 -3031 2256
rect -2997 2222 -2963 2256
rect -2929 2222 -2895 2256
rect -2861 2222 -2827 2256
rect -2793 2222 -2759 2256
rect -2725 2222 -2691 2256
rect -2657 2222 -2623 2256
rect -2589 2222 -2555 2256
rect -2521 2222 -2487 2256
rect -2453 2222 -2419 2256
rect -2385 2222 -2351 2256
rect -2317 2222 -2283 2256
rect -2249 2222 -2215 2256
rect -2181 2222 -2147 2256
rect -2113 2222 -2079 2256
rect -2045 2222 -2011 2256
rect -1977 2222 -1943 2256
rect -1909 2222 -1612 2256
rect -5926 2142 -5892 2222
rect -1885 2142 -1612 2222
rect -1394 2242 308 2260
rect -1394 2208 -1352 2242
rect -1308 2208 -1280 2242
rect -1240 2208 -1208 2242
rect -1172 2208 -1138 2242
rect -1102 2208 -1070 2242
rect -1030 2208 -1002 2242
rect -958 2208 -934 2242
rect -886 2208 -866 2242
rect -814 2208 -798 2242
rect -742 2208 -730 2242
rect -670 2208 -662 2242
rect -598 2208 -594 2242
rect -492 2208 -488 2242
rect -424 2208 -416 2242
rect -356 2208 -344 2242
rect -288 2208 -272 2242
rect -220 2208 -200 2242
rect -152 2208 -128 2242
rect -84 2208 -56 2242
rect -16 2208 16 2242
rect 52 2208 86 2242
rect 122 2208 154 2242
rect 194 2208 222 2242
rect 266 2208 308 2242
rect -1394 2190 308 2208
rect 782 2242 2484 2260
rect 782 2208 824 2242
rect 868 2208 896 2242
rect 936 2208 968 2242
rect 1004 2208 1038 2242
rect 1074 2208 1106 2242
rect 1146 2208 1174 2242
rect 1218 2208 1242 2242
rect 1290 2208 1310 2242
rect 1362 2208 1378 2242
rect 1434 2208 1446 2242
rect 1506 2208 1514 2242
rect 1578 2208 1582 2242
rect 1684 2208 1688 2242
rect 1752 2208 1760 2242
rect 1820 2208 1832 2242
rect 1888 2208 1904 2242
rect 1956 2208 1976 2242
rect 2024 2208 2048 2242
rect 2092 2208 2120 2242
rect 2160 2208 2192 2242
rect 2228 2208 2262 2242
rect 2298 2208 2330 2242
rect 2370 2208 2398 2242
rect 2442 2208 2484 2242
rect 782 2190 2484 2208
rect -5926 2074 -5892 2108
rect -1885 2108 -1836 2142
rect -1802 2118 -1612 2142
rect -1802 2108 -1666 2118
rect -1885 2084 -1666 2108
rect -1632 2084 -1612 2118
rect -1885 2074 -1612 2084
rect -5926 1960 -5892 2040
rect -1885 2040 -1836 2074
rect -1802 2050 -1612 2074
rect -1802 2040 -1666 2050
rect -1885 2016 -1666 2040
rect -1632 2016 -1612 2050
rect -1885 1982 -1612 2016
rect -1885 1960 -1666 1982
rect -5926 1926 -5819 1960
rect -5785 1926 -5751 1960
rect -5717 1926 -5683 1960
rect -5649 1926 -5615 1960
rect -5581 1926 -5547 1960
rect -5513 1926 -5479 1960
rect -5445 1926 -5411 1960
rect -5377 1926 -5343 1960
rect -5309 1926 -5275 1960
rect -5241 1926 -5207 1960
rect -5173 1926 -5139 1960
rect -5105 1926 -5071 1960
rect -5037 1926 -5003 1960
rect -4969 1926 -4935 1960
rect -4901 1926 -4867 1960
rect -4833 1926 -4799 1960
rect -4765 1926 -4731 1960
rect -4697 1926 -4663 1960
rect -4629 1926 -4595 1960
rect -4561 1926 -4527 1960
rect -4493 1926 -4459 1960
rect -4425 1926 -4391 1960
rect -4357 1926 -4323 1960
rect -4289 1926 -4255 1960
rect -4221 1926 -4187 1960
rect -4153 1926 -4119 1960
rect -4085 1926 -4051 1960
rect -4017 1926 -3983 1960
rect -3949 1926 -3915 1960
rect -3881 1926 -3847 1960
rect -3813 1926 -3779 1960
rect -3745 1926 -3711 1960
rect -3677 1926 -3643 1960
rect -3609 1926 -3575 1960
rect -3541 1926 -3507 1960
rect -3473 1926 -3439 1960
rect -3405 1926 -3371 1960
rect -3337 1926 -3303 1960
rect -3269 1926 -3235 1960
rect -3201 1926 -3167 1960
rect -3133 1926 -3099 1960
rect -3065 1926 -3031 1960
rect -2997 1926 -2963 1960
rect -2929 1926 -2895 1960
rect -2861 1926 -2827 1960
rect -2793 1926 -2759 1960
rect -2725 1926 -2691 1960
rect -2657 1926 -2623 1960
rect -2589 1926 -2555 1960
rect -2521 1926 -2487 1960
rect -2453 1926 -2419 1960
rect -2385 1926 -2351 1960
rect -2317 1926 -2283 1960
rect -2249 1926 -2215 1960
rect -2181 1926 -2147 1960
rect -2113 1926 -2079 1960
rect -2045 1926 -2011 1960
rect -1977 1926 -1943 1960
rect -1909 1948 -1666 1960
rect -1632 1948 -1612 1982
rect -1909 1926 -1612 1948
rect -4984 1747 -3029 1926
rect -1885 1914 -1612 1926
rect -1885 1880 -1666 1914
rect -1632 1880 -1612 1914
rect -1885 1846 -1612 1880
rect -1885 1812 -1666 1846
rect -1632 1812 -1612 1846
rect -1885 1778 -1612 1812
rect -1885 1747 -1666 1778
rect -5931 1713 -5824 1747
rect -5790 1713 -5756 1747
rect -5722 1713 -5688 1747
rect -5654 1713 -5620 1747
rect -5586 1713 -5552 1747
rect -5518 1713 -5484 1747
rect -5450 1713 -5416 1747
rect -5382 1713 -5348 1747
rect -5314 1713 -5280 1747
rect -5246 1713 -5212 1747
rect -5178 1713 -5144 1747
rect -5110 1713 -5076 1747
rect -5042 1713 -5008 1747
rect -4974 1713 -4940 1747
rect -4906 1713 -4872 1747
rect -4838 1713 -4804 1747
rect -4770 1713 -4736 1747
rect -4702 1713 -4668 1747
rect -4634 1713 -4600 1747
rect -4566 1713 -4532 1747
rect -4498 1713 -4464 1747
rect -4430 1713 -4396 1747
rect -4362 1713 -4328 1747
rect -4294 1713 -4260 1747
rect -4226 1713 -4192 1747
rect -4158 1713 -4124 1747
rect -4090 1713 -4056 1747
rect -4022 1713 -3988 1747
rect -3954 1713 -3920 1747
rect -3886 1713 -3852 1747
rect -3818 1713 -3784 1747
rect -3750 1713 -3716 1747
rect -3682 1713 -3648 1747
rect -3614 1713 -3580 1747
rect -3546 1713 -3512 1747
rect -3478 1713 -3444 1747
rect -3410 1713 -3376 1747
rect -3342 1713 -3308 1747
rect -3274 1713 -3240 1747
rect -3206 1713 -3172 1747
rect -3138 1713 -3104 1747
rect -3070 1713 -3036 1747
rect -3002 1713 -2968 1747
rect -2934 1713 -2900 1747
rect -2866 1713 -2832 1747
rect -2798 1713 -2764 1747
rect -2730 1713 -2696 1747
rect -2662 1713 -2628 1747
rect -2594 1713 -2560 1747
rect -2526 1713 -2492 1747
rect -2458 1713 -2424 1747
rect -2390 1713 -2356 1747
rect -2322 1713 -2288 1747
rect -2254 1713 -2220 1747
rect -2186 1713 -2152 1747
rect -2118 1713 -2084 1747
rect -2050 1713 -2016 1747
rect -1982 1713 -1948 1747
rect -1914 1744 -1666 1747
rect -1632 1744 -1612 1778
rect -1914 1713 -1612 1744
rect -5931 1633 -5897 1713
rect -5931 1565 -5897 1599
rect -5931 1451 -5897 1531
rect -4984 1451 -3029 1713
rect -1885 1710 -1612 1713
rect -1885 1676 -1666 1710
rect -1632 1676 -1612 1710
rect -1885 1642 -1612 1676
rect -1885 1633 -1666 1642
rect -1885 1599 -1841 1633
rect -1807 1608 -1666 1633
rect -1632 1608 -1612 1642
rect -1807 1599 -1612 1608
rect -1885 1574 -1612 1599
rect -1885 1565 -1666 1574
rect -1885 1531 -1841 1565
rect -1807 1540 -1666 1565
rect -1632 1540 -1612 1574
rect -1807 1531 -1612 1540
rect -1885 1506 -1612 1531
rect -1885 1472 -1666 1506
rect -1632 1472 -1612 1506
rect -1885 1451 -1612 1472
rect -5931 1417 -5824 1451
rect -5790 1417 -5756 1451
rect -5722 1417 -5688 1451
rect -5654 1417 -5620 1451
rect -5586 1417 -5552 1451
rect -5518 1417 -5484 1451
rect -5450 1417 -5416 1451
rect -5382 1417 -5348 1451
rect -5314 1417 -5280 1451
rect -5246 1417 -5212 1451
rect -5178 1417 -5144 1451
rect -5110 1417 -5076 1451
rect -5042 1417 -5008 1451
rect -4974 1417 -4940 1451
rect -4906 1417 -4872 1451
rect -4838 1417 -4804 1451
rect -4770 1417 -4736 1451
rect -4702 1417 -4668 1451
rect -4634 1417 -4600 1451
rect -4566 1417 -4532 1451
rect -4498 1417 -4464 1451
rect -4430 1417 -4396 1451
rect -4362 1417 -4328 1451
rect -4294 1417 -4260 1451
rect -4226 1417 -4192 1451
rect -4158 1417 -4124 1451
rect -4090 1417 -4056 1451
rect -4022 1417 -3988 1451
rect -3954 1417 -3920 1451
rect -3886 1417 -3852 1451
rect -3818 1417 -3784 1451
rect -3750 1417 -3716 1451
rect -3682 1417 -3648 1451
rect -3614 1417 -3580 1451
rect -3546 1417 -3512 1451
rect -3478 1417 -3444 1451
rect -3410 1417 -3376 1451
rect -3342 1417 -3308 1451
rect -3274 1417 -3240 1451
rect -3206 1417 -3172 1451
rect -3138 1417 -3104 1451
rect -3070 1417 -3036 1451
rect -3002 1417 -2968 1451
rect -2934 1417 -2900 1451
rect -2866 1417 -2832 1451
rect -2798 1417 -2764 1451
rect -2730 1417 -2696 1451
rect -2662 1417 -2628 1451
rect -2594 1417 -2560 1451
rect -2526 1417 -2492 1451
rect -2458 1417 -2424 1451
rect -2390 1417 -2356 1451
rect -2322 1417 -2288 1451
rect -2254 1417 -2220 1451
rect -2186 1417 -2152 1451
rect -2118 1417 -2084 1451
rect -2050 1417 -2016 1451
rect -1982 1417 -1948 1451
rect -1914 1438 -1612 1451
rect -1914 1417 -1666 1438
rect -4984 1208 -3029 1417
rect -1885 1404 -1666 1417
rect -1632 1404 -1612 1438
rect -1885 1370 -1612 1404
rect -1885 1336 -1666 1370
rect -1632 1336 -1612 1370
rect -1885 1302 -1612 1336
rect -1885 1268 -1666 1302
rect -1632 1268 -1612 1302
rect -1885 1234 -1612 1268
rect -1885 1208 -1666 1234
rect -5970 1174 -5863 1208
rect -5829 1174 -5795 1208
rect -5761 1174 -5727 1208
rect -5693 1174 -5659 1208
rect -5625 1174 -5591 1208
rect -5557 1174 -5523 1208
rect -5489 1174 -5455 1208
rect -5421 1174 -5387 1208
rect -5353 1174 -5319 1208
rect -5285 1174 -5251 1208
rect -5217 1174 -5183 1208
rect -5149 1174 -5115 1208
rect -5081 1174 -5047 1208
rect -5013 1174 -4979 1208
rect -4945 1174 -4911 1208
rect -4877 1174 -4843 1208
rect -4809 1174 -4775 1208
rect -4741 1174 -4707 1208
rect -4673 1174 -4639 1208
rect -4605 1174 -4571 1208
rect -4537 1174 -4503 1208
rect -4469 1174 -4435 1208
rect -4401 1174 -4367 1208
rect -4333 1174 -4299 1208
rect -4265 1174 -4231 1208
rect -4197 1174 -4163 1208
rect -4129 1174 -4095 1208
rect -4061 1174 -4027 1208
rect -3993 1174 -3959 1208
rect -3925 1174 -3891 1208
rect -3857 1174 -3823 1208
rect -3789 1174 -3755 1208
rect -3721 1174 -3687 1208
rect -3653 1174 -3619 1208
rect -3585 1174 -3551 1208
rect -3517 1174 -3483 1208
rect -3449 1174 -3415 1208
rect -3381 1174 -3347 1208
rect -3313 1174 -3279 1208
rect -3245 1174 -3211 1208
rect -3177 1174 -3143 1208
rect -3109 1174 -3075 1208
rect -3041 1174 -3007 1208
rect -2973 1174 -2939 1208
rect -2905 1174 -2871 1208
rect -2837 1174 -2803 1208
rect -2769 1174 -2735 1208
rect -2701 1174 -2667 1208
rect -2633 1174 -2599 1208
rect -2565 1174 -2531 1208
rect -2497 1174 -2463 1208
rect -2429 1174 -2395 1208
rect -2361 1174 -2327 1208
rect -2293 1174 -2259 1208
rect -2225 1174 -2191 1208
rect -2157 1174 -2123 1208
rect -2089 1174 -2055 1208
rect -2021 1174 -1987 1208
rect -1953 1200 -1666 1208
rect -1632 1200 -1612 1234
rect -1953 1174 -1612 1200
rect -5970 1094 -5936 1174
rect -1885 1166 -1612 1174
rect -1885 1132 -1666 1166
rect -1632 1132 -1612 1166
rect -1885 1098 -1612 1132
rect -1885 1094 -1666 1098
rect -5970 1026 -5936 1060
rect -1885 1060 -1880 1094
rect -1846 1064 -1666 1094
rect -1632 1064 -1612 1098
rect -1846 1060 -1612 1064
rect -1885 1030 -1612 1060
rect -1885 1026 -1666 1030
rect -5970 912 -5936 992
rect -1885 992 -1880 1026
rect -1846 996 -1666 1026
rect -1632 996 -1612 1030
rect -1846 992 -1612 996
rect -1885 962 -1612 992
rect -1885 928 -1666 962
rect -1632 928 -1612 962
rect -1885 912 -1612 928
rect -5970 878 -5863 912
rect -5829 878 -5795 912
rect -5761 878 -5727 912
rect -5693 878 -5659 912
rect -5625 878 -5591 912
rect -5557 878 -5523 912
rect -5489 878 -5455 912
rect -5421 878 -5387 912
rect -5353 878 -5319 912
rect -5285 878 -5251 912
rect -5217 878 -5183 912
rect -5149 878 -5115 912
rect -5081 878 -5047 912
rect -5013 878 -4979 912
rect -4945 878 -4911 912
rect -4877 878 -4843 912
rect -4809 878 -4775 912
rect -4741 878 -4707 912
rect -4673 878 -4639 912
rect -4605 878 -4571 912
rect -4537 878 -4503 912
rect -4469 878 -4435 912
rect -4401 878 -4367 912
rect -4333 878 -4299 912
rect -4265 878 -4231 912
rect -4197 878 -4163 912
rect -4129 878 -4095 912
rect -4061 878 -4027 912
rect -3993 878 -3959 912
rect -3925 878 -3891 912
rect -3857 878 -3823 912
rect -3789 878 -3755 912
rect -3721 878 -3687 912
rect -3653 878 -3619 912
rect -3585 878 -3551 912
rect -3517 878 -3483 912
rect -3449 878 -3415 912
rect -3381 878 -3347 912
rect -3313 878 -3279 912
rect -3245 878 -3211 912
rect -3177 878 -3143 912
rect -3109 878 -3075 912
rect -3041 878 -3007 912
rect -2973 878 -2939 912
rect -2905 878 -2871 912
rect -2837 878 -2803 912
rect -2769 878 -2735 912
rect -2701 878 -2667 912
rect -2633 878 -2599 912
rect -2565 878 -2531 912
rect -2497 878 -2463 912
rect -2429 878 -2395 912
rect -2361 878 -2327 912
rect -2293 878 -2259 912
rect -2225 878 -2191 912
rect -2157 878 -2123 912
rect -2089 878 -2055 912
rect -2021 878 -1987 912
rect -1953 878 -1612 912
rect -1440 2067 -1406 2110
rect -1440 1999 -1406 2029
rect -1440 1931 -1406 1957
rect -1440 1863 -1406 1885
rect -1440 1795 -1406 1813
rect -1440 1727 -1406 1741
rect -1440 1659 -1406 1669
rect -1440 1591 -1406 1597
rect -1440 1523 -1406 1525
rect -1440 1487 -1406 1489
rect -1440 1415 -1406 1421
rect -1440 1343 -1406 1353
rect -1440 1271 -1406 1285
rect -1440 1199 -1406 1217
rect -1440 1127 -1406 1149
rect -1440 1055 -1406 1081
rect -1440 983 -1406 1013
rect -1440 902 -1406 945
rect -1352 2067 -1318 2110
rect -1352 1999 -1318 2029
rect -1352 1931 -1318 1957
rect -1352 1863 -1318 1885
rect -1352 1795 -1318 1813
rect -1352 1727 -1318 1741
rect -1352 1659 -1318 1669
rect -1352 1591 -1318 1597
rect -1352 1523 -1318 1525
rect -1352 1487 -1318 1489
rect -1352 1415 -1318 1421
rect -1352 1343 -1318 1353
rect -1352 1271 -1318 1285
rect -1352 1199 -1318 1217
rect -1352 1127 -1318 1149
rect -1352 1055 -1318 1081
rect -1352 983 -1318 1013
rect -1352 902 -1318 945
rect -1264 2067 -1230 2110
rect -1264 1999 -1230 2029
rect -1264 1931 -1230 1957
rect -1264 1863 -1230 1885
rect -1264 1795 -1230 1813
rect -1264 1727 -1230 1741
rect -1264 1659 -1230 1669
rect -1264 1591 -1230 1597
rect -1264 1523 -1230 1525
rect -1264 1487 -1230 1489
rect -1264 1415 -1230 1421
rect -1264 1343 -1230 1353
rect -1264 1271 -1230 1285
rect -1264 1199 -1230 1217
rect -1264 1127 -1230 1149
rect -1264 1055 -1230 1081
rect -1264 983 -1230 1013
rect -1264 902 -1230 945
rect -1176 2067 -1142 2110
rect -1176 1999 -1142 2029
rect -1176 1931 -1142 1957
rect -1176 1863 -1142 1885
rect -1176 1795 -1142 1813
rect -1176 1727 -1142 1741
rect -1176 1659 -1142 1669
rect -1176 1591 -1142 1597
rect -1176 1523 -1142 1525
rect -1176 1487 -1142 1489
rect -1176 1415 -1142 1421
rect -1176 1343 -1142 1353
rect -1176 1271 -1142 1285
rect -1176 1199 -1142 1217
rect -1176 1127 -1142 1149
rect -1176 1055 -1142 1081
rect -1176 983 -1142 1013
rect -1176 902 -1142 945
rect -1088 2067 -1054 2110
rect -1088 1999 -1054 2029
rect -1088 1931 -1054 1957
rect -1088 1863 -1054 1885
rect -1088 1795 -1054 1813
rect -1088 1727 -1054 1741
rect -1088 1659 -1054 1669
rect -1088 1591 -1054 1597
rect -1088 1523 -1054 1525
rect -1088 1487 -1054 1489
rect -1088 1415 -1054 1421
rect -1088 1343 -1054 1353
rect -1088 1271 -1054 1285
rect -1088 1199 -1054 1217
rect -1088 1127 -1054 1149
rect -1088 1055 -1054 1081
rect -1088 983 -1054 1013
rect -1088 902 -1054 945
rect -1000 2067 -966 2110
rect -1000 1999 -966 2029
rect -1000 1931 -966 1957
rect -1000 1863 -966 1885
rect -1000 1795 -966 1813
rect -1000 1727 -966 1741
rect -1000 1659 -966 1669
rect -1000 1591 -966 1597
rect -1000 1523 -966 1525
rect -1000 1487 -966 1489
rect -1000 1415 -966 1421
rect -1000 1343 -966 1353
rect -1000 1271 -966 1285
rect -1000 1199 -966 1217
rect -1000 1127 -966 1149
rect -1000 1055 -966 1081
rect -1000 983 -966 1013
rect -1000 902 -966 945
rect -912 2067 -878 2110
rect -912 1999 -878 2029
rect -912 1931 -878 1957
rect -912 1863 -878 1885
rect -912 1795 -878 1813
rect -912 1727 -878 1741
rect -912 1659 -878 1669
rect -912 1591 -878 1597
rect -912 1523 -878 1525
rect -912 1487 -878 1489
rect -912 1415 -878 1421
rect -912 1343 -878 1353
rect -912 1271 -878 1285
rect -912 1199 -878 1217
rect -912 1127 -878 1149
rect -912 1055 -878 1081
rect -912 983 -878 1013
rect -912 902 -878 945
rect -824 2067 -790 2110
rect -824 1999 -790 2029
rect -824 1931 -790 1957
rect -824 1863 -790 1885
rect -824 1795 -790 1813
rect -824 1727 -790 1741
rect -824 1659 -790 1669
rect -824 1591 -790 1597
rect -824 1523 -790 1525
rect -824 1487 -790 1489
rect -824 1415 -790 1421
rect -824 1343 -790 1353
rect -824 1271 -790 1285
rect -824 1199 -790 1217
rect -824 1127 -790 1149
rect -824 1055 -790 1081
rect -824 983 -790 1013
rect -824 902 -790 945
rect -736 2067 -702 2110
rect -736 1999 -702 2029
rect -736 1931 -702 1957
rect -736 1863 -702 1885
rect -736 1795 -702 1813
rect -736 1727 -702 1741
rect -736 1659 -702 1669
rect -736 1591 -702 1597
rect -736 1523 -702 1525
rect -736 1487 -702 1489
rect -736 1415 -702 1421
rect -736 1343 -702 1353
rect -736 1271 -702 1285
rect -736 1199 -702 1217
rect -736 1127 -702 1149
rect -736 1055 -702 1081
rect -736 983 -702 1013
rect -736 902 -702 945
rect -648 2067 -614 2110
rect -648 1999 -614 2029
rect -648 1931 -614 1957
rect -648 1863 -614 1885
rect -648 1795 -614 1813
rect -648 1727 -614 1741
rect -648 1659 -614 1669
rect -648 1591 -614 1597
rect -648 1523 -614 1525
rect -648 1487 -614 1489
rect -648 1415 -614 1421
rect -648 1343 -614 1353
rect -648 1271 -614 1285
rect -648 1199 -614 1217
rect -648 1127 -614 1149
rect -648 1055 -614 1081
rect -648 983 -614 1013
rect -648 902 -614 945
rect -560 2067 -526 2110
rect -560 1999 -526 2029
rect -560 1931 -526 1957
rect -560 1863 -526 1885
rect -560 1795 -526 1813
rect -560 1727 -526 1741
rect -560 1659 -526 1669
rect -560 1591 -526 1597
rect -560 1523 -526 1525
rect -560 1487 -526 1489
rect -560 1415 -526 1421
rect -560 1343 -526 1353
rect -560 1271 -526 1285
rect -560 1199 -526 1217
rect -560 1127 -526 1149
rect -560 1055 -526 1081
rect -560 983 -526 1013
rect -560 902 -526 945
rect -472 2067 -438 2110
rect -472 1999 -438 2029
rect -472 1931 -438 1957
rect -472 1863 -438 1885
rect -472 1795 -438 1813
rect -472 1727 -438 1741
rect -472 1659 -438 1669
rect -472 1591 -438 1597
rect -472 1523 -438 1525
rect -472 1487 -438 1489
rect -472 1415 -438 1421
rect -472 1343 -438 1353
rect -472 1271 -438 1285
rect -472 1199 -438 1217
rect -472 1127 -438 1149
rect -472 1055 -438 1081
rect -472 983 -438 1013
rect -472 902 -438 945
rect -384 2067 -350 2110
rect -384 1999 -350 2029
rect -384 1931 -350 1957
rect -384 1863 -350 1885
rect -384 1795 -350 1813
rect -384 1727 -350 1741
rect -384 1659 -350 1669
rect -384 1591 -350 1597
rect -384 1523 -350 1525
rect -384 1487 -350 1489
rect -384 1415 -350 1421
rect -384 1343 -350 1353
rect -384 1271 -350 1285
rect -384 1199 -350 1217
rect -384 1127 -350 1149
rect -384 1055 -350 1081
rect -384 983 -350 1013
rect -384 902 -350 945
rect -296 2067 -262 2110
rect -296 1999 -262 2029
rect -296 1931 -262 1957
rect -296 1863 -262 1885
rect -296 1795 -262 1813
rect -296 1727 -262 1741
rect -296 1659 -262 1669
rect -296 1591 -262 1597
rect -296 1523 -262 1525
rect -296 1487 -262 1489
rect -296 1415 -262 1421
rect -296 1343 -262 1353
rect -296 1271 -262 1285
rect -296 1199 -262 1217
rect -296 1127 -262 1149
rect -296 1055 -262 1081
rect -296 983 -262 1013
rect -296 902 -262 945
rect -208 2067 -174 2110
rect -208 1999 -174 2029
rect -208 1931 -174 1957
rect -208 1863 -174 1885
rect -208 1795 -174 1813
rect -208 1727 -174 1741
rect -208 1659 -174 1669
rect -208 1591 -174 1597
rect -208 1523 -174 1525
rect -208 1487 -174 1489
rect -208 1415 -174 1421
rect -208 1343 -174 1353
rect -208 1271 -174 1285
rect -208 1199 -174 1217
rect -208 1127 -174 1149
rect -208 1055 -174 1081
rect -208 983 -174 1013
rect -208 902 -174 945
rect -120 2067 -86 2110
rect -120 1999 -86 2029
rect -120 1931 -86 1957
rect -120 1863 -86 1885
rect -120 1795 -86 1813
rect -120 1727 -86 1741
rect -120 1659 -86 1669
rect -120 1591 -86 1597
rect -120 1523 -86 1525
rect -120 1487 -86 1489
rect -120 1415 -86 1421
rect -120 1343 -86 1353
rect -120 1271 -86 1285
rect -120 1199 -86 1217
rect -120 1127 -86 1149
rect -120 1055 -86 1081
rect -120 983 -86 1013
rect -120 902 -86 945
rect -32 2067 2 2110
rect -32 1999 2 2029
rect -32 1931 2 1957
rect -32 1863 2 1885
rect -32 1795 2 1813
rect -32 1727 2 1741
rect -32 1659 2 1669
rect -32 1591 2 1597
rect -32 1523 2 1525
rect -32 1487 2 1489
rect -32 1415 2 1421
rect -32 1343 2 1353
rect -32 1271 2 1285
rect -32 1199 2 1217
rect -32 1127 2 1149
rect -32 1055 2 1081
rect -32 983 2 1013
rect -32 902 2 945
rect 56 2067 90 2110
rect 56 1999 90 2029
rect 56 1931 90 1957
rect 56 1863 90 1885
rect 56 1795 90 1813
rect 56 1727 90 1741
rect 56 1659 90 1669
rect 56 1591 90 1597
rect 56 1523 90 1525
rect 56 1487 90 1489
rect 56 1415 90 1421
rect 56 1343 90 1353
rect 56 1271 90 1285
rect 56 1199 90 1217
rect 56 1127 90 1149
rect 56 1055 90 1081
rect 56 983 90 1013
rect 56 902 90 945
rect 144 2067 178 2110
rect 144 1999 178 2029
rect 144 1931 178 1957
rect 144 1863 178 1885
rect 144 1795 178 1813
rect 144 1727 178 1741
rect 144 1659 178 1669
rect 144 1591 178 1597
rect 144 1523 178 1525
rect 144 1487 178 1489
rect 144 1415 178 1421
rect 144 1343 178 1353
rect 144 1271 178 1285
rect 144 1199 178 1217
rect 144 1127 178 1149
rect 144 1055 178 1081
rect 144 983 178 1013
rect 144 902 178 945
rect 232 2067 266 2110
rect 232 1999 266 2029
rect 232 1931 266 1957
rect 232 1863 266 1885
rect 232 1795 266 1813
rect 232 1727 266 1741
rect 232 1659 266 1669
rect 232 1591 266 1597
rect 232 1523 266 1525
rect 232 1487 266 1489
rect 232 1415 266 1421
rect 232 1343 266 1353
rect 232 1271 266 1285
rect 232 1199 266 1217
rect 232 1127 266 1149
rect 232 1055 266 1081
rect 232 983 266 1013
rect 232 902 266 945
rect 320 2067 354 2110
rect 320 1999 354 2029
rect 320 1931 354 1957
rect 320 1863 354 1885
rect 320 1795 354 1813
rect 320 1727 354 1741
rect 320 1659 354 1669
rect 320 1591 354 1597
rect 320 1523 354 1525
rect 320 1487 354 1489
rect 320 1415 354 1421
rect 320 1343 354 1353
rect 320 1271 354 1285
rect 320 1199 354 1217
rect 320 1127 354 1149
rect 320 1055 354 1081
rect 320 983 354 1013
rect 320 902 354 945
rect 2715 1973 3097 2293
rect 2715 1939 2734 1973
rect 2768 1939 3097 1973
rect 2715 1905 3097 1939
rect 2715 1871 2734 1905
rect 2768 1871 3097 1905
rect 2715 1837 3097 1871
rect 2715 1803 2734 1837
rect 2768 1803 3097 1837
rect 2715 1769 3097 1803
rect 2715 1735 2734 1769
rect 2768 1735 3097 1769
rect 2715 1701 3097 1735
rect 2715 1667 2734 1701
rect 2768 1667 3097 1701
rect 2715 1633 3097 1667
rect 2715 1599 2734 1633
rect 2768 1599 3097 1633
rect 2715 1565 3097 1599
rect 2715 1531 2734 1565
rect 2768 1531 3097 1565
rect 2715 1497 3097 1531
rect 2715 1463 2734 1497
rect 2768 1485 3097 1497
rect 2768 1463 3152 1485
rect 2715 1429 3152 1463
rect 2715 1395 2734 1429
rect 2768 1395 3152 1429
rect 2715 1361 3152 1395
rect 2715 1327 2734 1361
rect 2768 1327 3152 1361
rect 2715 1293 3152 1327
rect 2715 1259 2734 1293
rect 2768 1259 3152 1293
rect 2715 1225 3152 1259
rect 2715 1191 2734 1225
rect 2768 1191 3152 1225
rect 3921 1207 5740 1993
rect 2715 1157 3152 1191
rect 2715 1123 2734 1157
rect 2768 1123 3152 1157
rect 2715 1089 3152 1123
rect 2715 1055 2734 1089
rect 2768 1055 3152 1089
rect 2715 1021 3152 1055
rect 2715 987 2734 1021
rect 2768 987 3152 1021
rect 2715 953 3152 987
rect 2715 919 2734 953
rect 2768 919 3152 953
rect 2715 910 3152 919
rect -1885 848 -1612 878
rect -1685 437 -1612 848
rect 2715 885 2788 910
rect 2715 851 2734 885
rect 2768 851 2788 885
rect 2715 817 2788 851
rect -1306 778 220 796
rect -1306 744 -1273 778
rect -1233 744 -1201 778
rect -1165 744 -1131 778
rect -1095 744 -1063 778
rect -1023 744 -995 778
rect -951 744 -927 778
rect -879 744 -859 778
rect -807 744 -791 778
rect -735 744 -723 778
rect -663 744 -655 778
rect -591 744 -587 778
rect -485 744 -481 778
rect -417 744 -409 778
rect -349 744 -337 778
rect -281 744 -265 778
rect -213 744 -193 778
rect -145 744 -121 778
rect -77 744 -49 778
rect -9 744 23 778
rect 59 744 93 778
rect 129 744 161 778
rect 201 744 220 778
rect -1306 726 220 744
rect 870 778 2396 796
rect 870 744 889 778
rect 929 744 961 778
rect 997 744 1031 778
rect 1067 744 1099 778
rect 1139 744 1167 778
rect 1211 744 1235 778
rect 1283 744 1303 778
rect 1355 744 1371 778
rect 1427 744 1439 778
rect 1499 744 1507 778
rect 1571 744 1575 778
rect 1677 744 1681 778
rect 1745 744 1753 778
rect 1813 744 1825 778
rect 1881 744 1897 778
rect 1949 744 1969 778
rect 2017 744 2041 778
rect 2085 744 2113 778
rect 2153 744 2185 778
rect 2221 744 2255 778
rect 2291 744 2323 778
rect 2363 744 2396 778
rect 870 726 2396 744
rect 2715 783 2734 817
rect 2768 783 2788 817
rect 2715 437 2788 783
rect -1685 435 2788 437
rect -1685 333 -1454 435
rect 2524 333 2788 435
rect -1685 332 2788 333
<< viali >>
rect -1352 2208 -1342 2242
rect -1342 2208 -1318 2242
rect -1280 2208 -1274 2242
rect -1274 2208 -1246 2242
rect -1208 2208 -1206 2242
rect -1206 2208 -1174 2242
rect -1136 2208 -1104 2242
rect -1104 2208 -1102 2242
rect -1064 2208 -1036 2242
rect -1036 2208 -1030 2242
rect -992 2208 -968 2242
rect -968 2208 -958 2242
rect -920 2208 -900 2242
rect -900 2208 -886 2242
rect -848 2208 -832 2242
rect -832 2208 -814 2242
rect -776 2208 -764 2242
rect -764 2208 -742 2242
rect -704 2208 -696 2242
rect -696 2208 -670 2242
rect -632 2208 -628 2242
rect -628 2208 -598 2242
rect -560 2208 -526 2242
rect -488 2208 -458 2242
rect -458 2208 -454 2242
rect -416 2208 -390 2242
rect -390 2208 -382 2242
rect -344 2208 -322 2242
rect -322 2208 -310 2242
rect -272 2208 -254 2242
rect -254 2208 -238 2242
rect -200 2208 -186 2242
rect -186 2208 -166 2242
rect -128 2208 -118 2242
rect -118 2208 -94 2242
rect -56 2208 -50 2242
rect -50 2208 -22 2242
rect 16 2208 18 2242
rect 18 2208 50 2242
rect 88 2208 120 2242
rect 120 2208 122 2242
rect 160 2208 188 2242
rect 188 2208 194 2242
rect 232 2208 256 2242
rect 256 2208 266 2242
rect 824 2208 834 2242
rect 834 2208 858 2242
rect 896 2208 902 2242
rect 902 2208 930 2242
rect 968 2208 970 2242
rect 970 2208 1002 2242
rect 1040 2208 1072 2242
rect 1072 2208 1074 2242
rect 1112 2208 1140 2242
rect 1140 2208 1146 2242
rect 1184 2208 1208 2242
rect 1208 2208 1218 2242
rect 1256 2208 1276 2242
rect 1276 2208 1290 2242
rect 1328 2208 1344 2242
rect 1344 2208 1362 2242
rect 1400 2208 1412 2242
rect 1412 2208 1434 2242
rect 1472 2208 1480 2242
rect 1480 2208 1506 2242
rect 1544 2208 1548 2242
rect 1548 2208 1578 2242
rect 1616 2208 1650 2242
rect 1688 2208 1718 2242
rect 1718 2208 1722 2242
rect 1760 2208 1786 2242
rect 1786 2208 1794 2242
rect 1832 2208 1854 2242
rect 1854 2208 1866 2242
rect 1904 2208 1922 2242
rect 1922 2208 1938 2242
rect 1976 2208 1990 2242
rect 1990 2208 2010 2242
rect 2048 2208 2058 2242
rect 2058 2208 2082 2242
rect 2120 2208 2126 2242
rect 2126 2208 2154 2242
rect 2192 2208 2194 2242
rect 2194 2208 2226 2242
rect 2264 2208 2296 2242
rect 2296 2208 2298 2242
rect 2336 2208 2364 2242
rect 2364 2208 2370 2242
rect 2408 2208 2432 2242
rect 2432 2208 2442 2242
rect -5777 2074 -5743 2108
rect -5705 2074 -5671 2108
rect -5633 2074 -5599 2108
rect -5561 2074 -5527 2108
rect -5489 2074 -5455 2108
rect -5417 2074 -5383 2108
rect -2346 2074 -2312 2108
rect -2274 2074 -2240 2108
rect -2202 2074 -2168 2108
rect -2130 2074 -2096 2108
rect -2058 2074 -2024 2108
rect -1986 2074 -1952 2108
rect -5782 1565 -5748 1599
rect -5710 1565 -5676 1599
rect -5638 1565 -5604 1599
rect -5566 1565 -5532 1599
rect -5494 1565 -5460 1599
rect -5422 1565 -5388 1599
rect -2351 1565 -2317 1599
rect -2279 1565 -2245 1599
rect -2207 1565 -2173 1599
rect -2135 1565 -2101 1599
rect -2063 1565 -2029 1599
rect -1991 1565 -1957 1599
rect -5821 1026 -5787 1060
rect -5749 1026 -5715 1060
rect -5677 1026 -5643 1060
rect -5605 1026 -5571 1060
rect -5533 1026 -5499 1060
rect -5461 1026 -5427 1060
rect -2390 1026 -2356 1060
rect -2318 1026 -2284 1060
rect -2246 1026 -2212 1060
rect -2174 1026 -2140 1060
rect -2102 1026 -2068 1060
rect -2030 1026 -1996 1060
rect -1440 2033 -1406 2063
rect -1440 2029 -1406 2033
rect -1440 1965 -1406 1991
rect -1440 1957 -1406 1965
rect -1440 1897 -1406 1919
rect -1440 1885 -1406 1897
rect -1440 1829 -1406 1847
rect -1440 1813 -1406 1829
rect -1440 1761 -1406 1775
rect -1440 1741 -1406 1761
rect -1440 1693 -1406 1703
rect -1440 1669 -1406 1693
rect -1440 1625 -1406 1631
rect -1440 1597 -1406 1625
rect -1440 1557 -1406 1559
rect -1440 1525 -1406 1557
rect -1440 1455 -1406 1487
rect -1440 1453 -1406 1455
rect -1440 1387 -1406 1415
rect -1440 1381 -1406 1387
rect -1440 1319 -1406 1343
rect -1440 1309 -1406 1319
rect -1440 1251 -1406 1271
rect -1440 1237 -1406 1251
rect -1440 1183 -1406 1199
rect -1440 1165 -1406 1183
rect -1440 1115 -1406 1127
rect -1440 1093 -1406 1115
rect -1440 1047 -1406 1055
rect -1440 1021 -1406 1047
rect -1440 979 -1406 983
rect -1440 949 -1406 979
rect -1352 2033 -1318 2063
rect -1352 2029 -1318 2033
rect -1352 1965 -1318 1991
rect -1352 1957 -1318 1965
rect -1352 1897 -1318 1919
rect -1352 1885 -1318 1897
rect -1352 1829 -1318 1847
rect -1352 1813 -1318 1829
rect -1352 1761 -1318 1775
rect -1352 1741 -1318 1761
rect -1352 1693 -1318 1703
rect -1352 1669 -1318 1693
rect -1352 1625 -1318 1631
rect -1352 1597 -1318 1625
rect -1352 1557 -1318 1559
rect -1352 1525 -1318 1557
rect -1352 1455 -1318 1487
rect -1352 1453 -1318 1455
rect -1352 1387 -1318 1415
rect -1352 1381 -1318 1387
rect -1352 1319 -1318 1343
rect -1352 1309 -1318 1319
rect -1352 1251 -1318 1271
rect -1352 1237 -1318 1251
rect -1352 1183 -1318 1199
rect -1352 1165 -1318 1183
rect -1352 1115 -1318 1127
rect -1352 1093 -1318 1115
rect -1352 1047 -1318 1055
rect -1352 1021 -1318 1047
rect -1352 979 -1318 983
rect -1352 949 -1318 979
rect -1264 2033 -1230 2063
rect -1264 2029 -1230 2033
rect -1264 1965 -1230 1991
rect -1264 1957 -1230 1965
rect -1264 1897 -1230 1919
rect -1264 1885 -1230 1897
rect -1264 1829 -1230 1847
rect -1264 1813 -1230 1829
rect -1264 1761 -1230 1775
rect -1264 1741 -1230 1761
rect -1264 1693 -1230 1703
rect -1264 1669 -1230 1693
rect -1264 1625 -1230 1631
rect -1264 1597 -1230 1625
rect -1264 1557 -1230 1559
rect -1264 1525 -1230 1557
rect -1264 1455 -1230 1487
rect -1264 1453 -1230 1455
rect -1264 1387 -1230 1415
rect -1264 1381 -1230 1387
rect -1264 1319 -1230 1343
rect -1264 1309 -1230 1319
rect -1264 1251 -1230 1271
rect -1264 1237 -1230 1251
rect -1264 1183 -1230 1199
rect -1264 1165 -1230 1183
rect -1264 1115 -1230 1127
rect -1264 1093 -1230 1115
rect -1264 1047 -1230 1055
rect -1264 1021 -1230 1047
rect -1264 979 -1230 983
rect -1264 949 -1230 979
rect -1176 2033 -1142 2063
rect -1176 2029 -1142 2033
rect -1176 1965 -1142 1991
rect -1176 1957 -1142 1965
rect -1176 1897 -1142 1919
rect -1176 1885 -1142 1897
rect -1176 1829 -1142 1847
rect -1176 1813 -1142 1829
rect -1176 1761 -1142 1775
rect -1176 1741 -1142 1761
rect -1176 1693 -1142 1703
rect -1176 1669 -1142 1693
rect -1176 1625 -1142 1631
rect -1176 1597 -1142 1625
rect -1176 1557 -1142 1559
rect -1176 1525 -1142 1557
rect -1176 1455 -1142 1487
rect -1176 1453 -1142 1455
rect -1176 1387 -1142 1415
rect -1176 1381 -1142 1387
rect -1176 1319 -1142 1343
rect -1176 1309 -1142 1319
rect -1176 1251 -1142 1271
rect -1176 1237 -1142 1251
rect -1176 1183 -1142 1199
rect -1176 1165 -1142 1183
rect -1176 1115 -1142 1127
rect -1176 1093 -1142 1115
rect -1176 1047 -1142 1055
rect -1176 1021 -1142 1047
rect -1176 979 -1142 983
rect -1176 949 -1142 979
rect -1088 2033 -1054 2063
rect -1088 2029 -1054 2033
rect -1088 1965 -1054 1991
rect -1088 1957 -1054 1965
rect -1088 1897 -1054 1919
rect -1088 1885 -1054 1897
rect -1088 1829 -1054 1847
rect -1088 1813 -1054 1829
rect -1088 1761 -1054 1775
rect -1088 1741 -1054 1761
rect -1088 1693 -1054 1703
rect -1088 1669 -1054 1693
rect -1088 1625 -1054 1631
rect -1088 1597 -1054 1625
rect -1088 1557 -1054 1559
rect -1088 1525 -1054 1557
rect -1088 1455 -1054 1487
rect -1088 1453 -1054 1455
rect -1088 1387 -1054 1415
rect -1088 1381 -1054 1387
rect -1088 1319 -1054 1343
rect -1088 1309 -1054 1319
rect -1088 1251 -1054 1271
rect -1088 1237 -1054 1251
rect -1088 1183 -1054 1199
rect -1088 1165 -1054 1183
rect -1088 1115 -1054 1127
rect -1088 1093 -1054 1115
rect -1088 1047 -1054 1055
rect -1088 1021 -1054 1047
rect -1088 979 -1054 983
rect -1088 949 -1054 979
rect -1000 2033 -966 2063
rect -1000 2029 -966 2033
rect -1000 1965 -966 1991
rect -1000 1957 -966 1965
rect -1000 1897 -966 1919
rect -1000 1885 -966 1897
rect -1000 1829 -966 1847
rect -1000 1813 -966 1829
rect -1000 1761 -966 1775
rect -1000 1741 -966 1761
rect -1000 1693 -966 1703
rect -1000 1669 -966 1693
rect -1000 1625 -966 1631
rect -1000 1597 -966 1625
rect -1000 1557 -966 1559
rect -1000 1525 -966 1557
rect -1000 1455 -966 1487
rect -1000 1453 -966 1455
rect -1000 1387 -966 1415
rect -1000 1381 -966 1387
rect -1000 1319 -966 1343
rect -1000 1309 -966 1319
rect -1000 1251 -966 1271
rect -1000 1237 -966 1251
rect -1000 1183 -966 1199
rect -1000 1165 -966 1183
rect -1000 1115 -966 1127
rect -1000 1093 -966 1115
rect -1000 1047 -966 1055
rect -1000 1021 -966 1047
rect -1000 979 -966 983
rect -1000 949 -966 979
rect -912 2033 -878 2063
rect -912 2029 -878 2033
rect -912 1965 -878 1991
rect -912 1957 -878 1965
rect -912 1897 -878 1919
rect -912 1885 -878 1897
rect -912 1829 -878 1847
rect -912 1813 -878 1829
rect -912 1761 -878 1775
rect -912 1741 -878 1761
rect -912 1693 -878 1703
rect -912 1669 -878 1693
rect -912 1625 -878 1631
rect -912 1597 -878 1625
rect -912 1557 -878 1559
rect -912 1525 -878 1557
rect -912 1455 -878 1487
rect -912 1453 -878 1455
rect -912 1387 -878 1415
rect -912 1381 -878 1387
rect -912 1319 -878 1343
rect -912 1309 -878 1319
rect -912 1251 -878 1271
rect -912 1237 -878 1251
rect -912 1183 -878 1199
rect -912 1165 -878 1183
rect -912 1115 -878 1127
rect -912 1093 -878 1115
rect -912 1047 -878 1055
rect -912 1021 -878 1047
rect -912 979 -878 983
rect -912 949 -878 979
rect -824 2033 -790 2063
rect -824 2029 -790 2033
rect -824 1965 -790 1991
rect -824 1957 -790 1965
rect -824 1897 -790 1919
rect -824 1885 -790 1897
rect -824 1829 -790 1847
rect -824 1813 -790 1829
rect -824 1761 -790 1775
rect -824 1741 -790 1761
rect -824 1693 -790 1703
rect -824 1669 -790 1693
rect -824 1625 -790 1631
rect -824 1597 -790 1625
rect -824 1557 -790 1559
rect -824 1525 -790 1557
rect -824 1455 -790 1487
rect -824 1453 -790 1455
rect -824 1387 -790 1415
rect -824 1381 -790 1387
rect -824 1319 -790 1343
rect -824 1309 -790 1319
rect -824 1251 -790 1271
rect -824 1237 -790 1251
rect -824 1183 -790 1199
rect -824 1165 -790 1183
rect -824 1115 -790 1127
rect -824 1093 -790 1115
rect -824 1047 -790 1055
rect -824 1021 -790 1047
rect -824 979 -790 983
rect -824 949 -790 979
rect -736 2033 -702 2063
rect -736 2029 -702 2033
rect -736 1965 -702 1991
rect -736 1957 -702 1965
rect -736 1897 -702 1919
rect -736 1885 -702 1897
rect -736 1829 -702 1847
rect -736 1813 -702 1829
rect -736 1761 -702 1775
rect -736 1741 -702 1761
rect -736 1693 -702 1703
rect -736 1669 -702 1693
rect -736 1625 -702 1631
rect -736 1597 -702 1625
rect -736 1557 -702 1559
rect -736 1525 -702 1557
rect -736 1455 -702 1487
rect -736 1453 -702 1455
rect -736 1387 -702 1415
rect -736 1381 -702 1387
rect -736 1319 -702 1343
rect -736 1309 -702 1319
rect -736 1251 -702 1271
rect -736 1237 -702 1251
rect -736 1183 -702 1199
rect -736 1165 -702 1183
rect -736 1115 -702 1127
rect -736 1093 -702 1115
rect -736 1047 -702 1055
rect -736 1021 -702 1047
rect -736 979 -702 983
rect -736 949 -702 979
rect -648 2033 -614 2063
rect -648 2029 -614 2033
rect -648 1965 -614 1991
rect -648 1957 -614 1965
rect -648 1897 -614 1919
rect -648 1885 -614 1897
rect -648 1829 -614 1847
rect -648 1813 -614 1829
rect -648 1761 -614 1775
rect -648 1741 -614 1761
rect -648 1693 -614 1703
rect -648 1669 -614 1693
rect -648 1625 -614 1631
rect -648 1597 -614 1625
rect -648 1557 -614 1559
rect -648 1525 -614 1557
rect -648 1455 -614 1487
rect -648 1453 -614 1455
rect -648 1387 -614 1415
rect -648 1381 -614 1387
rect -648 1319 -614 1343
rect -648 1309 -614 1319
rect -648 1251 -614 1271
rect -648 1237 -614 1251
rect -648 1183 -614 1199
rect -648 1165 -614 1183
rect -648 1115 -614 1127
rect -648 1093 -614 1115
rect -648 1047 -614 1055
rect -648 1021 -614 1047
rect -648 979 -614 983
rect -648 949 -614 979
rect -560 2033 -526 2063
rect -560 2029 -526 2033
rect -560 1965 -526 1991
rect -560 1957 -526 1965
rect -560 1897 -526 1919
rect -560 1885 -526 1897
rect -560 1829 -526 1847
rect -560 1813 -526 1829
rect -560 1761 -526 1775
rect -560 1741 -526 1761
rect -560 1693 -526 1703
rect -560 1669 -526 1693
rect -560 1625 -526 1631
rect -560 1597 -526 1625
rect -560 1557 -526 1559
rect -560 1525 -526 1557
rect -560 1455 -526 1487
rect -560 1453 -526 1455
rect -560 1387 -526 1415
rect -560 1381 -526 1387
rect -560 1319 -526 1343
rect -560 1309 -526 1319
rect -560 1251 -526 1271
rect -560 1237 -526 1251
rect -560 1183 -526 1199
rect -560 1165 -526 1183
rect -560 1115 -526 1127
rect -560 1093 -526 1115
rect -560 1047 -526 1055
rect -560 1021 -526 1047
rect -560 979 -526 983
rect -560 949 -526 979
rect -472 2033 -438 2063
rect -472 2029 -438 2033
rect -472 1965 -438 1991
rect -472 1957 -438 1965
rect -472 1897 -438 1919
rect -472 1885 -438 1897
rect -472 1829 -438 1847
rect -472 1813 -438 1829
rect -472 1761 -438 1775
rect -472 1741 -438 1761
rect -472 1693 -438 1703
rect -472 1669 -438 1693
rect -472 1625 -438 1631
rect -472 1597 -438 1625
rect -472 1557 -438 1559
rect -472 1525 -438 1557
rect -472 1455 -438 1487
rect -472 1453 -438 1455
rect -472 1387 -438 1415
rect -472 1381 -438 1387
rect -472 1319 -438 1343
rect -472 1309 -438 1319
rect -472 1251 -438 1271
rect -472 1237 -438 1251
rect -472 1183 -438 1199
rect -472 1165 -438 1183
rect -472 1115 -438 1127
rect -472 1093 -438 1115
rect -472 1047 -438 1055
rect -472 1021 -438 1047
rect -472 979 -438 983
rect -472 949 -438 979
rect -384 2033 -350 2063
rect -384 2029 -350 2033
rect -384 1965 -350 1991
rect -384 1957 -350 1965
rect -384 1897 -350 1919
rect -384 1885 -350 1897
rect -384 1829 -350 1847
rect -384 1813 -350 1829
rect -384 1761 -350 1775
rect -384 1741 -350 1761
rect -384 1693 -350 1703
rect -384 1669 -350 1693
rect -384 1625 -350 1631
rect -384 1597 -350 1625
rect -384 1557 -350 1559
rect -384 1525 -350 1557
rect -384 1455 -350 1487
rect -384 1453 -350 1455
rect -384 1387 -350 1415
rect -384 1381 -350 1387
rect -384 1319 -350 1343
rect -384 1309 -350 1319
rect -384 1251 -350 1271
rect -384 1237 -350 1251
rect -384 1183 -350 1199
rect -384 1165 -350 1183
rect -384 1115 -350 1127
rect -384 1093 -350 1115
rect -384 1047 -350 1055
rect -384 1021 -350 1047
rect -384 979 -350 983
rect -384 949 -350 979
rect -296 2033 -262 2063
rect -296 2029 -262 2033
rect -296 1965 -262 1991
rect -296 1957 -262 1965
rect -296 1897 -262 1919
rect -296 1885 -262 1897
rect -296 1829 -262 1847
rect -296 1813 -262 1829
rect -296 1761 -262 1775
rect -296 1741 -262 1761
rect -296 1693 -262 1703
rect -296 1669 -262 1693
rect -296 1625 -262 1631
rect -296 1597 -262 1625
rect -296 1557 -262 1559
rect -296 1525 -262 1557
rect -296 1455 -262 1487
rect -296 1453 -262 1455
rect -296 1387 -262 1415
rect -296 1381 -262 1387
rect -296 1319 -262 1343
rect -296 1309 -262 1319
rect -296 1251 -262 1271
rect -296 1237 -262 1251
rect -296 1183 -262 1199
rect -296 1165 -262 1183
rect -296 1115 -262 1127
rect -296 1093 -262 1115
rect -296 1047 -262 1055
rect -296 1021 -262 1047
rect -296 979 -262 983
rect -296 949 -262 979
rect -208 2033 -174 2063
rect -208 2029 -174 2033
rect -208 1965 -174 1991
rect -208 1957 -174 1965
rect -208 1897 -174 1919
rect -208 1885 -174 1897
rect -208 1829 -174 1847
rect -208 1813 -174 1829
rect -208 1761 -174 1775
rect -208 1741 -174 1761
rect -208 1693 -174 1703
rect -208 1669 -174 1693
rect -208 1625 -174 1631
rect -208 1597 -174 1625
rect -208 1557 -174 1559
rect -208 1525 -174 1557
rect -208 1455 -174 1487
rect -208 1453 -174 1455
rect -208 1387 -174 1415
rect -208 1381 -174 1387
rect -208 1319 -174 1343
rect -208 1309 -174 1319
rect -208 1251 -174 1271
rect -208 1237 -174 1251
rect -208 1183 -174 1199
rect -208 1165 -174 1183
rect -208 1115 -174 1127
rect -208 1093 -174 1115
rect -208 1047 -174 1055
rect -208 1021 -174 1047
rect -208 979 -174 983
rect -208 949 -174 979
rect -120 2033 -86 2063
rect -120 2029 -86 2033
rect -120 1965 -86 1991
rect -120 1957 -86 1965
rect -120 1897 -86 1919
rect -120 1885 -86 1897
rect -120 1829 -86 1847
rect -120 1813 -86 1829
rect -120 1761 -86 1775
rect -120 1741 -86 1761
rect -120 1693 -86 1703
rect -120 1669 -86 1693
rect -120 1625 -86 1631
rect -120 1597 -86 1625
rect -120 1557 -86 1559
rect -120 1525 -86 1557
rect -120 1455 -86 1487
rect -120 1453 -86 1455
rect -120 1387 -86 1415
rect -120 1381 -86 1387
rect -120 1319 -86 1343
rect -120 1309 -86 1319
rect -120 1251 -86 1271
rect -120 1237 -86 1251
rect -120 1183 -86 1199
rect -120 1165 -86 1183
rect -120 1115 -86 1127
rect -120 1093 -86 1115
rect -120 1047 -86 1055
rect -120 1021 -86 1047
rect -120 979 -86 983
rect -120 949 -86 979
rect -32 2033 2 2063
rect -32 2029 2 2033
rect -32 1965 2 1991
rect -32 1957 2 1965
rect -32 1897 2 1919
rect -32 1885 2 1897
rect -32 1829 2 1847
rect -32 1813 2 1829
rect -32 1761 2 1775
rect -32 1741 2 1761
rect -32 1693 2 1703
rect -32 1669 2 1693
rect -32 1625 2 1631
rect -32 1597 2 1625
rect -32 1557 2 1559
rect -32 1525 2 1557
rect -32 1455 2 1487
rect -32 1453 2 1455
rect -32 1387 2 1415
rect -32 1381 2 1387
rect -32 1319 2 1343
rect -32 1309 2 1319
rect -32 1251 2 1271
rect -32 1237 2 1251
rect -32 1183 2 1199
rect -32 1165 2 1183
rect -32 1115 2 1127
rect -32 1093 2 1115
rect -32 1047 2 1055
rect -32 1021 2 1047
rect -32 979 2 983
rect -32 949 2 979
rect 56 2033 90 2063
rect 56 2029 90 2033
rect 56 1965 90 1991
rect 56 1957 90 1965
rect 56 1897 90 1919
rect 56 1885 90 1897
rect 56 1829 90 1847
rect 56 1813 90 1829
rect 56 1761 90 1775
rect 56 1741 90 1761
rect 56 1693 90 1703
rect 56 1669 90 1693
rect 56 1625 90 1631
rect 56 1597 90 1625
rect 56 1557 90 1559
rect 56 1525 90 1557
rect 56 1455 90 1487
rect 56 1453 90 1455
rect 56 1387 90 1415
rect 56 1381 90 1387
rect 56 1319 90 1343
rect 56 1309 90 1319
rect 56 1251 90 1271
rect 56 1237 90 1251
rect 56 1183 90 1199
rect 56 1165 90 1183
rect 56 1115 90 1127
rect 56 1093 90 1115
rect 56 1047 90 1055
rect 56 1021 90 1047
rect 56 979 90 983
rect 56 949 90 979
rect 144 2033 178 2063
rect 144 2029 178 2033
rect 144 1965 178 1991
rect 144 1957 178 1965
rect 144 1897 178 1919
rect 144 1885 178 1897
rect 144 1829 178 1847
rect 144 1813 178 1829
rect 144 1761 178 1775
rect 144 1741 178 1761
rect 144 1693 178 1703
rect 144 1669 178 1693
rect 144 1625 178 1631
rect 144 1597 178 1625
rect 144 1557 178 1559
rect 144 1525 178 1557
rect 144 1455 178 1487
rect 144 1453 178 1455
rect 144 1387 178 1415
rect 144 1381 178 1387
rect 144 1319 178 1343
rect 144 1309 178 1319
rect 144 1251 178 1271
rect 144 1237 178 1251
rect 144 1183 178 1199
rect 144 1165 178 1183
rect 144 1115 178 1127
rect 144 1093 178 1115
rect 144 1047 178 1055
rect 144 1021 178 1047
rect 144 979 178 983
rect 144 949 178 979
rect 232 2033 266 2063
rect 232 2029 266 2033
rect 232 1965 266 1991
rect 232 1957 266 1965
rect 232 1897 266 1919
rect 232 1885 266 1897
rect 232 1829 266 1847
rect 232 1813 266 1829
rect 232 1761 266 1775
rect 232 1741 266 1761
rect 232 1693 266 1703
rect 232 1669 266 1693
rect 232 1625 266 1631
rect 232 1597 266 1625
rect 232 1557 266 1559
rect 232 1525 266 1557
rect 232 1455 266 1487
rect 232 1453 266 1455
rect 232 1387 266 1415
rect 232 1381 266 1387
rect 232 1319 266 1343
rect 232 1309 266 1319
rect 232 1251 266 1271
rect 232 1237 266 1251
rect 232 1183 266 1199
rect 232 1165 266 1183
rect 232 1115 266 1127
rect 232 1093 266 1115
rect 232 1047 266 1055
rect 232 1021 266 1047
rect 232 979 266 983
rect 232 949 266 979
rect 320 2033 354 2063
rect 320 2029 354 2033
rect 320 1965 354 1991
rect 320 1957 354 1965
rect 320 1897 354 1919
rect 320 1885 354 1897
rect 320 1829 354 1847
rect 320 1813 354 1829
rect 320 1761 354 1775
rect 320 1741 354 1761
rect 320 1693 354 1703
rect 320 1669 354 1693
rect 320 1625 354 1631
rect 320 1597 354 1625
rect 320 1557 354 1559
rect 320 1525 354 1557
rect 320 1455 354 1487
rect 320 1453 354 1455
rect 320 1387 354 1415
rect 320 1381 354 1387
rect 320 1319 354 1343
rect 320 1309 354 1319
rect 320 1251 354 1271
rect 320 1237 354 1251
rect 320 1183 354 1199
rect 320 1165 354 1183
rect 320 1115 354 1127
rect 320 1093 354 1115
rect 320 1047 354 1055
rect 320 1021 354 1047
rect 320 979 354 983
rect 320 949 354 979
rect -1273 744 -1267 778
rect -1267 744 -1239 778
rect -1201 744 -1199 778
rect -1199 744 -1167 778
rect -1129 744 -1097 778
rect -1097 744 -1095 778
rect -1057 744 -1029 778
rect -1029 744 -1023 778
rect -985 744 -961 778
rect -961 744 -951 778
rect -913 744 -893 778
rect -893 744 -879 778
rect -841 744 -825 778
rect -825 744 -807 778
rect -769 744 -757 778
rect -757 744 -735 778
rect -697 744 -689 778
rect -689 744 -663 778
rect -625 744 -621 778
rect -621 744 -591 778
rect -553 744 -519 778
rect -481 744 -451 778
rect -451 744 -447 778
rect -409 744 -383 778
rect -383 744 -375 778
rect -337 744 -315 778
rect -315 744 -303 778
rect -265 744 -247 778
rect -247 744 -231 778
rect -193 744 -179 778
rect -179 744 -159 778
rect -121 744 -111 778
rect -111 744 -87 778
rect -49 744 -43 778
rect -43 744 -15 778
rect 23 744 25 778
rect 25 744 57 778
rect 95 744 127 778
rect 127 744 129 778
rect 167 744 195 778
rect 195 744 201 778
rect 889 744 895 778
rect 895 744 923 778
rect 961 744 963 778
rect 963 744 995 778
rect 1033 744 1065 778
rect 1065 744 1067 778
rect 1105 744 1133 778
rect 1133 744 1139 778
rect 1177 744 1201 778
rect 1201 744 1211 778
rect 1249 744 1269 778
rect 1269 744 1283 778
rect 1321 744 1337 778
rect 1337 744 1355 778
rect 1393 744 1405 778
rect 1405 744 1427 778
rect 1465 744 1473 778
rect 1473 744 1499 778
rect 1537 744 1541 778
rect 1541 744 1571 778
rect 1609 744 1643 778
rect 1681 744 1711 778
rect 1711 744 1715 778
rect 1753 744 1779 778
rect 1779 744 1787 778
rect 1825 744 1847 778
rect 1847 744 1859 778
rect 1897 744 1915 778
rect 1915 744 1931 778
rect 1969 744 1983 778
rect 1983 744 2003 778
rect 2041 744 2051 778
rect 2051 744 2075 778
rect 2113 744 2119 778
rect 2119 744 2147 778
rect 2185 744 2187 778
rect 2187 744 2219 778
rect 2257 744 2289 778
rect 2289 744 2291 778
rect 2329 744 2357 778
rect 2357 744 2363 778
<< metal1 >>
rect -2364 2242 308 2260
rect -2364 2208 -1352 2242
rect -1318 2208 -1280 2242
rect -1246 2208 -1208 2242
rect -1174 2208 -1136 2242
rect -1102 2208 -1064 2242
rect -1030 2208 -992 2242
rect -958 2208 -920 2242
rect -886 2208 -848 2242
rect -814 2208 -776 2242
rect -742 2208 -704 2242
rect -670 2208 -632 2242
rect -598 2208 -560 2242
rect -526 2208 -488 2242
rect -454 2208 -416 2242
rect -382 2208 -344 2242
rect -310 2208 -272 2242
rect -238 2208 -200 2242
rect -166 2208 -128 2242
rect -94 2208 -56 2242
rect -22 2208 16 2242
rect 50 2208 88 2242
rect 122 2208 160 2242
rect 194 2208 232 2242
rect 266 2208 308 2242
rect -2364 2190 308 2208
rect 782 2242 3635 2262
rect 782 2208 824 2242
rect 858 2208 896 2242
rect 930 2208 968 2242
rect 1002 2208 1040 2242
rect 1074 2208 1112 2242
rect 1146 2208 1184 2242
rect 1218 2208 1256 2242
rect 1290 2208 1328 2242
rect 1362 2208 1400 2242
rect 1434 2208 1472 2242
rect 1506 2208 1544 2242
rect 1578 2208 1616 2242
rect 1650 2208 1688 2242
rect 1722 2208 1760 2242
rect 1794 2208 1832 2242
rect 1866 2208 1904 2242
rect 1938 2208 1976 2242
rect 2010 2208 2048 2242
rect 2082 2208 2120 2242
rect 2154 2208 2192 2242
rect 2226 2208 2264 2242
rect 2298 2208 2336 2242
rect 2370 2208 2408 2242
rect 2442 2208 3635 2242
rect 782 2190 3635 2208
rect -5827 2116 -5374 2126
rect -5827 2108 -5369 2116
rect -5827 2074 -5777 2108
rect -5743 2074 -5705 2108
rect -5671 2074 -5633 2108
rect -5599 2074 -5561 2108
rect -5527 2074 -5489 2108
rect -5455 2074 -5417 2108
rect -5383 2074 -5369 2108
rect -5827 2066 -5369 2074
rect -2364 2108 -1932 2190
rect 2164 2189 3635 2190
rect -2364 2074 -2346 2108
rect -2312 2074 -2274 2108
rect -2240 2074 -2202 2108
rect -2168 2074 -2130 2108
rect -2096 2074 -2058 2108
rect -2024 2074 -1986 2108
rect -1952 2074 -1932 2108
rect -1446 2104 -1400 2106
rect -5827 1853 -5374 2066
rect -2364 2056 -1932 2074
rect -1557 2098 -1400 2104
rect -1557 2046 -1452 2098
rect -1557 2040 -1440 2046
rect -1446 2029 -1440 2040
rect -1406 2029 -1400 2046
rect -1446 1991 -1400 2029
rect -1446 1957 -1440 1991
rect -1406 1957 -1400 1991
rect -1446 1919 -1400 1957
rect -1446 1885 -1440 1919
rect -1406 1885 -1400 1919
rect -1358 2063 -1312 2106
rect -1358 2029 -1352 2063
rect -1318 2029 -1312 2063
rect -1358 1991 -1312 2029
rect -1358 1957 -1352 1991
rect -1318 1957 -1312 1991
rect -1358 1919 -1312 1957
rect -1358 1916 -1352 1919
rect -5827 1801 -5747 1853
rect -5695 1801 -5683 1853
rect -5631 1801 -5619 1853
rect -5567 1801 -5555 1853
rect -5503 1801 -5491 1853
rect -5439 1801 -5374 1853
rect -5827 1782 -5374 1801
rect -2370 1856 -1905 1878
rect -2370 1804 -2271 1856
rect -2219 1804 -2207 1856
rect -2155 1804 -2143 1856
rect -2091 1804 -2079 1856
rect -2027 1804 -2015 1856
rect -1963 1804 -1905 1856
rect -6207 1599 -5364 1657
rect -6207 1565 -5782 1599
rect -5748 1565 -5710 1599
rect -5676 1565 -5638 1599
rect -5604 1565 -5566 1599
rect -5532 1565 -5494 1599
rect -5460 1565 -5422 1599
rect -5388 1565 -5364 1599
rect -6207 1522 -5364 1565
rect -2370 1617 -1905 1804
rect -1446 1847 -1400 1885
rect -1364 1910 -1352 1916
rect -1318 1916 -1312 1919
rect -1270 2063 -1224 2106
rect -1270 2029 -1264 2063
rect -1230 2029 -1224 2063
rect -1270 1991 -1224 2029
rect -1270 1957 -1264 1991
rect -1230 1957 -1224 1991
rect -1270 1919 -1224 1957
rect -1318 1910 -1306 1916
rect -1312 1858 -1306 1910
rect -1364 1852 -1306 1858
rect -1270 1885 -1264 1919
rect -1230 1885 -1224 1919
rect -1182 2063 -1136 2106
rect -1094 2104 -1048 2106
rect -1182 2029 -1176 2063
rect -1142 2029 -1136 2063
rect -1106 2098 -1048 2104
rect -1106 2046 -1100 2098
rect -1106 2040 -1088 2046
rect -1182 1991 -1136 2029
rect -1182 1957 -1176 1991
rect -1142 1957 -1136 1991
rect -1182 1919 -1136 1957
rect -1182 1916 -1176 1919
rect -1446 1813 -1440 1847
rect -1406 1813 -1400 1847
rect -1446 1775 -1400 1813
rect -1446 1741 -1440 1775
rect -1406 1741 -1400 1775
rect -1446 1703 -1400 1741
rect -1446 1669 -1440 1703
rect -1406 1669 -1400 1703
rect -1446 1631 -1400 1669
rect -2370 1599 -1904 1617
rect -2370 1565 -2351 1599
rect -2317 1565 -2279 1599
rect -2245 1565 -2207 1599
rect -2173 1565 -2135 1599
rect -2101 1565 -2063 1599
rect -2029 1565 -1991 1599
rect -1957 1565 -1904 1599
rect -2370 1525 -1904 1565
rect -5841 1302 -5408 1328
rect -5841 1250 -5781 1302
rect -5729 1250 -5717 1302
rect -5665 1250 -5653 1302
rect -5601 1250 -5589 1302
rect -5537 1250 -5525 1302
rect -5473 1250 -5408 1302
rect -5841 1060 -5408 1250
rect -2369 1306 -1904 1525
rect -1446 1597 -1440 1631
rect -1406 1597 -1400 1631
rect -1446 1559 -1400 1597
rect -1446 1525 -1440 1559
rect -1406 1525 -1400 1559
rect -1446 1487 -1400 1525
rect -1446 1453 -1440 1487
rect -1406 1453 -1400 1487
rect -1446 1415 -1400 1453
rect -1446 1408 -1440 1415
rect -1458 1402 -1440 1408
rect -1406 1408 -1400 1415
rect -1358 1847 -1312 1852
rect -1358 1813 -1352 1847
rect -1318 1813 -1312 1847
rect -1358 1775 -1312 1813
rect -1358 1741 -1352 1775
rect -1318 1741 -1312 1775
rect -1358 1703 -1312 1741
rect -1358 1669 -1352 1703
rect -1318 1669 -1312 1703
rect -1358 1631 -1312 1669
rect -1270 1847 -1224 1885
rect -1188 1910 -1176 1916
rect -1142 1916 -1136 1919
rect -1094 2029 -1088 2040
rect -1054 2029 -1048 2046
rect -1094 1991 -1048 2029
rect -1094 1957 -1088 1991
rect -1054 1957 -1048 1991
rect -1094 1919 -1048 1957
rect -1142 1910 -1130 1916
rect -1136 1858 -1130 1910
rect -1188 1852 -1130 1858
rect -1094 1885 -1088 1919
rect -1054 1885 -1048 1919
rect -1006 2063 -960 2106
rect -1006 2029 -1000 2063
rect -966 2029 -960 2063
rect -1006 1991 -960 2029
rect -1006 1957 -1000 1991
rect -966 1957 -960 1991
rect -1006 1919 -960 1957
rect -1006 1916 -1000 1919
rect -1270 1813 -1264 1847
rect -1230 1813 -1224 1847
rect -1270 1775 -1224 1813
rect -1270 1741 -1264 1775
rect -1230 1741 -1224 1775
rect -1270 1703 -1224 1741
rect -1270 1669 -1264 1703
rect -1230 1669 -1224 1703
rect -1270 1650 -1224 1669
rect -1182 1847 -1136 1852
rect -1182 1813 -1176 1847
rect -1142 1813 -1136 1847
rect -1182 1775 -1136 1813
rect -1182 1741 -1176 1775
rect -1142 1741 -1136 1775
rect -1182 1703 -1136 1741
rect -1182 1669 -1176 1703
rect -1142 1669 -1136 1703
rect -1358 1597 -1352 1631
rect -1318 1597 -1312 1631
rect -1358 1559 -1312 1597
rect -1278 1644 -1214 1650
rect -1278 1592 -1272 1644
rect -1220 1592 -1214 1644
rect -1278 1586 -1214 1592
rect -1182 1631 -1136 1669
rect -1182 1597 -1176 1631
rect -1142 1597 -1136 1631
rect -1358 1525 -1352 1559
rect -1318 1525 -1312 1559
rect -1358 1487 -1312 1525
rect -1358 1453 -1352 1487
rect -1318 1453 -1312 1487
rect -1358 1415 -1312 1453
rect -1406 1402 -1394 1408
rect -1458 1350 -1452 1402
rect -1400 1350 -1394 1402
rect -1458 1344 -1394 1350
rect -1358 1381 -1352 1415
rect -1318 1381 -1312 1415
rect -2369 1254 -2272 1306
rect -2220 1254 -2208 1306
rect -2156 1254 -2144 1306
rect -2092 1254 -2080 1306
rect -2028 1254 -2016 1306
rect -1964 1254 -1904 1306
rect -2369 1232 -1904 1254
rect -1446 1343 -1400 1344
rect -1446 1309 -1440 1343
rect -1406 1309 -1400 1343
rect -1446 1271 -1400 1309
rect -1446 1237 -1440 1271
rect -1406 1237 -1400 1271
rect -1446 1199 -1400 1237
rect -1358 1343 -1312 1381
rect -1358 1309 -1352 1343
rect -1318 1309 -1312 1343
rect -1358 1271 -1312 1309
rect -1358 1237 -1352 1271
rect -1318 1237 -1312 1271
rect -1358 1218 -1312 1237
rect -1270 1559 -1224 1586
rect -1270 1525 -1264 1559
rect -1230 1525 -1224 1559
rect -1270 1487 -1224 1525
rect -1270 1453 -1264 1487
rect -1230 1453 -1224 1487
rect -1270 1415 -1224 1453
rect -1270 1381 -1264 1415
rect -1230 1381 -1224 1415
rect -1270 1343 -1224 1381
rect -1270 1309 -1264 1343
rect -1230 1309 -1224 1343
rect -1270 1271 -1224 1309
rect -1270 1237 -1264 1271
rect -1230 1237 -1224 1271
rect -1446 1165 -1440 1199
rect -1406 1165 -1400 1199
rect -1446 1127 -1400 1165
rect -1370 1212 -1306 1218
rect -1370 1160 -1364 1212
rect -1312 1160 -1306 1212
rect -1370 1154 -1306 1160
rect -1270 1199 -1224 1237
rect -1182 1559 -1136 1597
rect -1182 1525 -1176 1559
rect -1142 1525 -1136 1559
rect -1182 1487 -1136 1525
rect -1182 1453 -1176 1487
rect -1142 1453 -1136 1487
rect -1182 1415 -1136 1453
rect -1182 1381 -1176 1415
rect -1142 1381 -1136 1415
rect -1094 1847 -1048 1885
rect -1018 1910 -1000 1916
rect -966 1910 -960 1919
rect -1018 1858 -1012 1910
rect -1018 1852 -960 1858
rect -1094 1813 -1088 1847
rect -1054 1813 -1048 1847
rect -1094 1775 -1048 1813
rect -1094 1741 -1088 1775
rect -1054 1741 -1048 1775
rect -1094 1703 -1048 1741
rect -1094 1669 -1088 1703
rect -1054 1669 -1048 1703
rect -1094 1631 -1048 1669
rect -1094 1597 -1088 1631
rect -1054 1597 -1048 1631
rect -1094 1559 -1048 1597
rect -1094 1525 -1088 1559
rect -1054 1525 -1048 1559
rect -1094 1487 -1048 1525
rect -1094 1453 -1088 1487
rect -1054 1453 -1048 1487
rect -1094 1415 -1048 1453
rect -1094 1408 -1088 1415
rect -1182 1343 -1136 1381
rect -1106 1402 -1088 1408
rect -1054 1408 -1048 1415
rect -1006 1847 -960 1852
rect -1006 1813 -1000 1847
rect -966 1813 -960 1847
rect -1006 1775 -960 1813
rect -1006 1741 -1000 1775
rect -966 1741 -960 1775
rect -1006 1703 -960 1741
rect -1006 1669 -1000 1703
rect -966 1669 -960 1703
rect -1006 1631 -960 1669
rect -918 2063 -872 2106
rect -918 2029 -912 2063
rect -878 2029 -872 2063
rect -918 1991 -872 2029
rect -918 1957 -912 1991
rect -878 1957 -872 1991
rect -918 1919 -872 1957
rect -918 1885 -912 1919
rect -878 1885 -872 1919
rect -830 2063 -784 2106
rect -742 2104 -696 2106
rect -830 2029 -824 2063
rect -790 2029 -784 2063
rect -754 2098 -696 2104
rect -754 2046 -748 2098
rect -754 2040 -736 2046
rect -830 1991 -784 2029
rect -830 1957 -824 1991
rect -790 1957 -784 1991
rect -830 1919 -784 1957
rect -830 1916 -824 1919
rect -918 1847 -872 1885
rect -842 1910 -824 1916
rect -790 1910 -784 1919
rect -842 1858 -836 1910
rect -842 1852 -784 1858
rect -918 1813 -912 1847
rect -878 1813 -872 1847
rect -918 1775 -872 1813
rect -918 1741 -912 1775
rect -878 1741 -872 1775
rect -918 1703 -872 1741
rect -918 1669 -912 1703
rect -878 1669 -872 1703
rect -918 1650 -872 1669
rect -830 1847 -784 1852
rect -830 1813 -824 1847
rect -790 1813 -784 1847
rect -830 1775 -784 1813
rect -830 1741 -824 1775
rect -790 1741 -784 1775
rect -830 1703 -784 1741
rect -830 1669 -824 1703
rect -790 1669 -784 1703
rect -1006 1597 -1000 1631
rect -966 1597 -960 1631
rect -1006 1559 -960 1597
rect -926 1644 -862 1650
rect -926 1592 -920 1644
rect -868 1592 -862 1644
rect -926 1586 -862 1592
rect -830 1631 -784 1669
rect -830 1597 -824 1631
rect -790 1597 -784 1631
rect -1006 1525 -1000 1559
rect -966 1525 -960 1559
rect -1006 1487 -960 1525
rect -1006 1453 -1000 1487
rect -966 1453 -960 1487
rect -1006 1415 -960 1453
rect -1054 1402 -1042 1408
rect -1106 1350 -1100 1402
rect -1048 1350 -1042 1402
rect -1106 1344 -1042 1350
rect -1006 1381 -1000 1415
rect -966 1381 -960 1415
rect -1182 1309 -1176 1343
rect -1142 1309 -1136 1343
rect -1182 1271 -1136 1309
rect -1182 1237 -1176 1271
rect -1142 1237 -1136 1271
rect -1182 1218 -1136 1237
rect -1094 1343 -1048 1344
rect -1094 1309 -1088 1343
rect -1054 1309 -1048 1343
rect -1094 1271 -1048 1309
rect -1094 1237 -1088 1271
rect -1054 1237 -1048 1271
rect -1270 1165 -1264 1199
rect -1230 1165 -1224 1199
rect -1446 1093 -1440 1127
rect -1406 1093 -1400 1127
rect -5841 1026 -5821 1060
rect -5787 1026 -5749 1060
rect -5715 1026 -5677 1060
rect -5643 1026 -5605 1060
rect -5571 1026 -5533 1060
rect -5499 1026 -5461 1060
rect -5427 1026 -5408 1060
rect -5841 1008 -5408 1026
rect -2408 1060 -1976 1078
rect -2408 1026 -2390 1060
rect -2356 1026 -2318 1060
rect -2284 1026 -2246 1060
rect -2212 1026 -2174 1060
rect -2140 1026 -2102 1060
rect -2068 1026 -2030 1060
rect -1996 1026 -1976 1060
rect -2408 796 -1976 1026
rect -1446 1055 -1400 1093
rect -1446 1021 -1440 1055
rect -1406 1021 -1400 1055
rect -1446 983 -1400 1021
rect -1446 949 -1440 983
rect -1406 949 -1400 983
rect -1446 906 -1400 949
rect -1358 1127 -1312 1154
rect -1358 1093 -1352 1127
rect -1318 1093 -1312 1127
rect -1358 1055 -1312 1093
rect -1270 1127 -1224 1165
rect -1194 1212 -1130 1218
rect -1194 1160 -1188 1212
rect -1136 1160 -1130 1212
rect -1194 1154 -1130 1160
rect -1094 1199 -1048 1237
rect -1006 1343 -960 1381
rect -1006 1309 -1000 1343
rect -966 1309 -960 1343
rect -1006 1271 -960 1309
rect -1006 1237 -1000 1271
rect -966 1237 -960 1271
rect -1006 1218 -960 1237
rect -918 1559 -872 1586
rect -918 1525 -912 1559
rect -878 1525 -872 1559
rect -918 1487 -872 1525
rect -918 1453 -912 1487
rect -878 1453 -872 1487
rect -918 1415 -872 1453
rect -918 1381 -912 1415
rect -878 1381 -872 1415
rect -918 1343 -872 1381
rect -918 1309 -912 1343
rect -878 1309 -872 1343
rect -918 1271 -872 1309
rect -918 1237 -912 1271
rect -878 1237 -872 1271
rect -1094 1165 -1088 1199
rect -1054 1165 -1048 1199
rect -1270 1093 -1264 1127
rect -1230 1093 -1224 1127
rect -1270 1090 -1224 1093
rect -1182 1127 -1136 1154
rect -1182 1093 -1176 1127
rect -1142 1093 -1136 1127
rect -1358 1021 -1352 1055
rect -1318 1021 -1312 1055
rect -1279 1084 -1216 1090
rect -1279 1032 -1274 1084
rect -1222 1032 -1216 1084
rect -1279 1026 -1264 1032
rect -1358 983 -1312 1021
rect -1358 949 -1352 983
rect -1318 949 -1312 983
rect -1358 906 -1312 949
rect -1270 1021 -1264 1026
rect -1230 1026 -1216 1032
rect -1182 1055 -1136 1093
rect -1230 1021 -1224 1026
rect -1270 983 -1224 1021
rect -1270 949 -1264 983
rect -1230 949 -1224 983
rect -1270 906 -1224 949
rect -1182 1021 -1176 1055
rect -1142 1021 -1136 1055
rect -1182 983 -1136 1021
rect -1182 949 -1176 983
rect -1142 949 -1136 983
rect -1182 906 -1136 949
rect -1094 1127 -1048 1165
rect -1018 1212 -954 1218
rect -1018 1160 -1012 1212
rect -960 1160 -954 1212
rect -1018 1154 -954 1160
rect -918 1199 -872 1237
rect -830 1559 -784 1597
rect -830 1525 -824 1559
rect -790 1525 -784 1559
rect -830 1487 -784 1525
rect -830 1453 -824 1487
rect -790 1453 -784 1487
rect -830 1415 -784 1453
rect -830 1381 -824 1415
rect -790 1381 -784 1415
rect -742 2029 -736 2040
rect -702 2029 -696 2046
rect -742 1991 -696 2029
rect -742 1957 -736 1991
rect -702 1957 -696 1991
rect -742 1919 -696 1957
rect -742 1885 -736 1919
rect -702 1885 -696 1919
rect -654 2063 -608 2106
rect -654 2029 -648 2063
rect -614 2029 -608 2063
rect -654 1991 -608 2029
rect -654 1957 -648 1991
rect -614 1957 -608 1991
rect -654 1919 -608 1957
rect -654 1916 -648 1919
rect -742 1847 -696 1885
rect -666 1910 -648 1916
rect -614 1910 -608 1919
rect -666 1858 -660 1910
rect -666 1852 -608 1858
rect -742 1813 -736 1847
rect -702 1813 -696 1847
rect -742 1775 -696 1813
rect -742 1741 -736 1775
rect -702 1741 -696 1775
rect -742 1703 -696 1741
rect -742 1669 -736 1703
rect -702 1669 -696 1703
rect -742 1631 -696 1669
rect -742 1597 -736 1631
rect -702 1597 -696 1631
rect -742 1559 -696 1597
rect -742 1525 -736 1559
rect -702 1525 -696 1559
rect -742 1487 -696 1525
rect -742 1453 -736 1487
rect -702 1453 -696 1487
rect -742 1415 -696 1453
rect -742 1408 -736 1415
rect -830 1343 -784 1381
rect -754 1402 -736 1408
rect -702 1408 -696 1415
rect -654 1847 -608 1852
rect -654 1813 -648 1847
rect -614 1813 -608 1847
rect -654 1775 -608 1813
rect -654 1741 -648 1775
rect -614 1741 -608 1775
rect -654 1703 -608 1741
rect -654 1669 -648 1703
rect -614 1669 -608 1703
rect -654 1631 -608 1669
rect -566 2063 -520 2106
rect -566 2029 -560 2063
rect -526 2029 -520 2063
rect -566 1991 -520 2029
rect -566 1957 -560 1991
rect -526 1957 -520 1991
rect -566 1919 -520 1957
rect -566 1885 -560 1919
rect -526 1885 -520 1919
rect -478 2063 -432 2106
rect -390 2104 -344 2106
rect -478 2029 -472 2063
rect -438 2029 -432 2063
rect -402 2098 -344 2104
rect -402 2046 -396 2098
rect -402 2040 -384 2046
rect -478 1991 -432 2029
rect -478 1957 -472 1991
rect -438 1957 -432 1991
rect -478 1919 -432 1957
rect -478 1916 -472 1919
rect -566 1847 -520 1885
rect -490 1910 -472 1916
rect -438 1910 -432 1919
rect -490 1858 -484 1910
rect -490 1852 -432 1858
rect -566 1813 -560 1847
rect -526 1813 -520 1847
rect -566 1775 -520 1813
rect -566 1741 -560 1775
rect -526 1741 -520 1775
rect -566 1703 -520 1741
rect -566 1669 -560 1703
rect -526 1669 -520 1703
rect -566 1650 -520 1669
rect -478 1847 -432 1852
rect -478 1813 -472 1847
rect -438 1813 -432 1847
rect -478 1775 -432 1813
rect -478 1741 -472 1775
rect -438 1741 -432 1775
rect -478 1703 -432 1741
rect -478 1669 -472 1703
rect -438 1669 -432 1703
rect -654 1597 -648 1631
rect -614 1597 -608 1631
rect -654 1559 -608 1597
rect -574 1644 -510 1650
rect -574 1592 -568 1644
rect -516 1592 -510 1644
rect -574 1586 -510 1592
rect -478 1631 -432 1669
rect -478 1597 -472 1631
rect -438 1597 -432 1631
rect -654 1525 -648 1559
rect -614 1525 -608 1559
rect -654 1487 -608 1525
rect -654 1453 -648 1487
rect -614 1453 -608 1487
rect -654 1415 -608 1453
rect -702 1402 -690 1408
rect -754 1350 -748 1402
rect -696 1350 -690 1402
rect -754 1344 -690 1350
rect -654 1381 -648 1415
rect -614 1381 -608 1415
rect -830 1309 -824 1343
rect -790 1309 -784 1343
rect -830 1271 -784 1309
rect -830 1237 -824 1271
rect -790 1237 -784 1271
rect -830 1218 -784 1237
rect -742 1343 -696 1344
rect -742 1309 -736 1343
rect -702 1309 -696 1343
rect -742 1271 -696 1309
rect -742 1237 -736 1271
rect -702 1237 -696 1271
rect -918 1165 -912 1199
rect -878 1165 -872 1199
rect -1094 1093 -1088 1127
rect -1054 1093 -1048 1127
rect -1094 1055 -1048 1093
rect -1094 1021 -1088 1055
rect -1054 1021 -1048 1055
rect -1094 983 -1048 1021
rect -1094 949 -1088 983
rect -1054 949 -1048 983
rect -1094 906 -1048 949
rect -1006 1127 -960 1154
rect -1006 1093 -1000 1127
rect -966 1093 -960 1127
rect -1006 1055 -960 1093
rect -918 1127 -872 1165
rect -842 1212 -778 1218
rect -842 1160 -836 1212
rect -784 1160 -778 1212
rect -842 1154 -778 1160
rect -742 1199 -696 1237
rect -654 1343 -608 1381
rect -654 1309 -648 1343
rect -614 1309 -608 1343
rect -654 1271 -608 1309
rect -654 1237 -648 1271
rect -614 1237 -608 1271
rect -654 1218 -608 1237
rect -566 1559 -520 1586
rect -566 1525 -560 1559
rect -526 1525 -520 1559
rect -566 1487 -520 1525
rect -566 1453 -560 1487
rect -526 1453 -520 1487
rect -566 1415 -520 1453
rect -566 1381 -560 1415
rect -526 1381 -520 1415
rect -566 1343 -520 1381
rect -566 1309 -560 1343
rect -526 1309 -520 1343
rect -566 1271 -520 1309
rect -566 1237 -560 1271
rect -526 1237 -520 1271
rect -742 1165 -736 1199
rect -702 1165 -696 1199
rect -918 1093 -912 1127
rect -878 1093 -872 1127
rect -918 1090 -872 1093
rect -830 1127 -784 1154
rect -830 1093 -824 1127
rect -790 1093 -784 1127
rect -1006 1021 -1000 1055
rect -966 1021 -960 1055
rect -927 1084 -863 1090
rect -927 1032 -922 1084
rect -870 1032 -863 1084
rect -927 1026 -912 1032
rect -1006 983 -960 1021
rect -1006 949 -1000 983
rect -966 949 -960 983
rect -1006 906 -960 949
rect -918 1021 -912 1026
rect -878 1026 -863 1032
rect -830 1055 -784 1093
rect -878 1021 -872 1026
rect -918 983 -872 1021
rect -918 949 -912 983
rect -878 949 -872 983
rect -918 906 -872 949
rect -830 1021 -824 1055
rect -790 1021 -784 1055
rect -830 983 -784 1021
rect -830 949 -824 983
rect -790 949 -784 983
rect -830 906 -784 949
rect -742 1127 -696 1165
rect -666 1212 -602 1218
rect -666 1160 -660 1212
rect -608 1160 -602 1212
rect -666 1154 -602 1160
rect -566 1199 -520 1237
rect -478 1559 -432 1597
rect -478 1525 -472 1559
rect -438 1525 -432 1559
rect -478 1487 -432 1525
rect -478 1453 -472 1487
rect -438 1453 -432 1487
rect -478 1415 -432 1453
rect -478 1381 -472 1415
rect -438 1381 -432 1415
rect -390 2029 -384 2040
rect -350 2029 -344 2046
rect -390 1991 -344 2029
rect -390 1957 -384 1991
rect -350 1957 -344 1991
rect -390 1919 -344 1957
rect -390 1885 -384 1919
rect -350 1885 -344 1919
rect -302 2063 -256 2106
rect -302 2029 -296 2063
rect -262 2029 -256 2063
rect -302 1991 -256 2029
rect -302 1957 -296 1991
rect -262 1957 -256 1991
rect -302 1919 -256 1957
rect -302 1916 -296 1919
rect -390 1847 -344 1885
rect -314 1910 -296 1916
rect -262 1910 -256 1919
rect -314 1858 -308 1910
rect -314 1852 -256 1858
rect -390 1813 -384 1847
rect -350 1813 -344 1847
rect -390 1775 -344 1813
rect -390 1741 -384 1775
rect -350 1741 -344 1775
rect -390 1703 -344 1741
rect -390 1669 -384 1703
rect -350 1669 -344 1703
rect -390 1631 -344 1669
rect -390 1597 -384 1631
rect -350 1597 -344 1631
rect -390 1559 -344 1597
rect -390 1525 -384 1559
rect -350 1525 -344 1559
rect -390 1487 -344 1525
rect -390 1453 -384 1487
rect -350 1453 -344 1487
rect -390 1415 -344 1453
rect -390 1408 -384 1415
rect -478 1343 -432 1381
rect -402 1402 -384 1408
rect -350 1408 -344 1415
rect -302 1847 -256 1852
rect -302 1813 -296 1847
rect -262 1813 -256 1847
rect -302 1775 -256 1813
rect -302 1741 -296 1775
rect -262 1741 -256 1775
rect -302 1703 -256 1741
rect -302 1669 -296 1703
rect -262 1669 -256 1703
rect -302 1631 -256 1669
rect -214 2063 -168 2106
rect -214 2029 -208 2063
rect -174 2029 -168 2063
rect -214 1991 -168 2029
rect -214 1957 -208 1991
rect -174 1957 -168 1991
rect -214 1919 -168 1957
rect -214 1885 -208 1919
rect -174 1885 -168 1919
rect -126 2063 -80 2106
rect -38 2104 8 2106
rect -126 2029 -120 2063
rect -86 2029 -80 2063
rect -50 2098 8 2104
rect -50 2046 -44 2098
rect -50 2040 -32 2046
rect -126 1991 -80 2029
rect -126 1957 -120 1991
rect -86 1957 -80 1991
rect -126 1919 -80 1957
rect -126 1916 -120 1919
rect -214 1847 -168 1885
rect -138 1910 -120 1916
rect -86 1910 -80 1919
rect -138 1858 -132 1910
rect -138 1852 -80 1858
rect -214 1813 -208 1847
rect -174 1813 -168 1847
rect -214 1775 -168 1813
rect -214 1741 -208 1775
rect -174 1741 -168 1775
rect -214 1703 -168 1741
rect -214 1669 -208 1703
rect -174 1669 -168 1703
rect -214 1650 -168 1669
rect -126 1847 -80 1852
rect -126 1813 -120 1847
rect -86 1813 -80 1847
rect -126 1775 -80 1813
rect -126 1741 -120 1775
rect -86 1741 -80 1775
rect -126 1703 -80 1741
rect -126 1669 -120 1703
rect -86 1669 -80 1703
rect -302 1597 -296 1631
rect -262 1597 -256 1631
rect -302 1559 -256 1597
rect -222 1644 -158 1650
rect -222 1592 -216 1644
rect -164 1592 -158 1644
rect -222 1586 -158 1592
rect -126 1631 -80 1669
rect -126 1597 -120 1631
rect -86 1597 -80 1631
rect -302 1525 -296 1559
rect -262 1525 -256 1559
rect -302 1487 -256 1525
rect -302 1453 -296 1487
rect -262 1453 -256 1487
rect -302 1415 -256 1453
rect -350 1402 -338 1408
rect -402 1350 -396 1402
rect -344 1350 -338 1402
rect -402 1344 -338 1350
rect -302 1381 -296 1415
rect -262 1381 -256 1415
rect -478 1309 -472 1343
rect -438 1309 -432 1343
rect -478 1271 -432 1309
rect -478 1237 -472 1271
rect -438 1237 -432 1271
rect -478 1218 -432 1237
rect -390 1343 -344 1344
rect -390 1309 -384 1343
rect -350 1309 -344 1343
rect -390 1271 -344 1309
rect -390 1237 -384 1271
rect -350 1237 -344 1271
rect -566 1165 -560 1199
rect -526 1165 -520 1199
rect -742 1093 -736 1127
rect -702 1093 -696 1127
rect -742 1055 -696 1093
rect -742 1021 -736 1055
rect -702 1021 -696 1055
rect -742 983 -696 1021
rect -742 949 -736 983
rect -702 949 -696 983
rect -742 906 -696 949
rect -654 1127 -608 1154
rect -654 1093 -648 1127
rect -614 1093 -608 1127
rect -654 1055 -608 1093
rect -566 1127 -520 1165
rect -490 1212 -426 1218
rect -490 1160 -484 1212
rect -432 1160 -426 1212
rect -490 1154 -426 1160
rect -390 1199 -344 1237
rect -302 1343 -256 1381
rect -302 1309 -296 1343
rect -262 1309 -256 1343
rect -302 1271 -256 1309
rect -302 1237 -296 1271
rect -262 1237 -256 1271
rect -302 1218 -256 1237
rect -214 1559 -168 1586
rect -214 1525 -208 1559
rect -174 1525 -168 1559
rect -214 1487 -168 1525
rect -214 1453 -208 1487
rect -174 1453 -168 1487
rect -214 1415 -168 1453
rect -214 1381 -208 1415
rect -174 1381 -168 1415
rect -214 1343 -168 1381
rect -214 1309 -208 1343
rect -174 1309 -168 1343
rect -214 1271 -168 1309
rect -214 1237 -208 1271
rect -174 1237 -168 1271
rect -390 1165 -384 1199
rect -350 1165 -344 1199
rect -566 1093 -560 1127
rect -526 1093 -520 1127
rect -566 1090 -520 1093
rect -478 1127 -432 1154
rect -478 1093 -472 1127
rect -438 1093 -432 1127
rect -654 1021 -648 1055
rect -614 1021 -608 1055
rect -575 1084 -511 1090
rect -575 1032 -570 1084
rect -518 1032 -511 1084
rect -575 1026 -560 1032
rect -654 983 -608 1021
rect -654 949 -648 983
rect -614 949 -608 983
rect -654 906 -608 949
rect -566 1021 -560 1026
rect -526 1026 -511 1032
rect -478 1055 -432 1093
rect -526 1021 -520 1026
rect -566 983 -520 1021
rect -566 949 -560 983
rect -526 949 -520 983
rect -566 906 -520 949
rect -478 1021 -472 1055
rect -438 1021 -432 1055
rect -478 983 -432 1021
rect -478 949 -472 983
rect -438 949 -432 983
rect -478 906 -432 949
rect -390 1127 -344 1165
rect -314 1212 -250 1218
rect -314 1160 -308 1212
rect -256 1160 -250 1212
rect -314 1154 -250 1160
rect -214 1199 -168 1237
rect -126 1559 -80 1597
rect -126 1525 -120 1559
rect -86 1525 -80 1559
rect -126 1487 -80 1525
rect -126 1453 -120 1487
rect -86 1453 -80 1487
rect -126 1415 -80 1453
rect -126 1381 -120 1415
rect -86 1381 -80 1415
rect -38 2029 -32 2040
rect 2 2029 8 2046
rect -38 1991 8 2029
rect -38 1957 -32 1991
rect 2 1957 8 1991
rect -38 1919 8 1957
rect -38 1885 -32 1919
rect 2 1885 8 1919
rect 50 2063 96 2106
rect 50 2029 56 2063
rect 90 2029 96 2063
rect 50 1991 96 2029
rect 50 1957 56 1991
rect 90 1957 96 1991
rect 50 1919 96 1957
rect 50 1916 56 1919
rect -38 1847 8 1885
rect 38 1910 56 1916
rect 90 1910 96 1919
rect 38 1858 44 1910
rect 38 1852 96 1858
rect -38 1813 -32 1847
rect 2 1813 8 1847
rect -38 1775 8 1813
rect -38 1741 -32 1775
rect 2 1741 8 1775
rect -38 1703 8 1741
rect -38 1669 -32 1703
rect 2 1669 8 1703
rect -38 1631 8 1669
rect -38 1597 -32 1631
rect 2 1597 8 1631
rect -38 1559 8 1597
rect -38 1525 -32 1559
rect 2 1525 8 1559
rect -38 1487 8 1525
rect -38 1453 -32 1487
rect 2 1453 8 1487
rect -38 1415 8 1453
rect -38 1408 -32 1415
rect -126 1343 -80 1381
rect -50 1402 -32 1408
rect 2 1408 8 1415
rect 50 1847 96 1852
rect 50 1813 56 1847
rect 90 1813 96 1847
rect 50 1775 96 1813
rect 50 1741 56 1775
rect 90 1741 96 1775
rect 50 1703 96 1741
rect 50 1669 56 1703
rect 90 1669 96 1703
rect 50 1631 96 1669
rect 138 2063 184 2106
rect 138 2029 144 2063
rect 178 2029 184 2063
rect 138 1991 184 2029
rect 138 1957 144 1991
rect 178 1957 184 1991
rect 138 1919 184 1957
rect 138 1885 144 1919
rect 178 1885 184 1919
rect 226 2063 272 2106
rect 314 2104 360 2106
rect 226 2029 232 2063
rect 266 2029 272 2063
rect 302 2098 366 2104
rect 302 2046 308 2098
rect 360 2046 366 2098
rect 302 2040 320 2046
rect 226 1991 272 2029
rect 226 1957 232 1991
rect 266 1957 272 1991
rect 226 1919 272 1957
rect 226 1916 232 1919
rect 138 1847 184 1885
rect 214 1910 232 1916
rect 266 1910 272 1919
rect 214 1858 220 1910
rect 214 1852 272 1858
rect 138 1813 144 1847
rect 178 1813 184 1847
rect 138 1775 184 1813
rect 138 1741 144 1775
rect 178 1741 184 1775
rect 138 1703 184 1741
rect 138 1669 144 1703
rect 178 1669 184 1703
rect 138 1650 184 1669
rect 226 1847 272 1852
rect 226 1813 232 1847
rect 266 1813 272 1847
rect 226 1775 272 1813
rect 226 1741 232 1775
rect 266 1741 272 1775
rect 226 1703 272 1741
rect 226 1669 232 1703
rect 266 1669 272 1703
rect 50 1597 56 1631
rect 90 1597 96 1631
rect 50 1559 96 1597
rect 130 1644 194 1650
rect 130 1592 136 1644
rect 188 1592 194 1644
rect 130 1586 194 1592
rect 226 1631 272 1669
rect 226 1597 232 1631
rect 266 1597 272 1631
rect 50 1525 56 1559
rect 90 1525 96 1559
rect 50 1487 96 1525
rect 50 1453 56 1487
rect 90 1453 96 1487
rect 50 1415 96 1453
rect 2 1402 14 1408
rect -50 1350 -44 1402
rect 8 1350 14 1402
rect -50 1344 14 1350
rect 50 1381 56 1415
rect 90 1381 96 1415
rect -126 1309 -120 1343
rect -86 1309 -80 1343
rect -126 1271 -80 1309
rect -126 1237 -120 1271
rect -86 1237 -80 1271
rect -126 1218 -80 1237
rect -38 1343 8 1344
rect -38 1309 -32 1343
rect 2 1309 8 1343
rect -38 1271 8 1309
rect -38 1237 -32 1271
rect 2 1237 8 1271
rect -214 1165 -208 1199
rect -174 1165 -168 1199
rect -390 1093 -384 1127
rect -350 1093 -344 1127
rect -390 1055 -344 1093
rect -390 1021 -384 1055
rect -350 1021 -344 1055
rect -390 983 -344 1021
rect -390 949 -384 983
rect -350 949 -344 983
rect -390 906 -344 949
rect -302 1127 -256 1154
rect -302 1093 -296 1127
rect -262 1093 -256 1127
rect -302 1055 -256 1093
rect -214 1127 -168 1165
rect -138 1212 -74 1218
rect -138 1160 -132 1212
rect -80 1160 -74 1212
rect -138 1154 -74 1160
rect -38 1199 8 1237
rect 50 1343 96 1381
rect 50 1309 56 1343
rect 90 1309 96 1343
rect 50 1271 96 1309
rect 50 1237 56 1271
rect 90 1237 96 1271
rect 50 1218 96 1237
rect 138 1559 184 1586
rect 138 1525 144 1559
rect 178 1525 184 1559
rect 138 1487 184 1525
rect 138 1453 144 1487
rect 178 1453 184 1487
rect 138 1415 184 1453
rect 138 1381 144 1415
rect 178 1381 184 1415
rect 138 1343 184 1381
rect 138 1309 144 1343
rect 178 1309 184 1343
rect 138 1271 184 1309
rect 138 1237 144 1271
rect 178 1237 184 1271
rect -38 1165 -32 1199
rect 2 1165 8 1199
rect -214 1093 -208 1127
rect -174 1093 -168 1127
rect -214 1090 -168 1093
rect -126 1127 -80 1154
rect -126 1093 -120 1127
rect -86 1093 -80 1127
rect -302 1021 -296 1055
rect -262 1021 -256 1055
rect -223 1084 -159 1090
rect -223 1032 -218 1084
rect -166 1032 -159 1084
rect -223 1026 -208 1032
rect -302 983 -256 1021
rect -302 949 -296 983
rect -262 949 -256 983
rect -302 906 -256 949
rect -214 1021 -208 1026
rect -174 1026 -159 1032
rect -126 1055 -80 1093
rect -174 1021 -168 1026
rect -214 983 -168 1021
rect -214 949 -208 983
rect -174 949 -168 983
rect -214 906 -168 949
rect -126 1021 -120 1055
rect -86 1021 -80 1055
rect -126 983 -80 1021
rect -126 949 -120 983
rect -86 949 -80 983
rect -126 906 -80 949
rect -38 1127 8 1165
rect 38 1212 102 1218
rect 38 1160 44 1212
rect 96 1160 102 1212
rect 38 1154 102 1160
rect 138 1199 184 1237
rect 226 1559 272 1597
rect 226 1525 232 1559
rect 266 1525 272 1559
rect 226 1487 272 1525
rect 226 1453 232 1487
rect 266 1453 272 1487
rect 226 1415 272 1453
rect 226 1381 232 1415
rect 266 1381 272 1415
rect 314 2029 320 2040
rect 354 2040 366 2046
rect 724 2098 788 2104
rect 1084 2098 1140 2104
rect 724 2046 730 2098
rect 782 2046 788 2098
rect 1134 2046 1140 2098
rect 724 2040 788 2046
rect 1084 2040 1140 2046
rect 1434 2098 1492 2104
rect 1486 2046 1492 2098
rect 1434 2040 1492 2046
rect 1786 2098 1844 2104
rect 1838 2046 1844 2098
rect 1786 2040 1844 2046
rect 2138 2098 2196 2104
rect 2190 2046 2196 2098
rect 2138 2040 2196 2046
rect 2490 2098 2608 2104
rect 2542 2046 2608 2098
rect 3209 2089 3635 2189
rect 2490 2040 2608 2046
rect 354 2029 360 2040
rect 314 1991 360 2029
rect 314 1957 320 1991
rect 354 1957 360 1991
rect 314 1919 360 1957
rect 314 1885 320 1919
rect 354 1885 360 1919
rect 314 1847 360 1885
rect 818 1910 876 1916
rect 870 1858 876 1910
rect 818 1852 876 1858
rect 994 1910 1052 1916
rect 1046 1858 1052 1910
rect 994 1852 1052 1858
rect 1170 1910 1228 1916
rect 1222 1858 1228 1910
rect 1170 1852 1228 1858
rect 1346 1910 1404 1916
rect 1398 1858 1404 1910
rect 1346 1852 1404 1858
rect 1522 1910 1580 1916
rect 1574 1858 1580 1910
rect 1522 1852 1580 1858
rect 1698 1910 1756 1916
rect 1750 1858 1756 1910
rect 1698 1852 1756 1858
rect 1874 1910 1932 1916
rect 2086 1910 2108 1916
rect 1926 1858 1932 1910
rect 2102 1858 2108 1910
rect 1874 1852 1932 1858
rect 2086 1852 2108 1858
rect 2220 1910 2278 1916
rect 2220 1858 2226 1910
rect 2220 1852 2278 1858
rect 2396 1910 2454 1916
rect 2396 1858 2402 1910
rect 2396 1852 2454 1858
rect 3182 1889 3647 1911
rect 314 1813 320 1847
rect 354 1813 360 1847
rect 314 1775 360 1813
rect 314 1741 320 1775
rect 354 1741 360 1775
rect 314 1703 360 1741
rect 314 1669 320 1703
rect 354 1669 360 1703
rect 314 1631 360 1669
rect 3182 1837 3240 1889
rect 3292 1837 3304 1889
rect 3356 1837 3368 1889
rect 3420 1837 3432 1889
rect 3484 1837 3496 1889
rect 3548 1837 3647 1889
rect 3182 1650 3647 1837
rect 6651 1886 7104 2159
rect 6651 1834 6716 1886
rect 6768 1834 6780 1886
rect 6832 1834 6844 1886
rect 6896 1834 6908 1886
rect 6960 1834 6972 1886
rect 7024 1834 7104 1886
rect 6651 1815 7104 1834
rect 314 1597 320 1631
rect 354 1597 360 1631
rect 314 1559 360 1597
rect 896 1644 960 1650
rect 896 1592 902 1644
rect 954 1592 960 1644
rect 896 1586 960 1592
rect 1248 1644 1312 1650
rect 1248 1592 1254 1644
rect 1306 1592 1312 1644
rect 1248 1586 1312 1592
rect 1600 1644 1664 1650
rect 1600 1592 1606 1644
rect 1658 1592 1664 1644
rect 1600 1586 1664 1592
rect 1952 1644 2016 1650
rect 1952 1592 1958 1644
rect 2010 1592 2016 1644
rect 1952 1586 2016 1592
rect 2304 1644 2368 1650
rect 2304 1592 2310 1644
rect 2362 1592 2368 1644
rect 2304 1586 2368 1592
rect 314 1525 320 1559
rect 354 1525 360 1559
rect 314 1487 360 1525
rect 314 1453 320 1487
rect 354 1453 360 1487
rect 314 1415 360 1453
rect 314 1408 320 1415
rect 226 1343 272 1381
rect 302 1402 320 1408
rect 354 1408 360 1415
rect 3181 1558 3647 1650
rect 354 1402 366 1408
rect 302 1350 308 1402
rect 360 1350 366 1402
rect 302 1344 366 1350
rect 724 1402 788 1408
rect 724 1350 730 1402
rect 782 1350 788 1402
rect 724 1344 788 1350
rect 1076 1402 1140 1408
rect 1076 1350 1082 1402
rect 1134 1350 1140 1402
rect 1076 1344 1140 1350
rect 1428 1402 1492 1408
rect 1428 1350 1434 1402
rect 1486 1350 1492 1402
rect 1428 1344 1492 1350
rect 1780 1402 1844 1408
rect 1780 1350 1786 1402
rect 1838 1350 1844 1402
rect 1780 1344 1844 1350
rect 2132 1402 2196 1408
rect 2132 1350 2138 1402
rect 2190 1350 2196 1402
rect 2132 1344 2196 1350
rect 2484 1402 2548 1408
rect 2484 1350 2490 1402
rect 2542 1350 2548 1402
rect 2484 1344 2548 1350
rect 226 1309 232 1343
rect 266 1309 272 1343
rect 226 1271 272 1309
rect 226 1237 232 1271
rect 266 1237 272 1271
rect 226 1218 272 1237
rect 314 1343 360 1344
rect 314 1309 320 1343
rect 354 1309 360 1343
rect 314 1271 360 1309
rect 314 1237 320 1271
rect 354 1237 360 1271
rect 3181 1339 3646 1558
rect 6652 1539 7419 1720
rect 3181 1287 3241 1339
rect 3293 1287 3305 1339
rect 3357 1287 3369 1339
rect 3421 1287 3433 1339
rect 3485 1287 3497 1339
rect 3549 1287 3646 1339
rect 3181 1265 3646 1287
rect 6685 1335 7118 1361
rect 6685 1283 6750 1335
rect 6802 1283 6814 1335
rect 6866 1283 6878 1335
rect 6930 1283 6942 1335
rect 6994 1283 7006 1335
rect 7058 1283 7118 1335
rect 138 1165 144 1199
rect 178 1165 184 1199
rect -38 1093 -32 1127
rect 2 1093 8 1127
rect -38 1055 8 1093
rect -38 1021 -32 1055
rect 2 1021 8 1055
rect -38 983 8 1021
rect -38 949 -32 983
rect 2 949 8 983
rect -38 906 8 949
rect 50 1127 96 1154
rect 50 1093 56 1127
rect 90 1093 96 1127
rect 50 1055 96 1093
rect 138 1127 184 1165
rect 214 1212 278 1218
rect 214 1160 220 1212
rect 272 1160 278 1212
rect 214 1154 278 1160
rect 314 1199 360 1237
rect 314 1165 320 1199
rect 354 1165 360 1199
rect 138 1093 144 1127
rect 178 1093 184 1127
rect 138 1090 184 1093
rect 226 1127 272 1154
rect 226 1093 232 1127
rect 266 1093 272 1127
rect 50 1021 56 1055
rect 90 1021 96 1055
rect 129 1084 193 1090
rect 129 1032 134 1084
rect 186 1032 193 1084
rect 129 1026 144 1032
rect 50 983 96 1021
rect 50 949 56 983
rect 90 949 96 983
rect 50 906 96 949
rect 138 1021 144 1026
rect 178 1026 193 1032
rect 226 1055 272 1093
rect 178 1021 184 1026
rect 138 983 184 1021
rect 138 949 144 983
rect 178 949 184 983
rect 138 906 184 949
rect 226 1021 232 1055
rect 266 1021 272 1055
rect 226 983 272 1021
rect 226 949 232 983
rect 266 949 272 983
rect 226 906 272 949
rect 314 1127 360 1165
rect 812 1212 876 1218
rect 812 1160 818 1212
rect 870 1160 876 1212
rect 812 1154 876 1160
rect 988 1212 1052 1218
rect 988 1160 994 1212
rect 1046 1160 1052 1212
rect 988 1154 1052 1160
rect 1164 1212 1228 1218
rect 1164 1160 1170 1212
rect 1222 1160 1228 1212
rect 1164 1154 1228 1160
rect 1340 1212 1404 1218
rect 1340 1160 1346 1212
rect 1398 1160 1404 1212
rect 1340 1154 1404 1160
rect 1516 1212 1580 1218
rect 1516 1160 1522 1212
rect 1574 1160 1580 1212
rect 1516 1154 1580 1160
rect 1692 1212 1756 1218
rect 1692 1160 1698 1212
rect 1750 1160 1756 1212
rect 1692 1154 1756 1160
rect 1868 1212 1932 1218
rect 1868 1160 1874 1212
rect 1926 1160 1932 1212
rect 1868 1154 1932 1160
rect 2044 1212 2108 1218
rect 2044 1160 2050 1212
rect 2102 1160 2108 1212
rect 2044 1154 2108 1160
rect 2220 1212 2284 1218
rect 2220 1160 2226 1212
rect 2278 1160 2284 1212
rect 2220 1154 2284 1160
rect 2396 1212 2460 1218
rect 2396 1160 2402 1212
rect 2454 1160 2460 1212
rect 2396 1154 2460 1160
rect 314 1093 320 1127
rect 354 1093 360 1127
rect 314 1055 360 1093
rect 314 1021 320 1055
rect 354 1021 360 1055
rect 897 1084 961 1090
rect 897 1032 904 1084
rect 956 1032 961 1084
rect 897 1026 961 1032
rect 1249 1084 1313 1090
rect 1249 1032 1256 1084
rect 1308 1032 1313 1084
rect 1249 1026 1313 1032
rect 1601 1084 1665 1090
rect 1601 1032 1608 1084
rect 1660 1032 1665 1084
rect 1601 1026 1665 1032
rect 1953 1084 2017 1090
rect 1953 1032 1960 1084
rect 2012 1032 2017 1084
rect 1953 1026 2017 1032
rect 2306 1084 2369 1090
rect 2306 1032 2312 1084
rect 2364 1032 2369 1084
rect 2306 1026 2369 1032
rect 314 983 360 1021
rect 314 949 320 983
rect 354 949 360 983
rect 314 906 360 949
rect 3249 796 3685 1113
rect 6685 1041 7118 1283
rect -2408 778 220 796
rect -2408 744 -1273 778
rect -1239 744 -1201 778
rect -1167 744 -1129 778
rect -1095 744 -1057 778
rect -1023 744 -985 778
rect -951 744 -913 778
rect -879 744 -841 778
rect -807 744 -769 778
rect -735 744 -697 778
rect -663 744 -625 778
rect -591 744 -553 778
rect -519 744 -481 778
rect -447 744 -409 778
rect -375 744 -337 778
rect -303 744 -265 778
rect -231 744 -193 778
rect -159 744 -121 778
rect -87 744 -49 778
rect -15 744 23 778
rect 57 744 95 778
rect 129 744 167 778
rect 201 744 220 778
rect -2408 726 220 744
rect 870 778 3685 796
rect 870 744 889 778
rect 923 744 961 778
rect 995 744 1033 778
rect 1067 744 1105 778
rect 1139 744 1177 778
rect 1211 744 1249 778
rect 1283 744 1321 778
rect 1355 744 1393 778
rect 1427 744 1465 778
rect 1499 744 1537 778
rect 1571 744 1609 778
rect 1643 744 1681 778
rect 1715 744 1753 778
rect 1787 744 1825 778
rect 1859 744 1897 778
rect 1931 744 1969 778
rect 2003 744 2041 778
rect 2075 744 2113 778
rect 2147 744 2185 778
rect 2219 744 2257 778
rect 2291 744 2329 778
rect 2363 744 3685 778
rect 870 726 3685 744
<< via1 >>
rect -1452 2063 -1400 2098
rect -1452 2046 -1440 2063
rect -1440 2046 -1406 2063
rect -1406 2046 -1400 2063
rect -5747 1801 -5695 1853
rect -5683 1801 -5631 1853
rect -5619 1801 -5567 1853
rect -5555 1801 -5503 1853
rect -5491 1801 -5439 1853
rect -2271 1804 -2219 1856
rect -2207 1804 -2155 1856
rect -2143 1804 -2091 1856
rect -2079 1804 -2027 1856
rect -2015 1804 -1963 1856
rect -1364 1885 -1352 1910
rect -1352 1885 -1318 1910
rect -1318 1885 -1312 1910
rect -1364 1858 -1312 1885
rect -1100 2063 -1048 2098
rect -1100 2046 -1088 2063
rect -1088 2046 -1054 2063
rect -1054 2046 -1048 2063
rect -5781 1250 -5729 1302
rect -5717 1250 -5665 1302
rect -5653 1250 -5601 1302
rect -5589 1250 -5537 1302
rect -5525 1250 -5473 1302
rect -1188 1885 -1176 1910
rect -1176 1885 -1142 1910
rect -1142 1885 -1136 1910
rect -1188 1858 -1136 1885
rect -1272 1631 -1220 1644
rect -1272 1597 -1264 1631
rect -1264 1597 -1230 1631
rect -1230 1597 -1220 1631
rect -1272 1592 -1220 1597
rect -1452 1381 -1440 1402
rect -1440 1381 -1406 1402
rect -1406 1381 -1400 1402
rect -1452 1350 -1400 1381
rect -2272 1254 -2220 1306
rect -2208 1254 -2156 1306
rect -2144 1254 -2092 1306
rect -2080 1254 -2028 1306
rect -2016 1254 -1964 1306
rect -1364 1199 -1312 1212
rect -1364 1165 -1352 1199
rect -1352 1165 -1318 1199
rect -1318 1165 -1312 1199
rect -1364 1160 -1312 1165
rect -1012 1885 -1000 1910
rect -1000 1885 -966 1910
rect -966 1885 -960 1910
rect -1012 1858 -960 1885
rect -748 2063 -696 2098
rect -748 2046 -736 2063
rect -736 2046 -702 2063
rect -702 2046 -696 2063
rect -836 1885 -824 1910
rect -824 1885 -790 1910
rect -790 1885 -784 1910
rect -836 1858 -784 1885
rect -920 1631 -868 1644
rect -920 1597 -912 1631
rect -912 1597 -878 1631
rect -878 1597 -868 1631
rect -920 1592 -868 1597
rect -1100 1381 -1088 1402
rect -1088 1381 -1054 1402
rect -1054 1381 -1048 1402
rect -1100 1350 -1048 1381
rect -1188 1199 -1136 1212
rect -1188 1165 -1176 1199
rect -1176 1165 -1142 1199
rect -1142 1165 -1136 1199
rect -1188 1160 -1136 1165
rect -1274 1055 -1222 1084
rect -1274 1032 -1264 1055
rect -1264 1032 -1230 1055
rect -1230 1032 -1222 1055
rect -1012 1199 -960 1212
rect -1012 1165 -1000 1199
rect -1000 1165 -966 1199
rect -966 1165 -960 1199
rect -1012 1160 -960 1165
rect -660 1885 -648 1910
rect -648 1885 -614 1910
rect -614 1885 -608 1910
rect -660 1858 -608 1885
rect -396 2063 -344 2098
rect -396 2046 -384 2063
rect -384 2046 -350 2063
rect -350 2046 -344 2063
rect -484 1885 -472 1910
rect -472 1885 -438 1910
rect -438 1885 -432 1910
rect -484 1858 -432 1885
rect -568 1631 -516 1644
rect -568 1597 -560 1631
rect -560 1597 -526 1631
rect -526 1597 -516 1631
rect -568 1592 -516 1597
rect -748 1381 -736 1402
rect -736 1381 -702 1402
rect -702 1381 -696 1402
rect -748 1350 -696 1381
rect -836 1199 -784 1212
rect -836 1165 -824 1199
rect -824 1165 -790 1199
rect -790 1165 -784 1199
rect -836 1160 -784 1165
rect -922 1055 -870 1084
rect -922 1032 -912 1055
rect -912 1032 -878 1055
rect -878 1032 -870 1055
rect -660 1199 -608 1212
rect -660 1165 -648 1199
rect -648 1165 -614 1199
rect -614 1165 -608 1199
rect -660 1160 -608 1165
rect -308 1885 -296 1910
rect -296 1885 -262 1910
rect -262 1885 -256 1910
rect -308 1858 -256 1885
rect -44 2063 8 2098
rect -44 2046 -32 2063
rect -32 2046 2 2063
rect 2 2046 8 2063
rect -132 1885 -120 1910
rect -120 1885 -86 1910
rect -86 1885 -80 1910
rect -132 1858 -80 1885
rect -216 1631 -164 1644
rect -216 1597 -208 1631
rect -208 1597 -174 1631
rect -174 1597 -164 1631
rect -216 1592 -164 1597
rect -396 1381 -384 1402
rect -384 1381 -350 1402
rect -350 1381 -344 1402
rect -396 1350 -344 1381
rect -484 1199 -432 1212
rect -484 1165 -472 1199
rect -472 1165 -438 1199
rect -438 1165 -432 1199
rect -484 1160 -432 1165
rect -570 1055 -518 1084
rect -570 1032 -560 1055
rect -560 1032 -526 1055
rect -526 1032 -518 1055
rect -308 1199 -256 1212
rect -308 1165 -296 1199
rect -296 1165 -262 1199
rect -262 1165 -256 1199
rect -308 1160 -256 1165
rect 44 1885 56 1910
rect 56 1885 90 1910
rect 90 1885 96 1910
rect 44 1858 96 1885
rect 308 2063 360 2098
rect 308 2046 320 2063
rect 320 2046 354 2063
rect 354 2046 360 2063
rect 220 1885 232 1910
rect 232 1885 266 1910
rect 266 1885 272 1910
rect 220 1858 272 1885
rect 136 1631 188 1644
rect 136 1597 144 1631
rect 144 1597 178 1631
rect 178 1597 188 1631
rect 136 1592 188 1597
rect -44 1381 -32 1402
rect -32 1381 2 1402
rect 2 1381 8 1402
rect -44 1350 8 1381
rect -132 1199 -80 1212
rect -132 1165 -120 1199
rect -120 1165 -86 1199
rect -86 1165 -80 1199
rect -132 1160 -80 1165
rect -218 1055 -166 1084
rect -218 1032 -208 1055
rect -208 1032 -174 1055
rect -174 1032 -166 1055
rect 44 1199 96 1212
rect 44 1165 56 1199
rect 56 1165 90 1199
rect 90 1165 96 1199
rect 44 1160 96 1165
rect 730 2046 782 2098
rect 1082 2046 1134 2098
rect 1434 2046 1486 2098
rect 1786 2046 1838 2098
rect 2138 2046 2190 2098
rect 2490 2046 2542 2098
rect 818 1858 870 1910
rect 994 1858 1046 1910
rect 1170 1858 1222 1910
rect 1346 1858 1398 1910
rect 1522 1858 1574 1910
rect 1698 1858 1750 1910
rect 1874 1858 1926 1910
rect 2050 1858 2102 1910
rect 2226 1858 2278 1910
rect 2402 1858 2454 1910
rect 3240 1837 3292 1889
rect 3304 1837 3356 1889
rect 3368 1837 3420 1889
rect 3432 1837 3484 1889
rect 3496 1837 3548 1889
rect 6716 1834 6768 1886
rect 6780 1834 6832 1886
rect 6844 1834 6896 1886
rect 6908 1834 6960 1886
rect 6972 1834 7024 1886
rect 902 1592 954 1644
rect 1254 1592 1306 1644
rect 1606 1592 1658 1644
rect 1958 1592 2010 1644
rect 2310 1592 2362 1644
rect 308 1381 320 1402
rect 320 1381 354 1402
rect 354 1381 360 1402
rect 308 1350 360 1381
rect 730 1350 782 1402
rect 1082 1350 1134 1402
rect 1434 1350 1486 1402
rect 1786 1350 1838 1402
rect 2138 1350 2190 1402
rect 2490 1350 2542 1402
rect 3241 1287 3293 1339
rect 3305 1287 3357 1339
rect 3369 1287 3421 1339
rect 3433 1287 3485 1339
rect 3497 1287 3549 1339
rect 6750 1283 6802 1335
rect 6814 1283 6866 1335
rect 6878 1283 6930 1335
rect 6942 1283 6994 1335
rect 7006 1283 7058 1335
rect 220 1199 272 1212
rect 220 1165 232 1199
rect 232 1165 266 1199
rect 266 1165 272 1199
rect 220 1160 272 1165
rect 134 1055 186 1084
rect 134 1032 144 1055
rect 144 1032 178 1055
rect 178 1032 186 1055
rect 818 1160 870 1212
rect 994 1160 1046 1212
rect 1170 1160 1222 1212
rect 1346 1160 1398 1212
rect 1522 1160 1574 1212
rect 1698 1160 1750 1212
rect 1874 1160 1926 1212
rect 2050 1160 2102 1212
rect 2226 1160 2278 1212
rect 2402 1160 2454 1212
rect 904 1032 956 1084
rect 1256 1032 1308 1084
rect 1608 1032 1660 1084
rect 1960 1032 2012 1084
rect 2312 1032 2364 1084
<< metal2 >>
rect -1507 2104 314 3440
rect 696 2104 2517 3455
rect -1557 2098 387 2104
rect -1557 2046 -1452 2098
rect -1400 2046 -1100 2098
rect -1048 2046 -748 2098
rect -696 2046 -396 2098
rect -344 2046 -44 2098
rect 8 2046 308 2098
rect 360 2046 387 2098
rect -1557 2040 387 2046
rect 679 2098 2608 2104
rect 679 2046 730 2098
rect 782 2046 1082 2098
rect 1134 2046 1434 2098
rect 1486 2046 1786 2098
rect 1838 2046 2138 2098
rect 2190 2046 2490 2098
rect 2542 2046 2608 2098
rect 679 2040 2608 2046
rect -1370 1910 366 1916
rect -5842 1856 -1905 1878
rect -5842 1853 -2271 1856
rect -5842 1801 -5747 1853
rect -5695 1801 -5683 1853
rect -5631 1801 -5619 1853
rect -5567 1801 -5555 1853
rect -5503 1801 -5491 1853
rect -5439 1804 -2271 1853
rect -2219 1804 -2207 1856
rect -2155 1804 -2143 1856
rect -2091 1804 -2079 1856
rect -2027 1804 -2015 1856
rect -1963 1804 -1905 1856
rect -1370 1858 -1364 1910
rect -1312 1858 -1188 1910
rect -1136 1858 -1012 1910
rect -960 1858 -836 1910
rect -784 1858 -660 1910
rect -608 1858 -484 1910
rect -432 1858 -308 1910
rect -256 1858 -132 1910
rect -80 1858 44 1910
rect 96 1858 220 1910
rect 272 1858 366 1910
rect -1370 1852 366 1858
rect 724 1910 2460 1916
rect 724 1858 818 1910
rect 870 1858 994 1910
rect 1046 1858 1170 1910
rect 1222 1858 1346 1910
rect 1398 1858 1522 1910
rect 1574 1858 1698 1910
rect 1750 1858 1874 1910
rect 1926 1858 2050 1910
rect 2102 1858 2226 1910
rect 2278 1858 2402 1910
rect 2454 1858 2460 1910
rect 724 1852 2460 1858
rect 3182 1889 7119 1911
rect 3182 1837 3240 1889
rect 3292 1837 3304 1889
rect 3356 1837 3368 1889
rect 3420 1837 3432 1889
rect 3484 1837 3496 1889
rect 3548 1886 7119 1889
rect 3548 1837 6716 1886
rect 3182 1834 6716 1837
rect 6768 1834 6780 1886
rect 6832 1834 6844 1886
rect 6896 1834 6908 1886
rect 6960 1834 6972 1886
rect 7024 1834 7119 1886
rect 3182 1815 7119 1834
rect -5439 1801 -1905 1804
rect -5842 1782 -1905 1801
rect 374 1650 734 1651
rect -1278 1644 2368 1650
rect -1278 1592 -1272 1644
rect -1220 1592 -920 1644
rect -868 1592 -568 1644
rect -516 1592 -216 1644
rect -164 1592 136 1644
rect 188 1592 902 1644
rect 954 1592 1254 1644
rect 1306 1592 1606 1644
rect 1658 1592 1958 1644
rect 2010 1592 2310 1644
rect 2362 1592 2368 1644
rect -1278 1586 2368 1592
rect 374 1585 734 1586
rect -1458 1402 366 1408
rect -1458 1350 -1452 1402
rect -1400 1350 -1100 1402
rect -1048 1350 -748 1402
rect -696 1350 -396 1402
rect -344 1350 -44 1402
rect 8 1350 308 1402
rect 360 1350 366 1402
rect -1458 1344 366 1350
rect 724 1402 2548 1408
rect 724 1350 730 1402
rect 782 1350 1082 1402
rect 1134 1350 1434 1402
rect 1486 1350 1786 1402
rect 1838 1350 2138 1402
rect 2190 1350 2490 1402
rect 2542 1350 2548 1402
rect 724 1344 2548 1350
rect 3181 1339 7118 1361
rect -5841 1306 -1904 1328
rect -5841 1302 -2272 1306
rect -5841 1250 -5781 1302
rect -5729 1250 -5717 1302
rect -5665 1250 -5653 1302
rect -5601 1250 -5589 1302
rect -5537 1250 -5525 1302
rect -5473 1254 -2272 1302
rect -2220 1254 -2208 1306
rect -2156 1254 -2144 1306
rect -2092 1254 -2080 1306
rect -2028 1254 -2016 1306
rect -1964 1254 -1904 1306
rect 3181 1287 3241 1339
rect 3293 1287 3305 1339
rect 3357 1287 3369 1339
rect 3421 1287 3433 1339
rect 3485 1287 3497 1339
rect 3549 1335 7118 1339
rect 3549 1287 6750 1335
rect 3181 1283 6750 1287
rect 6802 1283 6814 1335
rect 6866 1283 6878 1335
rect 6930 1283 6942 1335
rect 6994 1283 7006 1335
rect 7058 1283 7118 1335
rect 3181 1265 7118 1283
rect -5473 1250 -1904 1254
rect -5841 1232 -1904 1250
rect -1370 1212 278 1218
rect -1370 1160 -1364 1212
rect -1312 1160 -1188 1212
rect -1136 1160 -1012 1212
rect -960 1160 -836 1212
rect -784 1160 -660 1212
rect -608 1160 -484 1212
rect -432 1160 -308 1212
rect -256 1160 -132 1212
rect -80 1160 44 1212
rect 96 1160 220 1212
rect 272 1160 278 1212
rect -1370 1154 278 1160
rect 812 1212 2460 1218
rect 812 1160 818 1212
rect 870 1160 994 1212
rect 1046 1160 1170 1212
rect 1222 1160 1346 1212
rect 1398 1160 1522 1212
rect 1574 1160 1698 1212
rect 1750 1160 1874 1212
rect 1926 1160 2050 1212
rect 2102 1160 2226 1212
rect 2278 1160 2402 1212
rect 2454 1160 2460 1212
rect 812 1154 2460 1160
rect -1279 1084 2369 1090
rect -1279 1032 -1274 1084
rect -1222 1032 -922 1084
rect -870 1032 -570 1084
rect -518 1032 -218 1084
rect -166 1032 134 1084
rect 186 1032 904 1084
rect 956 1032 1256 1084
rect 1308 1032 1608 1084
rect 1660 1032 1960 1084
rect 2012 1032 2312 1084
rect 2364 1032 2369 1084
rect -1279 1026 2369 1032
rect -441 -129 840 1026
use sky130_fd_pr__res_xhigh_po_0p35_9FS993  sky130_fd_pr__res_xhigh_po_0p35_9FS993_5
timestamp 1636132012
transform 0 1 -3869 -1 0 1582
box -191 -2088 191 2088
use sky130_fd_pr__res_xhigh_po_0p35_9FS993  sky130_fd_pr__res_xhigh_po_0p35_9FS993_4
timestamp 1636132012
transform 0 1 -3908 -1 0 1043
box -191 -2088 191 2088
use sky130_fd_pr__res_xhigh_po_0p35_9FS993  sky130_fd_pr__res_xhigh_po_0p35_9FS993_3
timestamp 1636132012
transform 0 1 -3864 -1 0 2091
box -191 -2088 191 2088
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_18
timestamp 1636132012
transform 1 0 885 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_19
timestamp 1636132012
transform 1 0 797 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_16
timestamp 1636132012
transform 1 0 1061 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_17
timestamp 1636132012
transform 1 0 973 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_13
timestamp 1636132012
transform 1 0 1237 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_14
timestamp 1636132012
transform 1 0 1149 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_15
timestamp 1636132012
transform 1 0 1325 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_11
timestamp 1636132012
transform 1 0 1413 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_12
timestamp 1636132012
transform 1 0 1501 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_8
timestamp 1636132012
transform 1 0 1589 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_9
timestamp 1636132012
transform 1 0 1677 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_10
timestamp 1636132012
transform 1 0 1765 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_6
timestamp 1636132012
transform 1 0 1941 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_7
timestamp 1636132012
transform 1 0 1853 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_3
timestamp 1636132012
transform 1 0 2029 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_4
timestamp 1636132012
transform 1 0 2117 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_5
timestamp 1636132012
transform 1 0 2205 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_1
timestamp 1636132012
transform 1 0 2293 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_2
timestamp 1636132012
transform 1 0 2381 0 1 1506
box -99 -626 99 626
use sky130_fd_pr__res_xhigh_po_0p35_9FS993  sky130_fd_pr__res_xhigh_po_0p35_9FS993_2
timestamp 1636132012
transform 0 1 5185 -1 0 1076
box -191 -2088 191 2088
use sky130_fd_pr__res_xhigh_po_0p35_9FS993  sky130_fd_pr__res_xhigh_po_0p35_9FS993_1
timestamp 1636132012
transform 0 1 5146 -1 0 1615
box -191 -2088 191 2088
use sky130_fd_pr__res_xhigh_po_0p35_9FS993  sky130_fd_pr__res_xhigh_po_0p35_9FS993_0
timestamp 1636132012
transform 0 1 5141 -1 0 2124
box -191 -2088 191 2088
use sky130_fd_pr__nfet_01v8_lvt_HYBPL5  sky130_fd_pr__nfet_01v8_lvt_HYBPL5_0
timestamp 1636132012
transform 1 0 2469 0 1 1506
box -99 -626 99 626
<< labels >>
rlabel metal1 s -6206 1584 -6206 1584 4 VSWN
port 1 nsew
rlabel metal1 s 7412 1617 7412 1617 4 VSWP
port 2 nsew
rlabel metal2 s -709 3384 -709 3384 4 VPA
port 3 nsew
rlabel metal2 s 1600 3435 1600 3435 4 VLNA
port 4 nsew
rlabel metal2 s 156 -127 156 -127 4 VO2
port 5 nsew
rlabel locali s 2981 2292 2981 2292 4 VSS
port 6 nsew
<< end >>
