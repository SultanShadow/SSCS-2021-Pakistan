magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< nwell >>
rect -738 -738 738 738
<< pwell >>
rect -866 780 866 866
rect -866 -780 -780 780
rect 780 -780 866 780
rect -866 -866 866 -780
<< psubdiff >>
rect -840 806 -731 840
rect -697 806 -663 840
rect -629 806 -595 840
rect -561 806 -527 840
rect -493 806 -459 840
rect -425 806 -391 840
rect -357 806 -323 840
rect -289 806 -255 840
rect -221 806 -187 840
rect -153 806 -119 840
rect -85 806 -51 840
rect -17 806 17 840
rect 51 806 85 840
rect 119 806 153 840
rect 187 806 221 840
rect 255 806 289 840
rect 323 806 357 840
rect 391 806 425 840
rect 459 806 493 840
rect 527 806 561 840
rect 595 806 629 840
rect 663 806 697 840
rect 731 806 840 840
rect -840 731 -806 806
rect 806 731 840 806
rect -840 663 -806 697
rect -840 595 -806 629
rect -840 527 -806 561
rect -840 459 -806 493
rect -840 391 -806 425
rect -840 323 -806 357
rect -840 255 -806 289
rect -840 187 -806 221
rect -840 119 -806 153
rect -840 51 -806 85
rect -840 -17 -806 17
rect -840 -85 -806 -51
rect -840 -153 -806 -119
rect -840 -221 -806 -187
rect -840 -289 -806 -255
rect -840 -357 -806 -323
rect -840 -425 -806 -391
rect -840 -493 -806 -459
rect -840 -561 -806 -527
rect -840 -629 -806 -595
rect -840 -697 -806 -663
rect 806 663 840 697
rect 806 595 840 629
rect 806 527 840 561
rect 806 459 840 493
rect 806 391 840 425
rect 806 323 840 357
rect 806 255 840 289
rect 806 187 840 221
rect 806 119 840 153
rect 806 51 840 85
rect 806 -17 840 17
rect 806 -85 840 -51
rect 806 -153 840 -119
rect 806 -221 840 -187
rect 806 -289 840 -255
rect 806 -357 840 -323
rect 806 -425 840 -391
rect 806 -493 840 -459
rect 806 -561 840 -527
rect 806 -629 840 -595
rect 806 -697 840 -663
rect -840 -806 -806 -731
rect 806 -806 840 -731
rect -840 -840 -731 -806
rect -697 -840 -663 -806
rect -629 -840 -595 -806
rect -561 -840 -527 -806
rect -493 -840 -459 -806
rect -425 -840 -391 -806
rect -357 -840 -323 -806
rect -289 -840 -255 -806
rect -221 -840 -187 -806
rect -153 -840 -119 -806
rect -85 -840 -51 -806
rect -17 -840 17 -806
rect 51 -840 85 -806
rect 119 -840 153 -806
rect 187 -840 221 -806
rect 255 -840 289 -806
rect 323 -840 357 -806
rect 391 -840 425 -806
rect 459 -840 493 -806
rect 527 -840 561 -806
rect 595 -840 629 -806
rect 663 -840 697 -806
rect 731 -840 840 -806
<< nsubdiff >>
rect -702 668 -595 702
rect -561 668 -527 702
rect -493 668 -459 702
rect -425 668 -391 702
rect -357 668 -323 702
rect -289 668 -255 702
rect -221 668 -187 702
rect -153 668 -119 702
rect -85 668 -51 702
rect -17 668 17 702
rect 51 668 85 702
rect 119 668 153 702
rect 187 668 221 702
rect 255 668 289 702
rect 323 668 357 702
rect 391 668 425 702
rect 459 668 493 702
rect 527 668 561 702
rect 595 668 702 702
rect -702 595 -668 668
rect -702 527 -668 561
rect -702 459 -668 493
rect -702 391 -668 425
rect -702 323 -668 357
rect -702 255 -668 289
rect -702 187 -668 221
rect -702 119 -668 153
rect -702 51 -668 85
rect -702 -17 -668 17
rect -702 -85 -668 -51
rect -702 -153 -668 -119
rect -702 -221 -668 -187
rect -702 -289 -668 -255
rect -702 -357 -668 -323
rect -702 -425 -668 -391
rect -702 -493 -668 -459
rect -702 -561 -668 -527
rect -702 -668 -668 -595
rect 668 595 702 668
rect 668 527 702 561
rect 668 459 702 493
rect 668 391 702 425
rect 668 323 702 357
rect 668 255 702 289
rect 668 187 702 221
rect 668 119 702 153
rect 668 51 702 85
rect 668 -17 702 17
rect 668 -85 702 -51
rect 668 -153 702 -119
rect 668 -221 702 -187
rect 668 -289 702 -255
rect 668 -357 702 -323
rect 668 -425 702 -391
rect 668 -493 702 -459
rect 668 -561 702 -527
rect 668 -668 702 -595
rect -702 -702 -595 -668
rect -561 -702 -527 -668
rect -493 -702 -459 -668
rect -425 -702 -391 -668
rect -357 -702 -323 -668
rect -289 -702 -255 -668
rect -221 -702 -187 -668
rect -153 -702 -119 -668
rect -85 -702 -51 -668
rect -17 -702 17 -668
rect 51 -702 85 -668
rect 119 -702 153 -668
rect 187 -702 221 -668
rect 255 -702 289 -668
rect 323 -702 357 -668
rect 391 -702 425 -668
rect 459 -702 493 -668
rect 527 -702 561 -668
rect 595 -702 702 -668
<< psubdiffcont >>
rect -731 806 -697 840
rect -663 806 -629 840
rect -595 806 -561 840
rect -527 806 -493 840
rect -459 806 -425 840
rect -391 806 -357 840
rect -323 806 -289 840
rect -255 806 -221 840
rect -187 806 -153 840
rect -119 806 -85 840
rect -51 806 -17 840
rect 17 806 51 840
rect 85 806 119 840
rect 153 806 187 840
rect 221 806 255 840
rect 289 806 323 840
rect 357 806 391 840
rect 425 806 459 840
rect 493 806 527 840
rect 561 806 595 840
rect 629 806 663 840
rect 697 806 731 840
rect -840 697 -806 731
rect -840 629 -806 663
rect -840 561 -806 595
rect -840 493 -806 527
rect -840 425 -806 459
rect -840 357 -806 391
rect -840 289 -806 323
rect -840 221 -806 255
rect -840 153 -806 187
rect -840 85 -806 119
rect -840 17 -806 51
rect -840 -51 -806 -17
rect -840 -119 -806 -85
rect -840 -187 -806 -153
rect -840 -255 -806 -221
rect -840 -323 -806 -289
rect -840 -391 -806 -357
rect -840 -459 -806 -425
rect -840 -527 -806 -493
rect -840 -595 -806 -561
rect -840 -663 -806 -629
rect -840 -731 -806 -697
rect 806 697 840 731
rect 806 629 840 663
rect 806 561 840 595
rect 806 493 840 527
rect 806 425 840 459
rect 806 357 840 391
rect 806 289 840 323
rect 806 221 840 255
rect 806 153 840 187
rect 806 85 840 119
rect 806 17 840 51
rect 806 -51 840 -17
rect 806 -119 840 -85
rect 806 -187 840 -153
rect 806 -255 840 -221
rect 806 -323 840 -289
rect 806 -391 840 -357
rect 806 -459 840 -425
rect 806 -527 840 -493
rect 806 -595 840 -561
rect 806 -663 840 -629
rect 806 -731 840 -697
rect -731 -840 -697 -806
rect -663 -840 -629 -806
rect -595 -840 -561 -806
rect -527 -840 -493 -806
rect -459 -840 -425 -806
rect -391 -840 -357 -806
rect -323 -840 -289 -806
rect -255 -840 -221 -806
rect -187 -840 -153 -806
rect -119 -840 -85 -806
rect -51 -840 -17 -806
rect 17 -840 51 -806
rect 85 -840 119 -806
rect 153 -840 187 -806
rect 221 -840 255 -806
rect 289 -840 323 -806
rect 357 -840 391 -806
rect 425 -840 459 -806
rect 493 -840 527 -806
rect 561 -840 595 -806
rect 629 -840 663 -806
rect 697 -840 731 -806
<< nsubdiffcont >>
rect -595 668 -561 702
rect -527 668 -493 702
rect -459 668 -425 702
rect -391 668 -357 702
rect -323 668 -289 702
rect -255 668 -221 702
rect -187 668 -153 702
rect -119 668 -85 702
rect -51 668 -17 702
rect 17 668 51 702
rect 85 668 119 702
rect 153 668 187 702
rect 221 668 255 702
rect 289 668 323 702
rect 357 668 391 702
rect 425 668 459 702
rect 493 668 527 702
rect 561 668 595 702
rect -702 561 -668 595
rect -702 493 -668 527
rect -702 425 -668 459
rect -702 357 -668 391
rect -702 289 -668 323
rect -702 221 -668 255
rect -702 153 -668 187
rect -702 85 -668 119
rect -702 17 -668 51
rect -702 -51 -668 -17
rect -702 -119 -668 -85
rect -702 -187 -668 -153
rect -702 -255 -668 -221
rect -702 -323 -668 -289
rect -702 -391 -668 -357
rect -702 -459 -668 -425
rect -702 -527 -668 -493
rect -702 -595 -668 -561
rect 668 561 702 595
rect 668 493 702 527
rect 668 425 702 459
rect 668 357 702 391
rect 668 289 702 323
rect 668 221 702 255
rect 668 153 702 187
rect 668 85 702 119
rect 668 17 702 51
rect 668 -51 702 -17
rect 668 -119 702 -85
rect 668 -187 702 -153
rect 668 -255 702 -221
rect 668 -323 702 -289
rect 668 -391 702 -357
rect 668 -459 702 -425
rect 668 -527 702 -493
rect 668 -595 702 -561
rect -595 -702 -561 -668
rect -527 -702 -493 -668
rect -459 -702 -425 -668
rect -391 -702 -357 -668
rect -323 -702 -289 -668
rect -255 -702 -221 -668
rect -187 -702 -153 -668
rect -119 -702 -85 -668
rect -51 -702 -17 -668
rect 17 -702 51 -668
rect 85 -702 119 -668
rect 153 -702 187 -668
rect 221 -702 255 -668
rect 289 -702 323 -668
rect 357 -702 391 -668
rect 425 -702 459 -668
rect 493 -702 527 -668
rect 561 -702 595 -668
<< pdiode >>
rect -600 561 600 600
rect -600 -561 -561 561
rect 561 -561 600 561
rect -600 -600 600 -561
<< pdiodec >>
rect -561 -561 561 561
<< locali >>
rect -840 806 -731 840
rect -697 806 -663 840
rect -629 806 -595 840
rect -561 806 -527 840
rect -493 806 -459 840
rect -425 806 -391 840
rect -357 806 -323 840
rect -289 806 -255 840
rect -221 806 -187 840
rect -153 806 -119 840
rect -85 806 -51 840
rect -17 806 17 840
rect 51 806 85 840
rect 119 806 153 840
rect 187 806 221 840
rect 255 806 289 840
rect 323 806 357 840
rect 391 806 425 840
rect 459 806 493 840
rect 527 806 561 840
rect 595 806 629 840
rect 663 806 697 840
rect 731 806 840 840
rect -840 731 -806 806
rect 806 731 840 806
rect -840 663 -806 697
rect -840 595 -806 629
rect -840 527 -806 561
rect -840 459 -806 493
rect -840 391 -806 425
rect -840 323 -806 357
rect -840 255 -806 289
rect -840 187 -806 221
rect -840 119 -806 153
rect -840 51 -806 85
rect -840 -17 -806 17
rect -840 -85 -806 -51
rect -840 -153 -806 -119
rect -840 -221 -806 -187
rect -840 -289 -806 -255
rect -840 -357 -806 -323
rect -840 -425 -806 -391
rect -840 -493 -806 -459
rect -840 -561 -806 -527
rect -840 -629 -806 -595
rect -840 -697 -806 -663
rect -702 668 -595 702
rect -561 668 -527 702
rect -493 668 -459 702
rect -425 668 -391 702
rect -357 668 -323 702
rect -289 668 -255 702
rect -221 668 -187 702
rect -153 668 -119 702
rect -85 668 -51 702
rect -17 668 17 702
rect 51 668 85 702
rect 119 668 153 702
rect 187 668 221 702
rect 255 668 289 702
rect 323 668 357 702
rect 391 668 425 702
rect 459 668 493 702
rect 527 668 561 702
rect 595 668 702 702
rect -702 595 -668 668
rect 668 595 702 668
rect -702 527 -668 561
rect -702 459 -668 493
rect -702 391 -668 425
rect -702 323 -668 357
rect -702 255 -668 289
rect -702 187 -668 221
rect -702 119 -668 153
rect -702 51 -668 85
rect -702 -17 -668 17
rect -702 -85 -668 -51
rect -702 -153 -668 -119
rect -702 -221 -668 -187
rect -702 -289 -668 -255
rect -702 -357 -668 -323
rect -702 -425 -668 -391
rect -702 -493 -668 -459
rect -702 -561 -668 -527
rect -604 561 604 588
rect -604 -561 -561 561
rect 561 -561 604 561
rect -604 -588 604 -561
rect 668 527 702 561
rect 668 459 702 493
rect 668 391 702 425
rect 668 323 702 357
rect 668 255 702 289
rect 668 187 702 221
rect 668 119 702 153
rect 668 51 702 85
rect 668 -17 702 17
rect 668 -85 702 -51
rect 668 -153 702 -119
rect 668 -221 702 -187
rect 668 -289 702 -255
rect 668 -357 702 -323
rect 668 -425 702 -391
rect 668 -493 702 -459
rect 668 -561 702 -527
rect -702 -668 -668 -595
rect 668 -668 702 -595
rect -702 -702 -595 -668
rect -561 -702 -527 -668
rect -493 -702 -459 -668
rect -425 -702 -391 -668
rect -357 -702 -323 -668
rect -289 -702 -255 -668
rect -221 -702 -187 -668
rect -153 -702 -119 -668
rect -85 -702 -51 -668
rect -17 -702 17 -668
rect 51 -702 85 -668
rect 119 -702 153 -668
rect 187 -702 221 -668
rect 255 -702 289 -668
rect 323 -702 357 -668
rect 391 -702 425 -668
rect 459 -702 493 -668
rect 527 -702 561 -668
rect 595 -702 702 -668
rect 806 663 840 697
rect 806 595 840 629
rect 806 527 840 561
rect 806 459 840 493
rect 806 391 840 425
rect 806 323 840 357
rect 806 255 840 289
rect 806 187 840 221
rect 806 119 840 153
rect 806 51 840 85
rect 806 -17 840 17
rect 806 -85 840 -51
rect 806 -153 840 -119
rect 806 -221 840 -187
rect 806 -289 840 -255
rect 806 -357 840 -323
rect 806 -425 840 -391
rect 806 -493 840 -459
rect 806 -561 840 -527
rect 806 -629 840 -595
rect 806 -697 840 -663
rect -840 -806 -806 -731
rect 806 -806 840 -731
rect -840 -840 -731 -806
rect -697 -840 -663 -806
rect -629 -840 -595 -806
rect -561 -840 -527 -806
rect -493 -840 -459 -806
rect -425 -840 -391 -806
rect -357 -840 -323 -806
rect -289 -840 -255 -806
rect -221 -840 -187 -806
rect -153 -840 -119 -806
rect -85 -840 -51 -806
rect -17 -840 17 -806
rect 51 -840 85 -806
rect 119 -840 153 -806
rect 187 -840 221 -806
rect 255 -840 289 -806
rect 323 -840 357 -806
rect 391 -840 425 -806
rect 459 -840 493 -806
rect 527 -840 561 -806
rect 595 -840 629 -806
rect 663 -840 697 -806
rect 731 -840 840 -806
<< viali >>
rect -557 -557 557 557
<< metal1 >>
rect -600 557 600 594
rect -600 -557 -557 557
rect 557 -557 600 557
rect -600 -594 600 -557
<< properties >>
string FIXED_BBOX -684 -684 684 684
<< end >>
