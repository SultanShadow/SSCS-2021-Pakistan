magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< error_s >>
rect 3964 12507 4500 12828
<< locali >>
rect 5324 29133 10352 29402
rect 5324 28163 6301 29133
rect 9647 28163 10352 29133
rect 5324 23200 10352 28163
rect 6226 23152 6638 23200
rect 3030 12461 4049 12511
rect 4383 12504 4864 12583
rect 4383 12470 4787 12504
rect 4821 12470 4864 12504
rect 3030 12389 3666 12461
rect 4383 12391 4864 12470
rect 3030 12283 3112 12389
rect 3578 12283 3666 12389
rect 3030 12228 3666 12283
rect 4001 12048 5024 12133
rect 4001 11798 4108 12048
rect 4358 11798 5024 12048
rect 4001 11734 5024 11798
rect -7302 10714 9516 10756
rect -7302 10300 23531 10714
rect -7302 8970 -6933 10300
rect -5675 8970 23531 10300
rect -7302 8618 23531 8970
rect 8218 8576 23531 8618
rect 7674 -288 8877 660
rect 7674 -1042 7858 -288
rect 8684 -1042 8877 -288
rect 7674 -1178 8877 -1042
rect 21480 108 22336 1455
rect 21480 -1078 21589 108
rect 22199 -1078 22336 108
rect 21480 -1179 22336 -1078
<< viali >>
rect 6301 28163 9647 29133
rect 4787 12470 4821 12504
rect 3112 12283 3578 12389
rect 4108 11798 4358 12048
rect -6933 8970 -5675 10300
rect 7858 -1042 8684 -288
rect 21589 -1078 22199 108
<< metal1 >>
rect 30188 29382 32214 29394
rect -7310 29152 32214 29382
rect -7310 28140 -6964 29152
rect -5824 29146 32214 29152
rect -5824 29133 30680 29146
rect -5824 28163 6301 29133
rect 9647 29108 30680 29133
rect 9647 28224 18979 29108
rect 21719 28224 30680 29108
rect 9647 28163 30680 28224
rect -5824 28140 30680 28163
rect -7310 28134 30680 28140
rect 31820 28134 32214 29146
rect -7310 27836 32214 28134
rect 15884 21135 16300 21189
rect 15884 20955 15969 21135
rect 16213 20955 16300 21135
rect 15884 20895 16300 20955
rect 20915 19274 22365 19634
rect 20915 16278 21273 19274
rect 22029 16278 22365 19274
rect 20915 15825 22365 16278
rect 2923 13188 4253 13272
rect 2923 12944 3142 13188
rect 4090 12944 4253 13188
rect 2923 12757 4253 12944
rect 18333 12758 18962 12797
rect 18333 12629 18963 12758
rect 4770 12504 4838 12537
rect 4770 12470 4787 12504
rect 4821 12470 4838 12504
rect 3030 12389 3666 12461
rect 4770 12437 4838 12470
rect 18333 12449 18531 12629
rect 18839 12449 18963 12629
rect 3030 12283 3112 12389
rect 3578 12283 3666 12389
rect 18333 12318 18963 12449
rect 3030 11511 3666 12283
rect 4001 12048 4459 12293
rect 4001 11798 4108 12048
rect 4358 11798 4459 12048
rect 4001 11734 4459 11798
rect 18333 11511 18962 12318
rect 3029 10886 18962 11511
rect 3029 10879 18943 10886
rect -7308 10301 -5274 10762
rect -7308 8969 -6938 10301
rect -5670 8969 -5274 10301
rect -7308 8618 -5274 8969
rect 27370 8966 28382 8974
rect 25680 8836 28382 8966
rect 25680 8208 27544 8836
rect 28236 8208 28382 8836
rect 25680 8082 28382 8208
rect 25680 8078 28024 8082
rect 6607 4555 7117 4655
rect 6607 4247 6677 4555
rect 7049 4247 7117 4555
rect 6607 4148 7117 4247
rect 11396 3724 12214 3838
rect 8172 3484 10959 3712
rect 8172 3242 8354 3484
rect 8171 3048 8354 3242
rect 10710 3048 10959 3484
rect 11396 3352 11567 3724
rect 12067 3352 12214 3724
rect 11396 3184 12214 3352
rect 8171 2840 10959 3048
rect 11397 3011 11958 3184
rect 11397 2526 11960 3011
rect 10473 1488 13158 1572
rect 10473 1308 12456 1488
rect 13020 1308 13158 1488
rect 10473 1218 13158 1308
rect 23378 1368 25246 1477
rect 23378 1124 23520 1368
rect 25044 1124 25246 1368
rect 23378 1019 25246 1124
rect 30190 372 32216 378
rect -7296 108 32216 372
rect -7296 100 21589 108
rect -7296 -912 -6904 100
rect -5764 -288 21589 100
rect -5764 -912 7858 -288
rect -7296 -1042 7858 -912
rect 8684 -1042 21589 -288
rect -7296 -1078 21589 -1042
rect 22199 72 32216 108
rect 22199 -940 30604 72
rect 31744 -940 32216 72
rect 22199 -1078 32216 -940
rect -7296 -1174 32216 -1078
rect 30190 -1180 32216 -1174
<< via1 >>
rect -6964 28140 -5824 29152
rect 18979 28224 21719 29108
rect 30680 28134 31820 29146
rect 15969 20955 16213 21135
rect 21273 16278 22029 19274
rect 3142 12944 4090 13188
rect 18531 12449 18839 12629
rect -6938 10300 -5670 10301
rect -6938 8970 -6933 10300
rect -6933 8970 -5675 10300
rect -5675 8970 -5670 10300
rect -6938 8969 -5670 8970
rect 27544 8208 28236 8836
rect 6677 4247 7049 4555
rect 8354 3048 10710 3484
rect 11567 3352 12067 3724
rect 12456 1308 13020 1488
rect 23520 1124 25044 1368
rect -6904 -912 -5764 100
rect 30604 -940 31744 72
<< metal2 >>
rect -7296 29152 -5274 29380
rect -7296 28140 -6964 29152
rect -5824 28140 -5274 29152
rect -7296 24953 -5274 28140
rect 18533 29108 22118 29379
rect 18533 28224 18979 29108
rect 21719 28224 22118 29108
rect 18533 27839 22118 28224
rect 30190 29146 32212 29374
rect 30190 28134 30680 29146
rect 31820 28134 32212 29146
rect -7296 24737 -7149 24953
rect -5413 24737 -5274 24953
rect -7296 18779 -5274 24737
rect 30190 26497 32212 28134
rect 11285 23133 14713 23535
rect 2743 22954 3419 23096
rect 2743 22018 2936 22954
rect 3232 22018 3419 22954
rect 2743 21850 3419 22018
rect 6660 21924 8416 21933
rect -7296 15203 -6705 18779
rect -5849 15203 -5274 18779
rect 1846 18900 2750 19395
rect 1846 16044 2200 18900
rect 2576 18496 2750 18900
rect 6716 18496 8416 21924
rect 11285 21797 11770 23133
rect 14386 21797 14713 23133
rect 18940 21933 22446 22596
rect 11285 21473 14713 21797
rect 18840 21887 22446 21933
rect 16636 21189 17625 21254
rect 15884 21135 16300 21189
rect 15884 21113 15969 21135
rect 16213 21113 16300 21135
rect 15884 20977 15943 21113
rect 16239 20977 16300 21113
rect 15884 20955 15969 20977
rect 16213 20955 16300 20977
rect 15884 20895 16300 20955
rect 16636 20973 16790 21189
rect 17486 20973 17625 21189
rect 16636 20914 17625 20973
rect 18840 20471 19520 21887
rect 21896 20471 22446 21887
rect 18840 20227 22446 20471
rect 18940 20156 22446 20227
rect 2576 16044 8416 18496
rect 1846 16008 8416 16044
rect 1846 15796 2750 16008
rect -7296 10301 -5274 15203
rect 2924 13188 4251 16008
rect 6716 16001 8416 16008
rect 20915 19284 22365 19634
rect 20915 16268 21263 19284
rect 22039 16268 22365 19284
rect 20915 15825 22365 16268
rect 30190 16121 30608 26497
rect 31784 16121 32212 26497
rect 2924 12944 3142 13188
rect 4090 12944 4251 13188
rect 2924 12846 4251 12944
rect 27161 12842 27959 13004
rect 27161 12781 27310 12842
rect 18388 12758 27310 12781
rect 18336 12629 27310 12758
rect 18336 12449 18531 12629
rect 18839 12449 27310 12629
rect 18336 12347 27310 12449
rect 18336 12318 18963 12347
rect 27161 12226 27310 12347
rect 27846 12226 27959 12842
rect 27161 12053 27959 12226
rect -7296 8969 -6938 10301
rect -5670 8969 -5274 10301
rect -7296 100 -5274 8969
rect 27370 8836 28382 8974
rect 27370 8830 27544 8836
rect 28236 8830 28382 8836
rect 27370 8214 27542 8830
rect 28238 8214 28382 8830
rect 27370 8208 27544 8214
rect 28236 8208 28382 8214
rect 27370 8082 28382 8208
rect -1767 4880 7109 5042
rect -1767 3784 -1614 4880
rect -838 4655 7109 4880
rect -838 4555 7117 4655
rect -838 4247 6677 4555
rect 7049 4247 7117 4555
rect -838 4148 7117 4247
rect -838 3784 7109 4148
rect -1767 3619 7109 3784
rect 11396 3726 12214 3838
rect 11396 3724 11589 3726
rect 12045 3724 12214 3726
rect 7879 3494 10928 3711
rect 7879 3038 8344 3494
rect 10720 3038 10928 3494
rect 11396 3352 11567 3724
rect 12067 3352 12214 3724
rect 11396 3350 11589 3352
rect 12045 3350 12214 3352
rect 11396 3184 12214 3350
rect 7879 2663 10928 3038
rect 12233 1506 13157 1581
rect 12233 1488 12470 1506
rect 13006 1488 13157 1506
rect 12233 1308 12456 1488
rect 13020 1308 13157 1488
rect 12233 1290 12470 1308
rect 13006 1290 13157 1308
rect 12233 1220 13157 1290
rect 23378 1368 25246 1477
rect 23378 1124 23520 1368
rect 25044 1124 25246 1368
rect 23378 1019 25246 1124
rect -7296 -912 -6904 100
rect -5764 -912 -5274 100
rect -7296 -1174 -5274 -912
rect 30190 72 32212 16121
rect 30190 -940 30604 72
rect 31744 -940 32212 72
rect 30190 -1180 32212 -940
<< via2 >>
rect 19001 28238 21697 29094
rect -7149 24737 -5413 24953
rect 2936 22018 3232 22954
rect -6705 15203 -5849 18779
rect 2200 16044 2576 18900
rect 11770 21797 14386 23133
rect 15943 20977 15969 21113
rect 15969 20977 16213 21113
rect 16213 20977 16239 21113
rect 16790 20973 17486 21189
rect 19520 20471 21896 21887
rect 21263 19274 22039 19284
rect 21263 16278 21273 19274
rect 21273 16278 22029 19274
rect 22029 16278 22039 19274
rect 21263 16268 22039 16278
rect 30608 16121 31784 26497
rect 27310 12226 27846 12842
rect 27542 8214 27544 8830
rect 27544 8214 28236 8830
rect 28236 8214 28238 8830
rect -1614 3784 -838 4880
rect 11589 3724 12045 3726
rect 8344 3484 10720 3494
rect 8344 3048 8354 3484
rect 8354 3048 10710 3484
rect 10710 3048 10720 3484
rect 8344 3038 10720 3048
rect 11589 3352 12045 3724
rect 11589 3350 12045 3352
rect 12470 1488 13006 1506
rect 12470 1308 13006 1488
rect 12470 1290 13006 1308
rect 23534 1138 25030 1354
<< metal3 >>
rect 18533 29098 22118 29379
rect 11285 27509 14736 29001
rect 11285 26245 12018 27509
rect 14402 26245 14736 27509
rect -7296 24957 -5274 25050
rect -7296 24733 -7153 24957
rect -5409 24733 -5274 24957
rect -7296 24640 -5274 24733
rect 11285 23133 14736 26245
rect 2743 22954 3419 23094
rect 2743 22918 2936 22954
rect 3232 22918 3419 22954
rect 2743 22054 2932 22918
rect 3236 22054 3419 22918
rect 2743 22018 2936 22054
rect 3232 22018 3419 22054
rect 2743 21856 3419 22018
rect 11285 21797 11770 23133
rect 14386 21797 14736 23133
rect 11285 21467 14736 21797
rect 15828 21113 16402 28964
rect 15828 20977 15943 21113
rect 16239 20977 16402 21113
rect 15828 20900 16402 20977
rect 16631 21189 17701 28953
rect 18533 28234 18997 29098
rect 21701 28234 22118 29098
rect 18533 27839 22118 28234
rect 30195 26501 32232 27059
rect 16631 20973 16790 21189
rect 17486 20973 17701 21189
rect 16631 20912 17701 20973
rect 18940 21891 22446 22596
rect 18940 20467 19516 21891
rect 21900 20467 22446 21891
rect 18940 20156 22446 20467
rect -7296 18783 -5277 19251
rect -7296 15199 -6709 18783
rect -5845 15199 -5277 18783
rect 1846 18904 2750 19395
rect 1846 18900 2236 18904
rect 2540 18900 2750 18904
rect 1846 16044 2200 18900
rect 2576 16044 2750 18900
rect 1846 16040 2236 16044
rect 2540 16040 2750 16044
rect 1846 15796 2750 16040
rect 20915 19284 22365 19634
rect 20915 19248 21263 19284
rect 22039 19248 22365 19284
rect 20915 16304 21259 19248
rect 22043 16304 22365 19248
rect 20915 16268 21263 16304
rect 22039 16268 22365 16304
rect 20915 15825 22365 16268
rect 30195 16117 30604 26501
rect 31788 16117 32232 26501
rect 30195 15560 32232 16117
rect -7296 14641 -5277 15199
rect 27161 12846 27959 13004
rect 27161 12222 27306 12846
rect 27850 12222 27959 12846
rect 27161 12053 27959 12222
rect 27370 8834 28382 8974
rect 27370 8210 27538 8834
rect 28242 8210 28382 8834
rect 27370 8082 28382 8210
rect -1767 4884 -687 5043
rect -1767 3780 -1618 4884
rect -834 3780 -687 4884
rect 14244 3938 16344 3956
rect -1767 3619 -687 3780
rect 7869 3494 10935 3746
rect 7869 3038 8344 3494
rect 10720 3038 10935 3494
rect 11366 3726 16344 3938
rect 11366 3350 11589 3726
rect 12045 3350 16344 3726
rect 11366 3118 16344 3350
rect 7869 660 10935 3038
rect 7674 -1178 10935 660
rect 7869 -3656 10935 -1178
rect 12232 1506 13156 1578
rect 12232 1290 12470 1506
rect 13006 1290 13156 1506
rect 12232 -3745 13156 1290
rect 14244 -3770 16344 3118
rect 22920 1354 26368 1458
rect 22920 1138 23534 1354
rect 25030 1138 26368 1354
rect 22920 -3837 26368 1138
<< via3 >>
rect 12018 26245 14402 27509
rect -7153 24953 -5409 24957
rect -7153 24737 -7149 24953
rect -7149 24737 -5413 24953
rect -5413 24737 -5409 24953
rect -7153 24733 -5409 24737
rect 2932 22054 2936 22918
rect 2936 22054 3232 22918
rect 3232 22054 3236 22918
rect 18997 29094 21701 29098
rect 18997 28238 19001 29094
rect 19001 28238 21697 29094
rect 21697 28238 21701 29094
rect 18997 28234 21701 28238
rect 19516 21887 21900 21891
rect 19516 20471 19520 21887
rect 19520 20471 21896 21887
rect 21896 20471 21900 21887
rect 19516 20467 21900 20471
rect -6709 18779 -5845 18783
rect -6709 15203 -6705 18779
rect -6705 15203 -5849 18779
rect -5849 15203 -5845 18779
rect -6709 15199 -5845 15203
rect 2236 18900 2540 18904
rect 2236 16044 2540 18900
rect 2236 16040 2540 16044
rect 21259 16304 21263 19248
rect 21263 16304 22039 19248
rect 22039 16304 22043 19248
rect 30604 26497 31788 26501
rect 30604 16121 30608 26497
rect 30608 16121 31784 26497
rect 31784 16121 31788 26497
rect 30604 16117 31788 16121
rect 27306 12842 27850 12846
rect 27306 12226 27310 12842
rect 27310 12226 27846 12842
rect 27846 12226 27850 12842
rect 27306 12222 27850 12226
rect 27538 8830 28242 8834
rect 27538 8214 27542 8830
rect 27542 8214 28238 8830
rect 28238 8214 28242 8830
rect 27538 8210 28242 8214
rect -1618 4880 -834 4884
rect -1618 3784 -1614 4880
rect -1614 3784 -838 4880
rect -838 3784 -834 4880
rect -1618 3780 -834 3784
<< metal4 >>
rect 18533 29104 22118 29379
rect 18533 29098 19111 29104
rect 21587 29098 22118 29104
rect 18533 28234 18997 29098
rect 21701 28234 22118 29098
rect 18533 28228 19111 28234
rect 21587 28228 22118 28234
rect 11285 27509 14693 27889
rect 18533 27839 22118 28228
rect 11285 26245 12018 27509
rect 14402 26245 14693 27509
rect 11285 25939 14693 26245
rect 29224 26501 32219 27078
rect -7296 25049 133 25050
rect -7296 24957 10919 25049
rect -7296 24733 -7153 24957
rect -5409 24733 10919 24957
rect -7296 24640 10919 24733
rect -2861 23094 3407 24203
rect -2861 22918 3419 23094
rect -2861 22054 2932 22918
rect 3236 22054 3419 22918
rect -2861 21856 3419 22054
rect 18940 21891 22446 22596
rect -2861 20918 3407 21856
rect 18940 20467 19516 21891
rect 21900 20467 22446 21891
rect 18940 20156 22446 20467
rect -7296 18783 -5277 19251
rect -7296 18709 -6709 18783
rect -5845 18709 -5277 18783
rect -7296 15273 -6715 18709
rect -5839 15273 -5277 18709
rect 1846 18904 2750 19395
rect 1846 16040 2236 18904
rect 2540 16040 2750 18904
rect 1846 15796 2750 16040
rect 20915 19248 22365 19634
rect 20915 16304 21259 19248
rect 22043 16304 22365 19248
rect 20915 15825 22365 16304
rect 29224 16117 30604 26501
rect 31788 16117 32219 26501
rect 29224 15568 32219 16117
rect -7296 15199 -6709 15273
rect -5845 15199 -5277 15273
rect -7296 14641 -5277 15199
rect 27146 12846 33376 13190
rect 27146 12222 27306 12846
rect 27850 12222 33376 12846
rect 27146 11933 33376 12222
rect 27376 8974 33458 9464
rect 27370 8834 33458 8974
rect 27370 8210 27538 8834
rect 28242 8210 33458 8834
rect 27370 8082 33458 8210
rect 27376 8068 33458 8082
rect -4578 4884 -529 5491
rect -4578 3780 -1618 4884
rect -834 3780 -529 4884
rect -4578 3318 -529 3780
<< via4 >>
rect 19111 29098 21587 29104
rect 19111 28234 21587 29098
rect 19111 28228 21587 28234
rect 12132 26279 14288 27475
rect -6715 15273 -6709 18709
rect -6709 15273 -5845 18709
rect -5845 15273 -5839 18709
rect 21373 16378 21929 19174
<< metal5 >>
rect 18533 29227 22118 29379
rect 18533 29104 22119 29227
rect 18533 28228 19111 29104
rect 21587 28228 22119 29104
rect -4127 27475 14692 27889
rect 18533 27839 22119 28228
rect -4127 26279 12132 27475
rect 14288 26279 14692 27475
rect -4127 25939 14692 26279
rect 18534 23739 22119 27839
rect 28057 23466 28108 25536
rect 23659 19638 28108 23466
rect 29226 21832 29546 22199
rect -7296 18709 -327 19251
rect -7296 15273 -6715 18709
rect -5839 15273 -327 18709
rect 20930 19174 28108 19638
rect 20930 16378 21373 19174
rect 21929 17032 28108 19174
rect 21929 16378 28099 17032
rect 20930 15826 28099 16378
rect -7296 14641 -327 15273
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1636132012
transform 1 0 4002 0 1 12246
box -38 -48 498 592
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_1
timestamp 1636132012
transform 1 0 -1294 0 1 17068
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1636132012
transform 1 0 26173 0 1 18811
box -3351 -3101 3373 3101
use sky130_fd_pr__cap_mim_m3_2_S6VVQT  sky130_fd_pr__cap_mim_m3_2_S6VVQT_0
timestamp 1636132012
transform 1 0 26173 0 1 24752
box -3351 -2601 3373 2601
use sky130_fd_pr__cap_mim_m3_2_WXTTNJ  sky130_fd_pr__cap_mim_m3_2_WXTTNJ_0
timestamp 1636132012
transform 0 1 20351 -1 0 24648
box -2351 -2101 2373 2101
use sky130_fd_pr__cap_mim_m3_2_D7CHNQ  sky130_fd_pr__cap_mim_m3_2_D7CHNQ_3
timestamp 1636132012
transform 0 1 5470 -1 0 26628
box -1851 -1601 1873 1601
use sky130_fd_pr__cap_mim_m3_2_D7CHNQ  sky130_fd_pr__cap_mim_m3_2_D7CHNQ_2
timestamp 1636132012
transform 0 1 9319 -1 0 26607
box -1851 -1601 1873 1601
use sky130_fd_pr__cap_mim_m3_2_D7CHNQ  sky130_fd_pr__cap_mim_m3_2_D7CHNQ_1
timestamp 1636132012
transform 0 1 -3143 -1 0 26622
box -1851 -1601 1873 1601
use sky130_fd_pr__cap_mim_m3_2_D7CHNQ  sky130_fd_pr__cap_mim_m3_2_D7CHNQ_0
timestamp 1636132012
transform 0 1 1008 -1 0 26603
box -1851 -1601 1873 1601
use Top  Top_0
timestamp 1636132012
transform 1 0 0 0 1 1008
box 0 -1008 27865 22304
<< labels >>
flabel metal4 s -4562 4270 -4562 4270 0 FreeSans 24413 0 0 0 VCASC1
port 1 nsew
flabel metal3 s 9434 -3609 9434 -3609 0 FreeSans 24413 0 0 0 RFIN
port 2 nsew
flabel metal4 s 33320 12505 33320 12505 0 FreeSans 24413 0 0 0 VSWP
port 3 nsew
flabel metal4 s -2814 22609 -2814 22609 0 FreeSans 24413 0 0 0 PAOUT
port 4 nsew
flabel metal3 s 17133 28906 17133 28906 0 FreeSans 24413 90 0 0 LNAOUT
port 5 nsew
flabel metal3 s 15986 28874 15986 28874 0 FreeSans 9765 90 0 0 VBIAS4
port 6 nsew
flabel metal3 s 12963 28355 12963 28355 0 FreeSans 24413 90 0 0 VDD
port 7 nsew
flabel metal3 s 24438 -3432 24438 -3432 0 FreeSans 24413 0 0 0 VBIAS3
port 8 nsew
flabel metal3 s 12730 -3549 12730 -3549 0 FreeSans 14647 0 0 0 VBIAS2
port 9 nsew
flabel metal3 s 15458 -3736 15458 -3736 0 FreeSans 14647 0 0 0 VBIAS1
port 10 nsew
flabel metal4 s 33022 8740 33022 8740 0 FreeSans 24413 0 0 0 VCASC2
port 11 nsew
flabel metal1 s -3366 -795 -3366 -795 0 FreeSans 24413 0 0 0 VSS
port 12 nsew
<< end >>
