magic
tech sky130A
magscale 1 2
timestamp 1635855079
<< pwell >>
rect -191 2002 191 2088
rect -191 -2002 -105 2002
rect 105 -2002 191 2002
rect -191 -2088 191 -2002
<< psubdiff >>
rect -165 2028 -51 2062
rect -17 2028 17 2062
rect 51 2028 165 2062
rect -165 1955 -131 2028
rect 131 1955 165 2028
rect -165 1887 -131 1921
rect -165 1819 -131 1853
rect -165 1751 -131 1785
rect -165 1683 -131 1717
rect -165 1615 -131 1649
rect -165 1547 -131 1581
rect -165 1479 -131 1513
rect -165 1411 -131 1445
rect -165 1343 -131 1377
rect -165 1275 -131 1309
rect -165 1207 -131 1241
rect -165 1139 -131 1173
rect -165 1071 -131 1105
rect -165 1003 -131 1037
rect -165 935 -131 969
rect -165 867 -131 901
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect -165 -901 -131 -867
rect -165 -969 -131 -935
rect -165 -1037 -131 -1003
rect -165 -1105 -131 -1071
rect -165 -1173 -131 -1139
rect -165 -1241 -131 -1207
rect -165 -1309 -131 -1275
rect -165 -1377 -131 -1343
rect -165 -1445 -131 -1411
rect -165 -1513 -131 -1479
rect -165 -1581 -131 -1547
rect -165 -1649 -131 -1615
rect -165 -1717 -131 -1683
rect -165 -1785 -131 -1751
rect -165 -1853 -131 -1819
rect -165 -1921 -131 -1887
rect 131 1887 165 1921
rect 131 1819 165 1853
rect 131 1751 165 1785
rect 131 1683 165 1717
rect 131 1615 165 1649
rect 131 1547 165 1581
rect 131 1479 165 1513
rect 131 1411 165 1445
rect 131 1343 165 1377
rect 131 1275 165 1309
rect 131 1207 165 1241
rect 131 1139 165 1173
rect 131 1071 165 1105
rect 131 1003 165 1037
rect 131 935 165 969
rect 131 867 165 901
rect 131 799 165 833
rect 131 731 165 765
rect 131 663 165 697
rect 131 595 165 629
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -663
rect 131 -765 165 -731
rect 131 -833 165 -799
rect 131 -901 165 -867
rect 131 -969 165 -935
rect 131 -1037 165 -1003
rect 131 -1105 165 -1071
rect 131 -1173 165 -1139
rect 131 -1241 165 -1207
rect 131 -1309 165 -1275
rect 131 -1377 165 -1343
rect 131 -1445 165 -1411
rect 131 -1513 165 -1479
rect 131 -1581 165 -1547
rect 131 -1649 165 -1615
rect 131 -1717 165 -1683
rect 131 -1785 165 -1751
rect 131 -1853 165 -1819
rect 131 -1921 165 -1887
rect -165 -2028 -131 -1955
rect 131 -2028 165 -1955
rect -165 -2062 -51 -2028
rect -17 -2062 17 -2028
rect 51 -2062 165 -2028
<< psubdiffcont >>
rect -51 2028 -17 2062
rect 17 2028 51 2062
rect -165 1921 -131 1955
rect -165 1853 -131 1887
rect -165 1785 -131 1819
rect -165 1717 -131 1751
rect -165 1649 -131 1683
rect -165 1581 -131 1615
rect -165 1513 -131 1547
rect -165 1445 -131 1479
rect -165 1377 -131 1411
rect -165 1309 -131 1343
rect -165 1241 -131 1275
rect -165 1173 -131 1207
rect -165 1105 -131 1139
rect -165 1037 -131 1071
rect -165 969 -131 1003
rect -165 901 -131 935
rect -165 833 -131 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect -165 -867 -131 -833
rect -165 -935 -131 -901
rect -165 -1003 -131 -969
rect -165 -1071 -131 -1037
rect -165 -1139 -131 -1105
rect -165 -1207 -131 -1173
rect -165 -1275 -131 -1241
rect -165 -1343 -131 -1309
rect -165 -1411 -131 -1377
rect -165 -1479 -131 -1445
rect -165 -1547 -131 -1513
rect -165 -1615 -131 -1581
rect -165 -1683 -131 -1649
rect -165 -1751 -131 -1717
rect -165 -1819 -131 -1785
rect -165 -1887 -131 -1853
rect -165 -1955 -131 -1921
rect 131 1921 165 1955
rect 131 1853 165 1887
rect 131 1785 165 1819
rect 131 1717 165 1751
rect 131 1649 165 1683
rect 131 1581 165 1615
rect 131 1513 165 1547
rect 131 1445 165 1479
rect 131 1377 165 1411
rect 131 1309 165 1343
rect 131 1241 165 1275
rect 131 1173 165 1207
rect 131 1105 165 1139
rect 131 1037 165 1071
rect 131 969 165 1003
rect 131 901 165 935
rect 131 833 165 867
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect 131 -867 165 -833
rect 131 -935 165 -901
rect 131 -1003 165 -969
rect 131 -1071 165 -1037
rect 131 -1139 165 -1105
rect 131 -1207 165 -1173
rect 131 -1275 165 -1241
rect 131 -1343 165 -1309
rect 131 -1411 165 -1377
rect 131 -1479 165 -1445
rect 131 -1547 165 -1513
rect 131 -1615 165 -1581
rect 131 -1683 165 -1649
rect 131 -1751 165 -1717
rect 131 -1819 165 -1785
rect 131 -1887 165 -1853
rect 131 -1955 165 -1921
rect -51 -2062 -17 -2028
rect 17 -2062 51 -2028
<< xpolycontact >>
rect -35 1500 35 1932
rect -35 -1932 35 -1500
<< ppolyres >>
rect -35 -1500 35 1500
<< locali >>
rect -165 2028 -51 2062
rect -17 2028 17 2062
rect 51 2028 165 2062
rect -165 1955 -131 2028
rect 131 1955 165 2028
rect -165 1887 -131 1921
rect -165 1819 -131 1853
rect -165 1751 -131 1785
rect -165 1683 -131 1717
rect -165 1615 -131 1649
rect -165 1547 -131 1581
rect -165 1479 -131 1513
rect 131 1887 165 1921
rect 131 1819 165 1853
rect 131 1751 165 1785
rect 131 1683 165 1717
rect 131 1615 165 1649
rect 131 1547 165 1581
rect -165 1411 -131 1445
rect -165 1343 -131 1377
rect -165 1275 -131 1309
rect -165 1207 -131 1241
rect -165 1139 -131 1173
rect -165 1071 -131 1105
rect -165 1003 -131 1037
rect -165 935 -131 969
rect -165 867 -131 901
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect -165 -901 -131 -867
rect -165 -969 -131 -935
rect -165 -1037 -131 -1003
rect -165 -1105 -131 -1071
rect -165 -1173 -131 -1139
rect -165 -1241 -131 -1207
rect -165 -1309 -131 -1275
rect -165 -1377 -131 -1343
rect -165 -1445 -131 -1411
rect -165 -1513 -131 -1479
rect 131 1479 165 1513
rect 131 1411 165 1445
rect 131 1343 165 1377
rect 131 1275 165 1309
rect 131 1207 165 1241
rect 131 1139 165 1173
rect 131 1071 165 1105
rect 131 1003 165 1037
rect 131 935 165 969
rect 131 867 165 901
rect 131 799 165 833
rect 131 731 165 765
rect 131 663 165 697
rect 131 595 165 629
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -663
rect 131 -765 165 -731
rect 131 -833 165 -799
rect 131 -901 165 -867
rect 131 -969 165 -935
rect 131 -1037 165 -1003
rect 131 -1105 165 -1071
rect 131 -1173 165 -1139
rect 131 -1241 165 -1207
rect 131 -1309 165 -1275
rect 131 -1377 165 -1343
rect 131 -1445 165 -1411
rect -165 -1581 -131 -1547
rect -165 -1649 -131 -1615
rect -165 -1717 -131 -1683
rect -165 -1785 -131 -1751
rect -165 -1853 -131 -1819
rect -165 -1921 -131 -1887
rect 131 -1513 165 -1479
rect 131 -1581 165 -1547
rect 131 -1649 165 -1615
rect 131 -1717 165 -1683
rect 131 -1785 165 -1751
rect 131 -1853 165 -1819
rect 131 -1921 165 -1887
rect -165 -2028 -131 -1955
rect 131 -2028 165 -1955
rect -165 -2062 -51 -2028
rect -17 -2062 17 -2028
rect 51 -2062 165 -2028
<< viali >>
rect -17 1878 17 1912
rect -17 1806 17 1840
rect -17 1734 17 1768
rect -17 1662 17 1696
rect -17 1590 17 1624
rect -17 1518 17 1552
rect -17 -1553 17 -1519
rect -17 -1625 17 -1591
rect -17 -1697 17 -1663
rect -17 -1769 17 -1735
rect -17 -1841 17 -1807
rect -17 -1913 17 -1879
<< metal1 >>
rect -25 1912 25 1926
rect -25 1878 -17 1912
rect 17 1878 25 1912
rect -25 1840 25 1878
rect -25 1806 -17 1840
rect 17 1806 25 1840
rect -25 1768 25 1806
rect -25 1734 -17 1768
rect 17 1734 25 1768
rect -25 1696 25 1734
rect -25 1662 -17 1696
rect 17 1662 25 1696
rect -25 1624 25 1662
rect -25 1590 -17 1624
rect 17 1590 25 1624
rect -25 1552 25 1590
rect -25 1518 -17 1552
rect 17 1518 25 1552
rect -25 1505 25 1518
rect -25 -1519 25 -1505
rect -25 -1553 -17 -1519
rect 17 -1553 25 -1519
rect -25 -1591 25 -1553
rect -25 -1625 -17 -1591
rect 17 -1625 25 -1591
rect -25 -1663 25 -1625
rect -25 -1697 -17 -1663
rect 17 -1697 25 -1663
rect -25 -1735 25 -1697
rect -25 -1769 -17 -1735
rect 17 -1769 25 -1735
rect -25 -1807 25 -1769
rect -25 -1841 -17 -1807
rect 17 -1841 25 -1807
rect -25 -1879 25 -1841
rect -25 -1913 -17 -1879
rect 17 -1913 25 -1879
rect -25 -1926 25 -1913
<< properties >>
string FIXED_BBOX -148 -2045 148 2045
<< end >>
