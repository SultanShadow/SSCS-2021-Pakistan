magic
tech sky130A
magscale 1 2
timestamp 1635855079
<< error_p >>
rect -31 2072 31 2078
rect -31 2038 -17 2072
rect -31 2032 31 2038
rect -31 -2038 31 -2032
rect -31 -2072 -17 -2038
rect -31 -2078 31 -2072
<< pwell >>
rect -221 -2200 221 2200
<< nmoslvt >>
rect -35 -2000 35 2000
<< ndiff >>
rect -93 1955 -35 2000
rect -93 1921 -81 1955
rect -47 1921 -35 1955
rect -93 1887 -35 1921
rect -93 1853 -81 1887
rect -47 1853 -35 1887
rect -93 1819 -35 1853
rect -93 1785 -81 1819
rect -47 1785 -35 1819
rect -93 1751 -35 1785
rect -93 1717 -81 1751
rect -47 1717 -35 1751
rect -93 1683 -35 1717
rect -93 1649 -81 1683
rect -47 1649 -35 1683
rect -93 1615 -35 1649
rect -93 1581 -81 1615
rect -47 1581 -35 1615
rect -93 1547 -35 1581
rect -93 1513 -81 1547
rect -47 1513 -35 1547
rect -93 1479 -35 1513
rect -93 1445 -81 1479
rect -47 1445 -35 1479
rect -93 1411 -35 1445
rect -93 1377 -81 1411
rect -47 1377 -35 1411
rect -93 1343 -35 1377
rect -93 1309 -81 1343
rect -47 1309 -35 1343
rect -93 1275 -35 1309
rect -93 1241 -81 1275
rect -47 1241 -35 1275
rect -93 1207 -35 1241
rect -93 1173 -81 1207
rect -47 1173 -35 1207
rect -93 1139 -35 1173
rect -93 1105 -81 1139
rect -47 1105 -35 1139
rect -93 1071 -35 1105
rect -93 1037 -81 1071
rect -47 1037 -35 1071
rect -93 1003 -35 1037
rect -93 969 -81 1003
rect -47 969 -35 1003
rect -93 935 -35 969
rect -93 901 -81 935
rect -47 901 -35 935
rect -93 867 -35 901
rect -93 833 -81 867
rect -47 833 -35 867
rect -93 799 -35 833
rect -93 765 -81 799
rect -47 765 -35 799
rect -93 731 -35 765
rect -93 697 -81 731
rect -47 697 -35 731
rect -93 663 -35 697
rect -93 629 -81 663
rect -47 629 -35 663
rect -93 595 -35 629
rect -93 561 -81 595
rect -47 561 -35 595
rect -93 527 -35 561
rect -93 493 -81 527
rect -47 493 -35 527
rect -93 459 -35 493
rect -93 425 -81 459
rect -47 425 -35 459
rect -93 391 -35 425
rect -93 357 -81 391
rect -47 357 -35 391
rect -93 323 -35 357
rect -93 289 -81 323
rect -47 289 -35 323
rect -93 255 -35 289
rect -93 221 -81 255
rect -47 221 -35 255
rect -93 187 -35 221
rect -93 153 -81 187
rect -47 153 -35 187
rect -93 119 -35 153
rect -93 85 -81 119
rect -47 85 -35 119
rect -93 51 -35 85
rect -93 17 -81 51
rect -47 17 -35 51
rect -93 -17 -35 17
rect -93 -51 -81 -17
rect -47 -51 -35 -17
rect -93 -85 -35 -51
rect -93 -119 -81 -85
rect -47 -119 -35 -85
rect -93 -153 -35 -119
rect -93 -187 -81 -153
rect -47 -187 -35 -153
rect -93 -221 -35 -187
rect -93 -255 -81 -221
rect -47 -255 -35 -221
rect -93 -289 -35 -255
rect -93 -323 -81 -289
rect -47 -323 -35 -289
rect -93 -357 -35 -323
rect -93 -391 -81 -357
rect -47 -391 -35 -357
rect -93 -425 -35 -391
rect -93 -459 -81 -425
rect -47 -459 -35 -425
rect -93 -493 -35 -459
rect -93 -527 -81 -493
rect -47 -527 -35 -493
rect -93 -561 -35 -527
rect -93 -595 -81 -561
rect -47 -595 -35 -561
rect -93 -629 -35 -595
rect -93 -663 -81 -629
rect -47 -663 -35 -629
rect -93 -697 -35 -663
rect -93 -731 -81 -697
rect -47 -731 -35 -697
rect -93 -765 -35 -731
rect -93 -799 -81 -765
rect -47 -799 -35 -765
rect -93 -833 -35 -799
rect -93 -867 -81 -833
rect -47 -867 -35 -833
rect -93 -901 -35 -867
rect -93 -935 -81 -901
rect -47 -935 -35 -901
rect -93 -969 -35 -935
rect -93 -1003 -81 -969
rect -47 -1003 -35 -969
rect -93 -1037 -35 -1003
rect -93 -1071 -81 -1037
rect -47 -1071 -35 -1037
rect -93 -1105 -35 -1071
rect -93 -1139 -81 -1105
rect -47 -1139 -35 -1105
rect -93 -1173 -35 -1139
rect -93 -1207 -81 -1173
rect -47 -1207 -35 -1173
rect -93 -1241 -35 -1207
rect -93 -1275 -81 -1241
rect -47 -1275 -35 -1241
rect -93 -1309 -35 -1275
rect -93 -1343 -81 -1309
rect -47 -1343 -35 -1309
rect -93 -1377 -35 -1343
rect -93 -1411 -81 -1377
rect -47 -1411 -35 -1377
rect -93 -1445 -35 -1411
rect -93 -1479 -81 -1445
rect -47 -1479 -35 -1445
rect -93 -1513 -35 -1479
rect -93 -1547 -81 -1513
rect -47 -1547 -35 -1513
rect -93 -1581 -35 -1547
rect -93 -1615 -81 -1581
rect -47 -1615 -35 -1581
rect -93 -1649 -35 -1615
rect -93 -1683 -81 -1649
rect -47 -1683 -35 -1649
rect -93 -1717 -35 -1683
rect -93 -1751 -81 -1717
rect -47 -1751 -35 -1717
rect -93 -1785 -35 -1751
rect -93 -1819 -81 -1785
rect -47 -1819 -35 -1785
rect -93 -1853 -35 -1819
rect -93 -1887 -81 -1853
rect -47 -1887 -35 -1853
rect -93 -1921 -35 -1887
rect -93 -1955 -81 -1921
rect -47 -1955 -35 -1921
rect -93 -2000 -35 -1955
rect 35 1955 93 2000
rect 35 1921 47 1955
rect 81 1921 93 1955
rect 35 1887 93 1921
rect 35 1853 47 1887
rect 81 1853 93 1887
rect 35 1819 93 1853
rect 35 1785 47 1819
rect 81 1785 93 1819
rect 35 1751 93 1785
rect 35 1717 47 1751
rect 81 1717 93 1751
rect 35 1683 93 1717
rect 35 1649 47 1683
rect 81 1649 93 1683
rect 35 1615 93 1649
rect 35 1581 47 1615
rect 81 1581 93 1615
rect 35 1547 93 1581
rect 35 1513 47 1547
rect 81 1513 93 1547
rect 35 1479 93 1513
rect 35 1445 47 1479
rect 81 1445 93 1479
rect 35 1411 93 1445
rect 35 1377 47 1411
rect 81 1377 93 1411
rect 35 1343 93 1377
rect 35 1309 47 1343
rect 81 1309 93 1343
rect 35 1275 93 1309
rect 35 1241 47 1275
rect 81 1241 93 1275
rect 35 1207 93 1241
rect 35 1173 47 1207
rect 81 1173 93 1207
rect 35 1139 93 1173
rect 35 1105 47 1139
rect 81 1105 93 1139
rect 35 1071 93 1105
rect 35 1037 47 1071
rect 81 1037 93 1071
rect 35 1003 93 1037
rect 35 969 47 1003
rect 81 969 93 1003
rect 35 935 93 969
rect 35 901 47 935
rect 81 901 93 935
rect 35 867 93 901
rect 35 833 47 867
rect 81 833 93 867
rect 35 799 93 833
rect 35 765 47 799
rect 81 765 93 799
rect 35 731 93 765
rect 35 697 47 731
rect 81 697 93 731
rect 35 663 93 697
rect 35 629 47 663
rect 81 629 93 663
rect 35 595 93 629
rect 35 561 47 595
rect 81 561 93 595
rect 35 527 93 561
rect 35 493 47 527
rect 81 493 93 527
rect 35 459 93 493
rect 35 425 47 459
rect 81 425 93 459
rect 35 391 93 425
rect 35 357 47 391
rect 81 357 93 391
rect 35 323 93 357
rect 35 289 47 323
rect 81 289 93 323
rect 35 255 93 289
rect 35 221 47 255
rect 81 221 93 255
rect 35 187 93 221
rect 35 153 47 187
rect 81 153 93 187
rect 35 119 93 153
rect 35 85 47 119
rect 81 85 93 119
rect 35 51 93 85
rect 35 17 47 51
rect 81 17 93 51
rect 35 -17 93 17
rect 35 -51 47 -17
rect 81 -51 93 -17
rect 35 -85 93 -51
rect 35 -119 47 -85
rect 81 -119 93 -85
rect 35 -153 93 -119
rect 35 -187 47 -153
rect 81 -187 93 -153
rect 35 -221 93 -187
rect 35 -255 47 -221
rect 81 -255 93 -221
rect 35 -289 93 -255
rect 35 -323 47 -289
rect 81 -323 93 -289
rect 35 -357 93 -323
rect 35 -391 47 -357
rect 81 -391 93 -357
rect 35 -425 93 -391
rect 35 -459 47 -425
rect 81 -459 93 -425
rect 35 -493 93 -459
rect 35 -527 47 -493
rect 81 -527 93 -493
rect 35 -561 93 -527
rect 35 -595 47 -561
rect 81 -595 93 -561
rect 35 -629 93 -595
rect 35 -663 47 -629
rect 81 -663 93 -629
rect 35 -697 93 -663
rect 35 -731 47 -697
rect 81 -731 93 -697
rect 35 -765 93 -731
rect 35 -799 47 -765
rect 81 -799 93 -765
rect 35 -833 93 -799
rect 35 -867 47 -833
rect 81 -867 93 -833
rect 35 -901 93 -867
rect 35 -935 47 -901
rect 81 -935 93 -901
rect 35 -969 93 -935
rect 35 -1003 47 -969
rect 81 -1003 93 -969
rect 35 -1037 93 -1003
rect 35 -1071 47 -1037
rect 81 -1071 93 -1037
rect 35 -1105 93 -1071
rect 35 -1139 47 -1105
rect 81 -1139 93 -1105
rect 35 -1173 93 -1139
rect 35 -1207 47 -1173
rect 81 -1207 93 -1173
rect 35 -1241 93 -1207
rect 35 -1275 47 -1241
rect 81 -1275 93 -1241
rect 35 -1309 93 -1275
rect 35 -1343 47 -1309
rect 81 -1343 93 -1309
rect 35 -1377 93 -1343
rect 35 -1411 47 -1377
rect 81 -1411 93 -1377
rect 35 -1445 93 -1411
rect 35 -1479 47 -1445
rect 81 -1479 93 -1445
rect 35 -1513 93 -1479
rect 35 -1547 47 -1513
rect 81 -1547 93 -1513
rect 35 -1581 93 -1547
rect 35 -1615 47 -1581
rect 81 -1615 93 -1581
rect 35 -1649 93 -1615
rect 35 -1683 47 -1649
rect 81 -1683 93 -1649
rect 35 -1717 93 -1683
rect 35 -1751 47 -1717
rect 81 -1751 93 -1717
rect 35 -1785 93 -1751
rect 35 -1819 47 -1785
rect 81 -1819 93 -1785
rect 35 -1853 93 -1819
rect 35 -1887 47 -1853
rect 81 -1887 93 -1853
rect 35 -1921 93 -1887
rect 35 -1955 47 -1921
rect 81 -1955 93 -1921
rect 35 -2000 93 -1955
<< ndiffc >>
rect -81 1921 -47 1955
rect -81 1853 -47 1887
rect -81 1785 -47 1819
rect -81 1717 -47 1751
rect -81 1649 -47 1683
rect -81 1581 -47 1615
rect -81 1513 -47 1547
rect -81 1445 -47 1479
rect -81 1377 -47 1411
rect -81 1309 -47 1343
rect -81 1241 -47 1275
rect -81 1173 -47 1207
rect -81 1105 -47 1139
rect -81 1037 -47 1071
rect -81 969 -47 1003
rect -81 901 -47 935
rect -81 833 -47 867
rect -81 765 -47 799
rect -81 697 -47 731
rect -81 629 -47 663
rect -81 561 -47 595
rect -81 493 -47 527
rect -81 425 -47 459
rect -81 357 -47 391
rect -81 289 -47 323
rect -81 221 -47 255
rect -81 153 -47 187
rect -81 85 -47 119
rect -81 17 -47 51
rect -81 -51 -47 -17
rect -81 -119 -47 -85
rect -81 -187 -47 -153
rect -81 -255 -47 -221
rect -81 -323 -47 -289
rect -81 -391 -47 -357
rect -81 -459 -47 -425
rect -81 -527 -47 -493
rect -81 -595 -47 -561
rect -81 -663 -47 -629
rect -81 -731 -47 -697
rect -81 -799 -47 -765
rect -81 -867 -47 -833
rect -81 -935 -47 -901
rect -81 -1003 -47 -969
rect -81 -1071 -47 -1037
rect -81 -1139 -47 -1105
rect -81 -1207 -47 -1173
rect -81 -1275 -47 -1241
rect -81 -1343 -47 -1309
rect -81 -1411 -47 -1377
rect -81 -1479 -47 -1445
rect -81 -1547 -47 -1513
rect -81 -1615 -47 -1581
rect -81 -1683 -47 -1649
rect -81 -1751 -47 -1717
rect -81 -1819 -47 -1785
rect -81 -1887 -47 -1853
rect -81 -1955 -47 -1921
rect 47 1921 81 1955
rect 47 1853 81 1887
rect 47 1785 81 1819
rect 47 1717 81 1751
rect 47 1649 81 1683
rect 47 1581 81 1615
rect 47 1513 81 1547
rect 47 1445 81 1479
rect 47 1377 81 1411
rect 47 1309 81 1343
rect 47 1241 81 1275
rect 47 1173 81 1207
rect 47 1105 81 1139
rect 47 1037 81 1071
rect 47 969 81 1003
rect 47 901 81 935
rect 47 833 81 867
rect 47 765 81 799
rect 47 697 81 731
rect 47 629 81 663
rect 47 561 81 595
rect 47 493 81 527
rect 47 425 81 459
rect 47 357 81 391
rect 47 289 81 323
rect 47 221 81 255
rect 47 153 81 187
rect 47 85 81 119
rect 47 17 81 51
rect 47 -51 81 -17
rect 47 -119 81 -85
rect 47 -187 81 -153
rect 47 -255 81 -221
rect 47 -323 81 -289
rect 47 -391 81 -357
rect 47 -459 81 -425
rect 47 -527 81 -493
rect 47 -595 81 -561
rect 47 -663 81 -629
rect 47 -731 81 -697
rect 47 -799 81 -765
rect 47 -867 81 -833
rect 47 -935 81 -901
rect 47 -1003 81 -969
rect 47 -1071 81 -1037
rect 47 -1139 81 -1105
rect 47 -1207 81 -1173
rect 47 -1275 81 -1241
rect 47 -1343 81 -1309
rect 47 -1411 81 -1377
rect 47 -1479 81 -1445
rect 47 -1547 81 -1513
rect 47 -1615 81 -1581
rect 47 -1683 81 -1649
rect 47 -1751 81 -1717
rect 47 -1819 81 -1785
rect 47 -1887 81 -1853
rect 47 -1955 81 -1921
<< psubdiff >>
rect -195 2140 -85 2174
rect -51 2140 -17 2174
rect 17 2140 51 2174
rect 85 2140 195 2174
rect -195 2057 -161 2140
rect -195 1989 -161 2023
rect 161 2057 195 2140
rect -195 1921 -161 1955
rect -195 1853 -161 1887
rect -195 1785 -161 1819
rect -195 1717 -161 1751
rect -195 1649 -161 1683
rect -195 1581 -161 1615
rect -195 1513 -161 1547
rect -195 1445 -161 1479
rect -195 1377 -161 1411
rect -195 1309 -161 1343
rect -195 1241 -161 1275
rect -195 1173 -161 1207
rect -195 1105 -161 1139
rect -195 1037 -161 1071
rect -195 969 -161 1003
rect -195 901 -161 935
rect -195 833 -161 867
rect -195 765 -161 799
rect -195 697 -161 731
rect -195 629 -161 663
rect -195 561 -161 595
rect -195 493 -161 527
rect -195 425 -161 459
rect -195 357 -161 391
rect -195 289 -161 323
rect -195 221 -161 255
rect -195 153 -161 187
rect -195 85 -161 119
rect -195 17 -161 51
rect -195 -51 -161 -17
rect -195 -119 -161 -85
rect -195 -187 -161 -153
rect -195 -255 -161 -221
rect -195 -323 -161 -289
rect -195 -391 -161 -357
rect -195 -459 -161 -425
rect -195 -527 -161 -493
rect -195 -595 -161 -561
rect -195 -663 -161 -629
rect -195 -731 -161 -697
rect -195 -799 -161 -765
rect -195 -867 -161 -833
rect -195 -935 -161 -901
rect -195 -1003 -161 -969
rect -195 -1071 -161 -1037
rect -195 -1139 -161 -1105
rect -195 -1207 -161 -1173
rect -195 -1275 -161 -1241
rect -195 -1343 -161 -1309
rect -195 -1411 -161 -1377
rect -195 -1479 -161 -1445
rect -195 -1547 -161 -1513
rect -195 -1615 -161 -1581
rect -195 -1683 -161 -1649
rect -195 -1751 -161 -1717
rect -195 -1819 -161 -1785
rect -195 -1887 -161 -1853
rect -195 -1955 -161 -1921
rect -195 -2023 -161 -1989
rect 161 1989 195 2023
rect 161 1921 195 1955
rect 161 1853 195 1887
rect 161 1785 195 1819
rect 161 1717 195 1751
rect 161 1649 195 1683
rect 161 1581 195 1615
rect 161 1513 195 1547
rect 161 1445 195 1479
rect 161 1377 195 1411
rect 161 1309 195 1343
rect 161 1241 195 1275
rect 161 1173 195 1207
rect 161 1105 195 1139
rect 161 1037 195 1071
rect 161 969 195 1003
rect 161 901 195 935
rect 161 833 195 867
rect 161 765 195 799
rect 161 697 195 731
rect 161 629 195 663
rect 161 561 195 595
rect 161 493 195 527
rect 161 425 195 459
rect 161 357 195 391
rect 161 289 195 323
rect 161 221 195 255
rect 161 153 195 187
rect 161 85 195 119
rect 161 17 195 51
rect 161 -51 195 -17
rect 161 -119 195 -85
rect 161 -187 195 -153
rect 161 -255 195 -221
rect 161 -323 195 -289
rect 161 -391 195 -357
rect 161 -459 195 -425
rect 161 -527 195 -493
rect 161 -595 195 -561
rect 161 -663 195 -629
rect 161 -731 195 -697
rect 161 -799 195 -765
rect 161 -867 195 -833
rect 161 -935 195 -901
rect 161 -1003 195 -969
rect 161 -1071 195 -1037
rect 161 -1139 195 -1105
rect 161 -1207 195 -1173
rect 161 -1275 195 -1241
rect 161 -1343 195 -1309
rect 161 -1411 195 -1377
rect 161 -1479 195 -1445
rect 161 -1547 195 -1513
rect 161 -1615 195 -1581
rect 161 -1683 195 -1649
rect 161 -1751 195 -1717
rect 161 -1819 195 -1785
rect 161 -1887 195 -1853
rect 161 -1955 195 -1921
rect -195 -2140 -161 -2057
rect 161 -2023 195 -1989
rect 161 -2140 195 -2057
rect -195 -2174 -85 -2140
rect -51 -2174 -17 -2140
rect 17 -2174 51 -2140
rect 85 -2174 195 -2140
<< psubdiffcont >>
rect -85 2140 -51 2174
rect -17 2140 17 2174
rect 51 2140 85 2174
rect -195 2023 -161 2057
rect 161 2023 195 2057
rect -195 1955 -161 1989
rect -195 1887 -161 1921
rect -195 1819 -161 1853
rect -195 1751 -161 1785
rect -195 1683 -161 1717
rect -195 1615 -161 1649
rect -195 1547 -161 1581
rect -195 1479 -161 1513
rect -195 1411 -161 1445
rect -195 1343 -161 1377
rect -195 1275 -161 1309
rect -195 1207 -161 1241
rect -195 1139 -161 1173
rect -195 1071 -161 1105
rect -195 1003 -161 1037
rect -195 935 -161 969
rect -195 867 -161 901
rect -195 799 -161 833
rect -195 731 -161 765
rect -195 663 -161 697
rect -195 595 -161 629
rect -195 527 -161 561
rect -195 459 -161 493
rect -195 391 -161 425
rect -195 323 -161 357
rect -195 255 -161 289
rect -195 187 -161 221
rect -195 119 -161 153
rect -195 51 -161 85
rect -195 -17 -161 17
rect -195 -85 -161 -51
rect -195 -153 -161 -119
rect -195 -221 -161 -187
rect -195 -289 -161 -255
rect -195 -357 -161 -323
rect -195 -425 -161 -391
rect -195 -493 -161 -459
rect -195 -561 -161 -527
rect -195 -629 -161 -595
rect -195 -697 -161 -663
rect -195 -765 -161 -731
rect -195 -833 -161 -799
rect -195 -901 -161 -867
rect -195 -969 -161 -935
rect -195 -1037 -161 -1003
rect -195 -1105 -161 -1071
rect -195 -1173 -161 -1139
rect -195 -1241 -161 -1207
rect -195 -1309 -161 -1275
rect -195 -1377 -161 -1343
rect -195 -1445 -161 -1411
rect -195 -1513 -161 -1479
rect -195 -1581 -161 -1547
rect -195 -1649 -161 -1615
rect -195 -1717 -161 -1683
rect -195 -1785 -161 -1751
rect -195 -1853 -161 -1819
rect -195 -1921 -161 -1887
rect -195 -1989 -161 -1955
rect 161 1955 195 1989
rect 161 1887 195 1921
rect 161 1819 195 1853
rect 161 1751 195 1785
rect 161 1683 195 1717
rect 161 1615 195 1649
rect 161 1547 195 1581
rect 161 1479 195 1513
rect 161 1411 195 1445
rect 161 1343 195 1377
rect 161 1275 195 1309
rect 161 1207 195 1241
rect 161 1139 195 1173
rect 161 1071 195 1105
rect 161 1003 195 1037
rect 161 935 195 969
rect 161 867 195 901
rect 161 799 195 833
rect 161 731 195 765
rect 161 663 195 697
rect 161 595 195 629
rect 161 527 195 561
rect 161 459 195 493
rect 161 391 195 425
rect 161 323 195 357
rect 161 255 195 289
rect 161 187 195 221
rect 161 119 195 153
rect 161 51 195 85
rect 161 -17 195 17
rect 161 -85 195 -51
rect 161 -153 195 -119
rect 161 -221 195 -187
rect 161 -289 195 -255
rect 161 -357 195 -323
rect 161 -425 195 -391
rect 161 -493 195 -459
rect 161 -561 195 -527
rect 161 -629 195 -595
rect 161 -697 195 -663
rect 161 -765 195 -731
rect 161 -833 195 -799
rect 161 -901 195 -867
rect 161 -969 195 -935
rect 161 -1037 195 -1003
rect 161 -1105 195 -1071
rect 161 -1173 195 -1139
rect 161 -1241 195 -1207
rect 161 -1309 195 -1275
rect 161 -1377 195 -1343
rect 161 -1445 195 -1411
rect 161 -1513 195 -1479
rect 161 -1581 195 -1547
rect 161 -1649 195 -1615
rect 161 -1717 195 -1683
rect 161 -1785 195 -1751
rect 161 -1853 195 -1819
rect 161 -1921 195 -1887
rect 161 -1989 195 -1955
rect -195 -2057 -161 -2023
rect 161 -2057 195 -2023
rect -85 -2174 -51 -2140
rect -17 -2174 17 -2140
rect 51 -2174 85 -2140
<< poly >>
rect -35 2072 35 2088
rect -35 2038 -17 2072
rect 17 2038 35 2072
rect -35 2000 35 2038
rect -35 -2038 35 -2000
rect -35 -2072 -17 -2038
rect 17 -2072 35 -2038
rect -35 -2088 35 -2072
<< polycont >>
rect -17 2038 17 2072
rect -17 -2072 17 -2038
<< locali >>
rect -195 2140 -85 2174
rect -51 2140 -17 2174
rect 17 2140 51 2174
rect 85 2140 195 2174
rect -195 2057 -161 2140
rect -35 2038 -17 2072
rect 17 2038 35 2072
rect 161 2057 195 2140
rect -195 1989 -161 2023
rect -195 1921 -161 1955
rect -195 1853 -161 1887
rect -195 1785 -161 1819
rect -195 1717 -161 1751
rect -195 1649 -161 1683
rect -195 1581 -161 1615
rect -195 1513 -161 1547
rect -195 1445 -161 1479
rect -195 1377 -161 1411
rect -195 1309 -161 1343
rect -195 1241 -161 1275
rect -195 1173 -161 1207
rect -195 1105 -161 1139
rect -195 1037 -161 1071
rect -195 969 -161 1003
rect -195 901 -161 935
rect -195 833 -161 867
rect -195 765 -161 799
rect -195 697 -161 731
rect -195 629 -161 663
rect -195 561 -161 595
rect -195 493 -161 527
rect -195 425 -161 459
rect -195 357 -161 391
rect -195 289 -161 323
rect -195 221 -161 255
rect -195 153 -161 187
rect -195 85 -161 119
rect -195 17 -161 51
rect -195 -51 -161 -17
rect -195 -119 -161 -85
rect -195 -187 -161 -153
rect -195 -255 -161 -221
rect -195 -323 -161 -289
rect -195 -391 -161 -357
rect -195 -459 -161 -425
rect -195 -527 -161 -493
rect -195 -595 -161 -561
rect -195 -663 -161 -629
rect -195 -731 -161 -697
rect -195 -799 -161 -765
rect -195 -867 -161 -833
rect -195 -935 -161 -901
rect -195 -1003 -161 -969
rect -195 -1071 -161 -1037
rect -195 -1139 -161 -1105
rect -195 -1207 -161 -1173
rect -195 -1275 -161 -1241
rect -195 -1343 -161 -1309
rect -195 -1411 -161 -1377
rect -195 -1479 -161 -1445
rect -195 -1547 -161 -1513
rect -195 -1615 -161 -1581
rect -195 -1683 -161 -1649
rect -195 -1751 -161 -1717
rect -195 -1819 -161 -1785
rect -195 -1887 -161 -1853
rect -195 -1955 -161 -1921
rect -195 -2023 -161 -1989
rect -81 1961 -47 2004
rect -81 1889 -47 1921
rect -81 1819 -47 1853
rect -81 1751 -47 1783
rect -81 1683 -47 1711
rect -81 1615 -47 1639
rect -81 1547 -47 1567
rect -81 1479 -47 1495
rect -81 1411 -47 1423
rect -81 1343 -47 1351
rect -81 1275 -47 1279
rect -81 1169 -47 1173
rect -81 1097 -47 1105
rect -81 1025 -47 1037
rect -81 953 -47 969
rect -81 881 -47 901
rect -81 809 -47 833
rect -81 737 -47 765
rect -81 665 -47 697
rect -81 595 -47 629
rect -81 527 -47 559
rect -81 459 -47 487
rect -81 391 -47 415
rect -81 323 -47 343
rect -81 255 -47 271
rect -81 187 -47 199
rect -81 119 -47 127
rect -81 51 -47 55
rect -81 -55 -47 -51
rect -81 -127 -47 -119
rect -81 -199 -47 -187
rect -81 -271 -47 -255
rect -81 -343 -47 -323
rect -81 -415 -47 -391
rect -81 -487 -47 -459
rect -81 -559 -47 -527
rect -81 -629 -47 -595
rect -81 -697 -47 -665
rect -81 -765 -47 -737
rect -81 -833 -47 -809
rect -81 -901 -47 -881
rect -81 -969 -47 -953
rect -81 -1037 -47 -1025
rect -81 -1105 -47 -1097
rect -81 -1173 -47 -1169
rect -81 -1279 -47 -1275
rect -81 -1351 -47 -1343
rect -81 -1423 -47 -1411
rect -81 -1495 -47 -1479
rect -81 -1567 -47 -1547
rect -81 -1639 -47 -1615
rect -81 -1711 -47 -1683
rect -81 -1783 -47 -1751
rect -81 -1853 -47 -1819
rect -81 -1921 -47 -1889
rect -81 -2004 -47 -1961
rect 47 1961 81 2004
rect 47 1889 81 1921
rect 47 1819 81 1853
rect 47 1751 81 1783
rect 47 1683 81 1711
rect 47 1615 81 1639
rect 47 1547 81 1567
rect 47 1479 81 1495
rect 47 1411 81 1423
rect 47 1343 81 1351
rect 47 1275 81 1279
rect 47 1169 81 1173
rect 47 1097 81 1105
rect 47 1025 81 1037
rect 47 953 81 969
rect 47 881 81 901
rect 47 809 81 833
rect 47 737 81 765
rect 47 665 81 697
rect 47 595 81 629
rect 47 527 81 559
rect 47 459 81 487
rect 47 391 81 415
rect 47 323 81 343
rect 47 255 81 271
rect 47 187 81 199
rect 47 119 81 127
rect 47 51 81 55
rect 47 -55 81 -51
rect 47 -127 81 -119
rect 47 -199 81 -187
rect 47 -271 81 -255
rect 47 -343 81 -323
rect 47 -415 81 -391
rect 47 -487 81 -459
rect 47 -559 81 -527
rect 47 -629 81 -595
rect 47 -697 81 -665
rect 47 -765 81 -737
rect 47 -833 81 -809
rect 47 -901 81 -881
rect 47 -969 81 -953
rect 47 -1037 81 -1025
rect 47 -1105 81 -1097
rect 47 -1173 81 -1169
rect 47 -1279 81 -1275
rect 47 -1351 81 -1343
rect 47 -1423 81 -1411
rect 47 -1495 81 -1479
rect 47 -1567 81 -1547
rect 47 -1639 81 -1615
rect 47 -1711 81 -1683
rect 47 -1783 81 -1751
rect 47 -1853 81 -1819
rect 47 -1921 81 -1889
rect 47 -2004 81 -1961
rect 161 1989 195 2023
rect 161 1921 195 1955
rect 161 1853 195 1887
rect 161 1785 195 1819
rect 161 1717 195 1751
rect 161 1649 195 1683
rect 161 1581 195 1615
rect 161 1513 195 1547
rect 161 1445 195 1479
rect 161 1377 195 1411
rect 161 1309 195 1343
rect 161 1241 195 1275
rect 161 1173 195 1207
rect 161 1105 195 1139
rect 161 1037 195 1071
rect 161 969 195 1003
rect 161 901 195 935
rect 161 833 195 867
rect 161 765 195 799
rect 161 697 195 731
rect 161 629 195 663
rect 161 561 195 595
rect 161 493 195 527
rect 161 425 195 459
rect 161 357 195 391
rect 161 289 195 323
rect 161 221 195 255
rect 161 153 195 187
rect 161 85 195 119
rect 161 17 195 51
rect 161 -51 195 -17
rect 161 -119 195 -85
rect 161 -187 195 -153
rect 161 -255 195 -221
rect 161 -323 195 -289
rect 161 -391 195 -357
rect 161 -459 195 -425
rect 161 -527 195 -493
rect 161 -595 195 -561
rect 161 -663 195 -629
rect 161 -731 195 -697
rect 161 -799 195 -765
rect 161 -867 195 -833
rect 161 -935 195 -901
rect 161 -1003 195 -969
rect 161 -1071 195 -1037
rect 161 -1139 195 -1105
rect 161 -1207 195 -1173
rect 161 -1275 195 -1241
rect 161 -1343 195 -1309
rect 161 -1411 195 -1377
rect 161 -1479 195 -1445
rect 161 -1547 195 -1513
rect 161 -1615 195 -1581
rect 161 -1683 195 -1649
rect 161 -1751 195 -1717
rect 161 -1819 195 -1785
rect 161 -1887 195 -1853
rect 161 -1955 195 -1921
rect 161 -2023 195 -1989
rect -195 -2140 -161 -2057
rect -35 -2072 -17 -2038
rect 17 -2072 35 -2038
rect 161 -2140 195 -2057
rect -195 -2174 -85 -2140
rect -51 -2174 -17 -2140
rect 17 -2174 51 -2140
rect 85 -2174 195 -2140
<< viali >>
rect -17 2038 17 2072
rect -81 1955 -47 1961
rect -81 1927 -47 1955
rect -81 1887 -47 1889
rect -81 1855 -47 1887
rect -81 1785 -47 1817
rect -81 1783 -47 1785
rect -81 1717 -47 1745
rect -81 1711 -47 1717
rect -81 1649 -47 1673
rect -81 1639 -47 1649
rect -81 1581 -47 1601
rect -81 1567 -47 1581
rect -81 1513 -47 1529
rect -81 1495 -47 1513
rect -81 1445 -47 1457
rect -81 1423 -47 1445
rect -81 1377 -47 1385
rect -81 1351 -47 1377
rect -81 1309 -47 1313
rect -81 1279 -47 1309
rect -81 1207 -47 1241
rect -81 1139 -47 1169
rect -81 1135 -47 1139
rect -81 1071 -47 1097
rect -81 1063 -47 1071
rect -81 1003 -47 1025
rect -81 991 -47 1003
rect -81 935 -47 953
rect -81 919 -47 935
rect -81 867 -47 881
rect -81 847 -47 867
rect -81 799 -47 809
rect -81 775 -47 799
rect -81 731 -47 737
rect -81 703 -47 731
rect -81 663 -47 665
rect -81 631 -47 663
rect -81 561 -47 593
rect -81 559 -47 561
rect -81 493 -47 521
rect -81 487 -47 493
rect -81 425 -47 449
rect -81 415 -47 425
rect -81 357 -47 377
rect -81 343 -47 357
rect -81 289 -47 305
rect -81 271 -47 289
rect -81 221 -47 233
rect -81 199 -47 221
rect -81 153 -47 161
rect -81 127 -47 153
rect -81 85 -47 89
rect -81 55 -47 85
rect -81 -17 -47 17
rect -81 -85 -47 -55
rect -81 -89 -47 -85
rect -81 -153 -47 -127
rect -81 -161 -47 -153
rect -81 -221 -47 -199
rect -81 -233 -47 -221
rect -81 -289 -47 -271
rect -81 -305 -47 -289
rect -81 -357 -47 -343
rect -81 -377 -47 -357
rect -81 -425 -47 -415
rect -81 -449 -47 -425
rect -81 -493 -47 -487
rect -81 -521 -47 -493
rect -81 -561 -47 -559
rect -81 -593 -47 -561
rect -81 -663 -47 -631
rect -81 -665 -47 -663
rect -81 -731 -47 -703
rect -81 -737 -47 -731
rect -81 -799 -47 -775
rect -81 -809 -47 -799
rect -81 -867 -47 -847
rect -81 -881 -47 -867
rect -81 -935 -47 -919
rect -81 -953 -47 -935
rect -81 -1003 -47 -991
rect -81 -1025 -47 -1003
rect -81 -1071 -47 -1063
rect -81 -1097 -47 -1071
rect -81 -1139 -47 -1135
rect -81 -1169 -47 -1139
rect -81 -1241 -47 -1207
rect -81 -1309 -47 -1279
rect -81 -1313 -47 -1309
rect -81 -1377 -47 -1351
rect -81 -1385 -47 -1377
rect -81 -1445 -47 -1423
rect -81 -1457 -47 -1445
rect -81 -1513 -47 -1495
rect -81 -1529 -47 -1513
rect -81 -1581 -47 -1567
rect -81 -1601 -47 -1581
rect -81 -1649 -47 -1639
rect -81 -1673 -47 -1649
rect -81 -1717 -47 -1711
rect -81 -1745 -47 -1717
rect -81 -1785 -47 -1783
rect -81 -1817 -47 -1785
rect -81 -1887 -47 -1855
rect -81 -1889 -47 -1887
rect -81 -1955 -47 -1927
rect -81 -1961 -47 -1955
rect 47 1955 81 1961
rect 47 1927 81 1955
rect 47 1887 81 1889
rect 47 1855 81 1887
rect 47 1785 81 1817
rect 47 1783 81 1785
rect 47 1717 81 1745
rect 47 1711 81 1717
rect 47 1649 81 1673
rect 47 1639 81 1649
rect 47 1581 81 1601
rect 47 1567 81 1581
rect 47 1513 81 1529
rect 47 1495 81 1513
rect 47 1445 81 1457
rect 47 1423 81 1445
rect 47 1377 81 1385
rect 47 1351 81 1377
rect 47 1309 81 1313
rect 47 1279 81 1309
rect 47 1207 81 1241
rect 47 1139 81 1169
rect 47 1135 81 1139
rect 47 1071 81 1097
rect 47 1063 81 1071
rect 47 1003 81 1025
rect 47 991 81 1003
rect 47 935 81 953
rect 47 919 81 935
rect 47 867 81 881
rect 47 847 81 867
rect 47 799 81 809
rect 47 775 81 799
rect 47 731 81 737
rect 47 703 81 731
rect 47 663 81 665
rect 47 631 81 663
rect 47 561 81 593
rect 47 559 81 561
rect 47 493 81 521
rect 47 487 81 493
rect 47 425 81 449
rect 47 415 81 425
rect 47 357 81 377
rect 47 343 81 357
rect 47 289 81 305
rect 47 271 81 289
rect 47 221 81 233
rect 47 199 81 221
rect 47 153 81 161
rect 47 127 81 153
rect 47 85 81 89
rect 47 55 81 85
rect 47 -17 81 17
rect 47 -85 81 -55
rect 47 -89 81 -85
rect 47 -153 81 -127
rect 47 -161 81 -153
rect 47 -221 81 -199
rect 47 -233 81 -221
rect 47 -289 81 -271
rect 47 -305 81 -289
rect 47 -357 81 -343
rect 47 -377 81 -357
rect 47 -425 81 -415
rect 47 -449 81 -425
rect 47 -493 81 -487
rect 47 -521 81 -493
rect 47 -561 81 -559
rect 47 -593 81 -561
rect 47 -663 81 -631
rect 47 -665 81 -663
rect 47 -731 81 -703
rect 47 -737 81 -731
rect 47 -799 81 -775
rect 47 -809 81 -799
rect 47 -867 81 -847
rect 47 -881 81 -867
rect 47 -935 81 -919
rect 47 -953 81 -935
rect 47 -1003 81 -991
rect 47 -1025 81 -1003
rect 47 -1071 81 -1063
rect 47 -1097 81 -1071
rect 47 -1139 81 -1135
rect 47 -1169 81 -1139
rect 47 -1241 81 -1207
rect 47 -1309 81 -1279
rect 47 -1313 81 -1309
rect 47 -1377 81 -1351
rect 47 -1385 81 -1377
rect 47 -1445 81 -1423
rect 47 -1457 81 -1445
rect 47 -1513 81 -1495
rect 47 -1529 81 -1513
rect 47 -1581 81 -1567
rect 47 -1601 81 -1581
rect 47 -1649 81 -1639
rect 47 -1673 81 -1649
rect 47 -1717 81 -1711
rect 47 -1745 81 -1717
rect 47 -1785 81 -1783
rect 47 -1817 81 -1785
rect 47 -1887 81 -1855
rect 47 -1889 81 -1887
rect 47 -1955 81 -1927
rect 47 -1961 81 -1955
rect -17 -2072 17 -2038
<< metal1 >>
rect -31 2072 31 2078
rect -31 2038 -17 2072
rect 17 2038 31 2072
rect -31 2032 31 2038
rect -87 1961 -41 2000
rect -87 1927 -81 1961
rect -47 1927 -41 1961
rect -87 1889 -41 1927
rect -87 1855 -81 1889
rect -47 1855 -41 1889
rect -87 1817 -41 1855
rect -87 1783 -81 1817
rect -47 1783 -41 1817
rect -87 1745 -41 1783
rect -87 1711 -81 1745
rect -47 1711 -41 1745
rect -87 1673 -41 1711
rect -87 1639 -81 1673
rect -47 1639 -41 1673
rect -87 1601 -41 1639
rect -87 1567 -81 1601
rect -47 1567 -41 1601
rect -87 1529 -41 1567
rect -87 1495 -81 1529
rect -47 1495 -41 1529
rect -87 1457 -41 1495
rect -87 1423 -81 1457
rect -47 1423 -41 1457
rect -87 1385 -41 1423
rect -87 1351 -81 1385
rect -47 1351 -41 1385
rect -87 1313 -41 1351
rect -87 1279 -81 1313
rect -47 1279 -41 1313
rect -87 1241 -41 1279
rect -87 1207 -81 1241
rect -47 1207 -41 1241
rect -87 1169 -41 1207
rect -87 1135 -81 1169
rect -47 1135 -41 1169
rect -87 1097 -41 1135
rect -87 1063 -81 1097
rect -47 1063 -41 1097
rect -87 1025 -41 1063
rect -87 991 -81 1025
rect -47 991 -41 1025
rect -87 953 -41 991
rect -87 919 -81 953
rect -47 919 -41 953
rect -87 881 -41 919
rect -87 847 -81 881
rect -47 847 -41 881
rect -87 809 -41 847
rect -87 775 -81 809
rect -47 775 -41 809
rect -87 737 -41 775
rect -87 703 -81 737
rect -47 703 -41 737
rect -87 665 -41 703
rect -87 631 -81 665
rect -47 631 -41 665
rect -87 593 -41 631
rect -87 559 -81 593
rect -47 559 -41 593
rect -87 521 -41 559
rect -87 487 -81 521
rect -47 487 -41 521
rect -87 449 -41 487
rect -87 415 -81 449
rect -47 415 -41 449
rect -87 377 -41 415
rect -87 343 -81 377
rect -47 343 -41 377
rect -87 305 -41 343
rect -87 271 -81 305
rect -47 271 -41 305
rect -87 233 -41 271
rect -87 199 -81 233
rect -47 199 -41 233
rect -87 161 -41 199
rect -87 127 -81 161
rect -47 127 -41 161
rect -87 89 -41 127
rect -87 55 -81 89
rect -47 55 -41 89
rect -87 17 -41 55
rect -87 -17 -81 17
rect -47 -17 -41 17
rect -87 -55 -41 -17
rect -87 -89 -81 -55
rect -47 -89 -41 -55
rect -87 -127 -41 -89
rect -87 -161 -81 -127
rect -47 -161 -41 -127
rect -87 -199 -41 -161
rect -87 -233 -81 -199
rect -47 -233 -41 -199
rect -87 -271 -41 -233
rect -87 -305 -81 -271
rect -47 -305 -41 -271
rect -87 -343 -41 -305
rect -87 -377 -81 -343
rect -47 -377 -41 -343
rect -87 -415 -41 -377
rect -87 -449 -81 -415
rect -47 -449 -41 -415
rect -87 -487 -41 -449
rect -87 -521 -81 -487
rect -47 -521 -41 -487
rect -87 -559 -41 -521
rect -87 -593 -81 -559
rect -47 -593 -41 -559
rect -87 -631 -41 -593
rect -87 -665 -81 -631
rect -47 -665 -41 -631
rect -87 -703 -41 -665
rect -87 -737 -81 -703
rect -47 -737 -41 -703
rect -87 -775 -41 -737
rect -87 -809 -81 -775
rect -47 -809 -41 -775
rect -87 -847 -41 -809
rect -87 -881 -81 -847
rect -47 -881 -41 -847
rect -87 -919 -41 -881
rect -87 -953 -81 -919
rect -47 -953 -41 -919
rect -87 -991 -41 -953
rect -87 -1025 -81 -991
rect -47 -1025 -41 -991
rect -87 -1063 -41 -1025
rect -87 -1097 -81 -1063
rect -47 -1097 -41 -1063
rect -87 -1135 -41 -1097
rect -87 -1169 -81 -1135
rect -47 -1169 -41 -1135
rect -87 -1207 -41 -1169
rect -87 -1241 -81 -1207
rect -47 -1241 -41 -1207
rect -87 -1279 -41 -1241
rect -87 -1313 -81 -1279
rect -47 -1313 -41 -1279
rect -87 -1351 -41 -1313
rect -87 -1385 -81 -1351
rect -47 -1385 -41 -1351
rect -87 -1423 -41 -1385
rect -87 -1457 -81 -1423
rect -47 -1457 -41 -1423
rect -87 -1495 -41 -1457
rect -87 -1529 -81 -1495
rect -47 -1529 -41 -1495
rect -87 -1567 -41 -1529
rect -87 -1601 -81 -1567
rect -47 -1601 -41 -1567
rect -87 -1639 -41 -1601
rect -87 -1673 -81 -1639
rect -47 -1673 -41 -1639
rect -87 -1711 -41 -1673
rect -87 -1745 -81 -1711
rect -47 -1745 -41 -1711
rect -87 -1783 -41 -1745
rect -87 -1817 -81 -1783
rect -47 -1817 -41 -1783
rect -87 -1855 -41 -1817
rect -87 -1889 -81 -1855
rect -47 -1889 -41 -1855
rect -87 -1927 -41 -1889
rect -87 -1961 -81 -1927
rect -47 -1961 -41 -1927
rect -87 -2000 -41 -1961
rect 41 1961 87 2000
rect 41 1927 47 1961
rect 81 1927 87 1961
rect 41 1889 87 1927
rect 41 1855 47 1889
rect 81 1855 87 1889
rect 41 1817 87 1855
rect 41 1783 47 1817
rect 81 1783 87 1817
rect 41 1745 87 1783
rect 41 1711 47 1745
rect 81 1711 87 1745
rect 41 1673 87 1711
rect 41 1639 47 1673
rect 81 1639 87 1673
rect 41 1601 87 1639
rect 41 1567 47 1601
rect 81 1567 87 1601
rect 41 1529 87 1567
rect 41 1495 47 1529
rect 81 1495 87 1529
rect 41 1457 87 1495
rect 41 1423 47 1457
rect 81 1423 87 1457
rect 41 1385 87 1423
rect 41 1351 47 1385
rect 81 1351 87 1385
rect 41 1313 87 1351
rect 41 1279 47 1313
rect 81 1279 87 1313
rect 41 1241 87 1279
rect 41 1207 47 1241
rect 81 1207 87 1241
rect 41 1169 87 1207
rect 41 1135 47 1169
rect 81 1135 87 1169
rect 41 1097 87 1135
rect 41 1063 47 1097
rect 81 1063 87 1097
rect 41 1025 87 1063
rect 41 991 47 1025
rect 81 991 87 1025
rect 41 953 87 991
rect 41 919 47 953
rect 81 919 87 953
rect 41 881 87 919
rect 41 847 47 881
rect 81 847 87 881
rect 41 809 87 847
rect 41 775 47 809
rect 81 775 87 809
rect 41 737 87 775
rect 41 703 47 737
rect 81 703 87 737
rect 41 665 87 703
rect 41 631 47 665
rect 81 631 87 665
rect 41 593 87 631
rect 41 559 47 593
rect 81 559 87 593
rect 41 521 87 559
rect 41 487 47 521
rect 81 487 87 521
rect 41 449 87 487
rect 41 415 47 449
rect 81 415 87 449
rect 41 377 87 415
rect 41 343 47 377
rect 81 343 87 377
rect 41 305 87 343
rect 41 271 47 305
rect 81 271 87 305
rect 41 233 87 271
rect 41 199 47 233
rect 81 199 87 233
rect 41 161 87 199
rect 41 127 47 161
rect 81 127 87 161
rect 41 89 87 127
rect 41 55 47 89
rect 81 55 87 89
rect 41 17 87 55
rect 41 -17 47 17
rect 81 -17 87 17
rect 41 -55 87 -17
rect 41 -89 47 -55
rect 81 -89 87 -55
rect 41 -127 87 -89
rect 41 -161 47 -127
rect 81 -161 87 -127
rect 41 -199 87 -161
rect 41 -233 47 -199
rect 81 -233 87 -199
rect 41 -271 87 -233
rect 41 -305 47 -271
rect 81 -305 87 -271
rect 41 -343 87 -305
rect 41 -377 47 -343
rect 81 -377 87 -343
rect 41 -415 87 -377
rect 41 -449 47 -415
rect 81 -449 87 -415
rect 41 -487 87 -449
rect 41 -521 47 -487
rect 81 -521 87 -487
rect 41 -559 87 -521
rect 41 -593 47 -559
rect 81 -593 87 -559
rect 41 -631 87 -593
rect 41 -665 47 -631
rect 81 -665 87 -631
rect 41 -703 87 -665
rect 41 -737 47 -703
rect 81 -737 87 -703
rect 41 -775 87 -737
rect 41 -809 47 -775
rect 81 -809 87 -775
rect 41 -847 87 -809
rect 41 -881 47 -847
rect 81 -881 87 -847
rect 41 -919 87 -881
rect 41 -953 47 -919
rect 81 -953 87 -919
rect 41 -991 87 -953
rect 41 -1025 47 -991
rect 81 -1025 87 -991
rect 41 -1063 87 -1025
rect 41 -1097 47 -1063
rect 81 -1097 87 -1063
rect 41 -1135 87 -1097
rect 41 -1169 47 -1135
rect 81 -1169 87 -1135
rect 41 -1207 87 -1169
rect 41 -1241 47 -1207
rect 81 -1241 87 -1207
rect 41 -1279 87 -1241
rect 41 -1313 47 -1279
rect 81 -1313 87 -1279
rect 41 -1351 87 -1313
rect 41 -1385 47 -1351
rect 81 -1385 87 -1351
rect 41 -1423 87 -1385
rect 41 -1457 47 -1423
rect 81 -1457 87 -1423
rect 41 -1495 87 -1457
rect 41 -1529 47 -1495
rect 81 -1529 87 -1495
rect 41 -1567 87 -1529
rect 41 -1601 47 -1567
rect 81 -1601 87 -1567
rect 41 -1639 87 -1601
rect 41 -1673 47 -1639
rect 81 -1673 87 -1639
rect 41 -1711 87 -1673
rect 41 -1745 47 -1711
rect 81 -1745 87 -1711
rect 41 -1783 87 -1745
rect 41 -1817 47 -1783
rect 81 -1817 87 -1783
rect 41 -1855 87 -1817
rect 41 -1889 47 -1855
rect 81 -1889 87 -1855
rect 41 -1927 87 -1889
rect 41 -1961 47 -1927
rect 81 -1961 87 -1927
rect 41 -2000 87 -1961
rect -31 -2038 31 -2032
rect -31 -2072 -17 -2038
rect 17 -2072 31 -2038
rect -31 -2078 31 -2072
<< properties >>
string FIXED_BBOX -178 -2157 178 2157
<< end >>
