magic
tech sky130A
magscale 1 2
timestamp 1637060811
<< pwell >>
rect -425 2547 3221 2834
rect -425 2052 -152 2547
rect -425 0 2724 2052
rect -425 -366 -152 0
rect 2948 -366 3221 2547
rect -425 -583 3221 -366
rect -425 -653 3220 -583
<< nmoslvt >>
rect 58 26 88 2026
rect 146 26 176 2026
rect 234 26 264 2026
rect 322 26 352 2026
rect 410 26 440 2026
rect 498 26 528 2026
rect 586 26 616 2026
rect 674 26 704 2026
rect 762 26 792 2026
rect 850 26 880 2026
rect 938 26 968 2026
rect 1026 26 1056 2026
rect 1114 26 1144 2026
rect 1202 26 1232 2026
rect 1290 26 1320 2026
rect 1378 26 1408 2026
rect 1466 26 1496 2026
rect 1554 26 1584 2026
rect 1642 26 1672 2026
rect 1730 26 1760 2026
rect 1818 26 1848 2026
rect 1906 26 1936 2026
rect 1994 26 2024 2026
rect 2082 26 2112 2026
rect 2170 26 2200 2026
rect 2258 26 2288 2026
rect 2346 26 2376 2026
rect 2434 26 2464 2026
rect 2522 26 2552 2026
rect 2610 26 2640 2026
<< ndiff >>
rect 0 1995 58 2026
rect 0 1961 12 1995
rect 46 1961 58 1995
rect 0 1927 58 1961
rect 0 1893 12 1927
rect 46 1893 58 1927
rect 0 1859 58 1893
rect 0 1825 12 1859
rect 46 1825 58 1859
rect 0 1791 58 1825
rect 0 1757 12 1791
rect 46 1757 58 1791
rect 0 1723 58 1757
rect 0 1689 12 1723
rect 46 1689 58 1723
rect 0 1655 58 1689
rect 0 1621 12 1655
rect 46 1621 58 1655
rect 0 1587 58 1621
rect 0 1553 12 1587
rect 46 1553 58 1587
rect 0 1519 58 1553
rect 0 1485 12 1519
rect 46 1485 58 1519
rect 0 1451 58 1485
rect 0 1417 12 1451
rect 46 1417 58 1451
rect 0 1383 58 1417
rect 0 1349 12 1383
rect 46 1349 58 1383
rect 0 1315 58 1349
rect 0 1281 12 1315
rect 46 1281 58 1315
rect 0 1247 58 1281
rect 0 1213 12 1247
rect 46 1213 58 1247
rect 0 1179 58 1213
rect 0 1145 12 1179
rect 46 1145 58 1179
rect 0 1111 58 1145
rect 0 1077 12 1111
rect 46 1077 58 1111
rect 0 1043 58 1077
rect 0 1009 12 1043
rect 46 1009 58 1043
rect 0 975 58 1009
rect 0 941 12 975
rect 46 941 58 975
rect 0 907 58 941
rect 0 873 12 907
rect 46 873 58 907
rect 0 839 58 873
rect 0 805 12 839
rect 46 805 58 839
rect 0 771 58 805
rect 0 737 12 771
rect 46 737 58 771
rect 0 703 58 737
rect 0 669 12 703
rect 46 669 58 703
rect 0 635 58 669
rect 0 601 12 635
rect 46 601 58 635
rect 0 567 58 601
rect 0 533 12 567
rect 46 533 58 567
rect 0 499 58 533
rect 0 465 12 499
rect 46 465 58 499
rect 0 431 58 465
rect 0 397 12 431
rect 46 397 58 431
rect 0 363 58 397
rect 0 329 12 363
rect 46 329 58 363
rect 0 295 58 329
rect 0 261 12 295
rect 46 261 58 295
rect 0 227 58 261
rect 0 193 12 227
rect 46 193 58 227
rect 0 159 58 193
rect 0 125 12 159
rect 46 125 58 159
rect 0 91 58 125
rect 0 57 12 91
rect 46 57 58 91
rect 0 26 58 57
rect 88 1995 146 2026
rect 88 1961 100 1995
rect 134 1961 146 1995
rect 88 1927 146 1961
rect 88 1893 100 1927
rect 134 1893 146 1927
rect 88 1859 146 1893
rect 88 1825 100 1859
rect 134 1825 146 1859
rect 88 1791 146 1825
rect 88 1757 100 1791
rect 134 1757 146 1791
rect 88 1723 146 1757
rect 88 1689 100 1723
rect 134 1689 146 1723
rect 88 1655 146 1689
rect 88 1621 100 1655
rect 134 1621 146 1655
rect 88 1587 146 1621
rect 88 1553 100 1587
rect 134 1553 146 1587
rect 88 1519 146 1553
rect 88 1485 100 1519
rect 134 1485 146 1519
rect 88 1451 146 1485
rect 88 1417 100 1451
rect 134 1417 146 1451
rect 88 1383 146 1417
rect 88 1349 100 1383
rect 134 1349 146 1383
rect 88 1315 146 1349
rect 88 1281 100 1315
rect 134 1281 146 1315
rect 88 1247 146 1281
rect 88 1213 100 1247
rect 134 1213 146 1247
rect 88 1179 146 1213
rect 88 1145 100 1179
rect 134 1145 146 1179
rect 88 1111 146 1145
rect 88 1077 100 1111
rect 134 1077 146 1111
rect 88 1043 146 1077
rect 88 1009 100 1043
rect 134 1009 146 1043
rect 88 975 146 1009
rect 88 941 100 975
rect 134 941 146 975
rect 88 907 146 941
rect 88 873 100 907
rect 134 873 146 907
rect 88 839 146 873
rect 88 805 100 839
rect 134 805 146 839
rect 88 771 146 805
rect 88 737 100 771
rect 134 737 146 771
rect 88 703 146 737
rect 88 669 100 703
rect 134 669 146 703
rect 88 635 146 669
rect 88 601 100 635
rect 134 601 146 635
rect 88 567 146 601
rect 88 533 100 567
rect 134 533 146 567
rect 88 499 146 533
rect 88 465 100 499
rect 134 465 146 499
rect 88 431 146 465
rect 88 397 100 431
rect 134 397 146 431
rect 88 363 146 397
rect 88 329 100 363
rect 134 329 146 363
rect 88 295 146 329
rect 88 261 100 295
rect 134 261 146 295
rect 88 227 146 261
rect 88 193 100 227
rect 134 193 146 227
rect 88 159 146 193
rect 88 125 100 159
rect 134 125 146 159
rect 88 91 146 125
rect 88 57 100 91
rect 134 57 146 91
rect 88 26 146 57
rect 176 1995 234 2026
rect 176 1961 188 1995
rect 222 1961 234 1995
rect 176 1927 234 1961
rect 176 1893 188 1927
rect 222 1893 234 1927
rect 176 1859 234 1893
rect 176 1825 188 1859
rect 222 1825 234 1859
rect 176 1791 234 1825
rect 176 1757 188 1791
rect 222 1757 234 1791
rect 176 1723 234 1757
rect 176 1689 188 1723
rect 222 1689 234 1723
rect 176 1655 234 1689
rect 176 1621 188 1655
rect 222 1621 234 1655
rect 176 1587 234 1621
rect 176 1553 188 1587
rect 222 1553 234 1587
rect 176 1519 234 1553
rect 176 1485 188 1519
rect 222 1485 234 1519
rect 176 1451 234 1485
rect 176 1417 188 1451
rect 222 1417 234 1451
rect 176 1383 234 1417
rect 176 1349 188 1383
rect 222 1349 234 1383
rect 176 1315 234 1349
rect 176 1281 188 1315
rect 222 1281 234 1315
rect 176 1247 234 1281
rect 176 1213 188 1247
rect 222 1213 234 1247
rect 176 1179 234 1213
rect 176 1145 188 1179
rect 222 1145 234 1179
rect 176 1111 234 1145
rect 176 1077 188 1111
rect 222 1077 234 1111
rect 176 1043 234 1077
rect 176 1009 188 1043
rect 222 1009 234 1043
rect 176 975 234 1009
rect 176 941 188 975
rect 222 941 234 975
rect 176 907 234 941
rect 176 873 188 907
rect 222 873 234 907
rect 176 839 234 873
rect 176 805 188 839
rect 222 805 234 839
rect 176 771 234 805
rect 176 737 188 771
rect 222 737 234 771
rect 176 703 234 737
rect 176 669 188 703
rect 222 669 234 703
rect 176 635 234 669
rect 176 601 188 635
rect 222 601 234 635
rect 176 567 234 601
rect 176 533 188 567
rect 222 533 234 567
rect 176 499 234 533
rect 176 465 188 499
rect 222 465 234 499
rect 176 431 234 465
rect 176 397 188 431
rect 222 397 234 431
rect 176 363 234 397
rect 176 329 188 363
rect 222 329 234 363
rect 176 295 234 329
rect 176 261 188 295
rect 222 261 234 295
rect 176 227 234 261
rect 176 193 188 227
rect 222 193 234 227
rect 176 159 234 193
rect 176 125 188 159
rect 222 125 234 159
rect 176 91 234 125
rect 176 57 188 91
rect 222 57 234 91
rect 176 26 234 57
rect 264 1995 322 2026
rect 264 1961 276 1995
rect 310 1961 322 1995
rect 264 1927 322 1961
rect 264 1893 276 1927
rect 310 1893 322 1927
rect 264 1859 322 1893
rect 264 1825 276 1859
rect 310 1825 322 1859
rect 264 1791 322 1825
rect 264 1757 276 1791
rect 310 1757 322 1791
rect 264 1723 322 1757
rect 264 1689 276 1723
rect 310 1689 322 1723
rect 264 1655 322 1689
rect 264 1621 276 1655
rect 310 1621 322 1655
rect 264 1587 322 1621
rect 264 1553 276 1587
rect 310 1553 322 1587
rect 264 1519 322 1553
rect 264 1485 276 1519
rect 310 1485 322 1519
rect 264 1451 322 1485
rect 264 1417 276 1451
rect 310 1417 322 1451
rect 264 1383 322 1417
rect 264 1349 276 1383
rect 310 1349 322 1383
rect 264 1315 322 1349
rect 264 1281 276 1315
rect 310 1281 322 1315
rect 264 1247 322 1281
rect 264 1213 276 1247
rect 310 1213 322 1247
rect 264 1179 322 1213
rect 264 1145 276 1179
rect 310 1145 322 1179
rect 264 1111 322 1145
rect 264 1077 276 1111
rect 310 1077 322 1111
rect 264 1043 322 1077
rect 264 1009 276 1043
rect 310 1009 322 1043
rect 264 975 322 1009
rect 264 941 276 975
rect 310 941 322 975
rect 264 907 322 941
rect 264 873 276 907
rect 310 873 322 907
rect 264 839 322 873
rect 264 805 276 839
rect 310 805 322 839
rect 264 771 322 805
rect 264 737 276 771
rect 310 737 322 771
rect 264 703 322 737
rect 264 669 276 703
rect 310 669 322 703
rect 264 635 322 669
rect 264 601 276 635
rect 310 601 322 635
rect 264 567 322 601
rect 264 533 276 567
rect 310 533 322 567
rect 264 499 322 533
rect 264 465 276 499
rect 310 465 322 499
rect 264 431 322 465
rect 264 397 276 431
rect 310 397 322 431
rect 264 363 322 397
rect 264 329 276 363
rect 310 329 322 363
rect 264 295 322 329
rect 264 261 276 295
rect 310 261 322 295
rect 264 227 322 261
rect 264 193 276 227
rect 310 193 322 227
rect 264 159 322 193
rect 264 125 276 159
rect 310 125 322 159
rect 264 91 322 125
rect 264 57 276 91
rect 310 57 322 91
rect 264 26 322 57
rect 352 1995 410 2026
rect 352 1961 364 1995
rect 398 1961 410 1995
rect 352 1927 410 1961
rect 352 1893 364 1927
rect 398 1893 410 1927
rect 352 1859 410 1893
rect 352 1825 364 1859
rect 398 1825 410 1859
rect 352 1791 410 1825
rect 352 1757 364 1791
rect 398 1757 410 1791
rect 352 1723 410 1757
rect 352 1689 364 1723
rect 398 1689 410 1723
rect 352 1655 410 1689
rect 352 1621 364 1655
rect 398 1621 410 1655
rect 352 1587 410 1621
rect 352 1553 364 1587
rect 398 1553 410 1587
rect 352 1519 410 1553
rect 352 1485 364 1519
rect 398 1485 410 1519
rect 352 1451 410 1485
rect 352 1417 364 1451
rect 398 1417 410 1451
rect 352 1383 410 1417
rect 352 1349 364 1383
rect 398 1349 410 1383
rect 352 1315 410 1349
rect 352 1281 364 1315
rect 398 1281 410 1315
rect 352 1247 410 1281
rect 352 1213 364 1247
rect 398 1213 410 1247
rect 352 1179 410 1213
rect 352 1145 364 1179
rect 398 1145 410 1179
rect 352 1111 410 1145
rect 352 1077 364 1111
rect 398 1077 410 1111
rect 352 1043 410 1077
rect 352 1009 364 1043
rect 398 1009 410 1043
rect 352 975 410 1009
rect 352 941 364 975
rect 398 941 410 975
rect 352 907 410 941
rect 352 873 364 907
rect 398 873 410 907
rect 352 839 410 873
rect 352 805 364 839
rect 398 805 410 839
rect 352 771 410 805
rect 352 737 364 771
rect 398 737 410 771
rect 352 703 410 737
rect 352 669 364 703
rect 398 669 410 703
rect 352 635 410 669
rect 352 601 364 635
rect 398 601 410 635
rect 352 567 410 601
rect 352 533 364 567
rect 398 533 410 567
rect 352 499 410 533
rect 352 465 364 499
rect 398 465 410 499
rect 352 431 410 465
rect 352 397 364 431
rect 398 397 410 431
rect 352 363 410 397
rect 352 329 364 363
rect 398 329 410 363
rect 352 295 410 329
rect 352 261 364 295
rect 398 261 410 295
rect 352 227 410 261
rect 352 193 364 227
rect 398 193 410 227
rect 352 159 410 193
rect 352 125 364 159
rect 398 125 410 159
rect 352 91 410 125
rect 352 57 364 91
rect 398 57 410 91
rect 352 26 410 57
rect 440 1995 498 2026
rect 440 1961 452 1995
rect 486 1961 498 1995
rect 440 1927 498 1961
rect 440 1893 452 1927
rect 486 1893 498 1927
rect 440 1859 498 1893
rect 440 1825 452 1859
rect 486 1825 498 1859
rect 440 1791 498 1825
rect 440 1757 452 1791
rect 486 1757 498 1791
rect 440 1723 498 1757
rect 440 1689 452 1723
rect 486 1689 498 1723
rect 440 1655 498 1689
rect 440 1621 452 1655
rect 486 1621 498 1655
rect 440 1587 498 1621
rect 440 1553 452 1587
rect 486 1553 498 1587
rect 440 1519 498 1553
rect 440 1485 452 1519
rect 486 1485 498 1519
rect 440 1451 498 1485
rect 440 1417 452 1451
rect 486 1417 498 1451
rect 440 1383 498 1417
rect 440 1349 452 1383
rect 486 1349 498 1383
rect 440 1315 498 1349
rect 440 1281 452 1315
rect 486 1281 498 1315
rect 440 1247 498 1281
rect 440 1213 452 1247
rect 486 1213 498 1247
rect 440 1179 498 1213
rect 440 1145 452 1179
rect 486 1145 498 1179
rect 440 1111 498 1145
rect 440 1077 452 1111
rect 486 1077 498 1111
rect 440 1043 498 1077
rect 440 1009 452 1043
rect 486 1009 498 1043
rect 440 975 498 1009
rect 440 941 452 975
rect 486 941 498 975
rect 440 907 498 941
rect 440 873 452 907
rect 486 873 498 907
rect 440 839 498 873
rect 440 805 452 839
rect 486 805 498 839
rect 440 771 498 805
rect 440 737 452 771
rect 486 737 498 771
rect 440 703 498 737
rect 440 669 452 703
rect 486 669 498 703
rect 440 635 498 669
rect 440 601 452 635
rect 486 601 498 635
rect 440 567 498 601
rect 440 533 452 567
rect 486 533 498 567
rect 440 499 498 533
rect 440 465 452 499
rect 486 465 498 499
rect 440 431 498 465
rect 440 397 452 431
rect 486 397 498 431
rect 440 363 498 397
rect 440 329 452 363
rect 486 329 498 363
rect 440 295 498 329
rect 440 261 452 295
rect 486 261 498 295
rect 440 227 498 261
rect 440 193 452 227
rect 486 193 498 227
rect 440 159 498 193
rect 440 125 452 159
rect 486 125 498 159
rect 440 91 498 125
rect 440 57 452 91
rect 486 57 498 91
rect 440 26 498 57
rect 528 1995 586 2026
rect 528 1961 540 1995
rect 574 1961 586 1995
rect 528 1927 586 1961
rect 528 1893 540 1927
rect 574 1893 586 1927
rect 528 1859 586 1893
rect 528 1825 540 1859
rect 574 1825 586 1859
rect 528 1791 586 1825
rect 528 1757 540 1791
rect 574 1757 586 1791
rect 528 1723 586 1757
rect 528 1689 540 1723
rect 574 1689 586 1723
rect 528 1655 586 1689
rect 528 1621 540 1655
rect 574 1621 586 1655
rect 528 1587 586 1621
rect 528 1553 540 1587
rect 574 1553 586 1587
rect 528 1519 586 1553
rect 528 1485 540 1519
rect 574 1485 586 1519
rect 528 1451 586 1485
rect 528 1417 540 1451
rect 574 1417 586 1451
rect 528 1383 586 1417
rect 528 1349 540 1383
rect 574 1349 586 1383
rect 528 1315 586 1349
rect 528 1281 540 1315
rect 574 1281 586 1315
rect 528 1247 586 1281
rect 528 1213 540 1247
rect 574 1213 586 1247
rect 528 1179 586 1213
rect 528 1145 540 1179
rect 574 1145 586 1179
rect 528 1111 586 1145
rect 528 1077 540 1111
rect 574 1077 586 1111
rect 528 1043 586 1077
rect 528 1009 540 1043
rect 574 1009 586 1043
rect 528 975 586 1009
rect 528 941 540 975
rect 574 941 586 975
rect 528 907 586 941
rect 528 873 540 907
rect 574 873 586 907
rect 528 839 586 873
rect 528 805 540 839
rect 574 805 586 839
rect 528 771 586 805
rect 528 737 540 771
rect 574 737 586 771
rect 528 703 586 737
rect 528 669 540 703
rect 574 669 586 703
rect 528 635 586 669
rect 528 601 540 635
rect 574 601 586 635
rect 528 567 586 601
rect 528 533 540 567
rect 574 533 586 567
rect 528 499 586 533
rect 528 465 540 499
rect 574 465 586 499
rect 528 431 586 465
rect 528 397 540 431
rect 574 397 586 431
rect 528 363 586 397
rect 528 329 540 363
rect 574 329 586 363
rect 528 295 586 329
rect 528 261 540 295
rect 574 261 586 295
rect 528 227 586 261
rect 528 193 540 227
rect 574 193 586 227
rect 528 159 586 193
rect 528 125 540 159
rect 574 125 586 159
rect 528 91 586 125
rect 528 57 540 91
rect 574 57 586 91
rect 528 26 586 57
rect 616 1995 674 2026
rect 616 1961 628 1995
rect 662 1961 674 1995
rect 616 1927 674 1961
rect 616 1893 628 1927
rect 662 1893 674 1927
rect 616 1859 674 1893
rect 616 1825 628 1859
rect 662 1825 674 1859
rect 616 1791 674 1825
rect 616 1757 628 1791
rect 662 1757 674 1791
rect 616 1723 674 1757
rect 616 1689 628 1723
rect 662 1689 674 1723
rect 616 1655 674 1689
rect 616 1621 628 1655
rect 662 1621 674 1655
rect 616 1587 674 1621
rect 616 1553 628 1587
rect 662 1553 674 1587
rect 616 1519 674 1553
rect 616 1485 628 1519
rect 662 1485 674 1519
rect 616 1451 674 1485
rect 616 1417 628 1451
rect 662 1417 674 1451
rect 616 1383 674 1417
rect 616 1349 628 1383
rect 662 1349 674 1383
rect 616 1315 674 1349
rect 616 1281 628 1315
rect 662 1281 674 1315
rect 616 1247 674 1281
rect 616 1213 628 1247
rect 662 1213 674 1247
rect 616 1179 674 1213
rect 616 1145 628 1179
rect 662 1145 674 1179
rect 616 1111 674 1145
rect 616 1077 628 1111
rect 662 1077 674 1111
rect 616 1043 674 1077
rect 616 1009 628 1043
rect 662 1009 674 1043
rect 616 975 674 1009
rect 616 941 628 975
rect 662 941 674 975
rect 616 907 674 941
rect 616 873 628 907
rect 662 873 674 907
rect 616 839 674 873
rect 616 805 628 839
rect 662 805 674 839
rect 616 771 674 805
rect 616 737 628 771
rect 662 737 674 771
rect 616 703 674 737
rect 616 669 628 703
rect 662 669 674 703
rect 616 635 674 669
rect 616 601 628 635
rect 662 601 674 635
rect 616 567 674 601
rect 616 533 628 567
rect 662 533 674 567
rect 616 499 674 533
rect 616 465 628 499
rect 662 465 674 499
rect 616 431 674 465
rect 616 397 628 431
rect 662 397 674 431
rect 616 363 674 397
rect 616 329 628 363
rect 662 329 674 363
rect 616 295 674 329
rect 616 261 628 295
rect 662 261 674 295
rect 616 227 674 261
rect 616 193 628 227
rect 662 193 674 227
rect 616 159 674 193
rect 616 125 628 159
rect 662 125 674 159
rect 616 91 674 125
rect 616 57 628 91
rect 662 57 674 91
rect 616 26 674 57
rect 704 1995 762 2026
rect 704 1961 716 1995
rect 750 1961 762 1995
rect 704 1927 762 1961
rect 704 1893 716 1927
rect 750 1893 762 1927
rect 704 1859 762 1893
rect 704 1825 716 1859
rect 750 1825 762 1859
rect 704 1791 762 1825
rect 704 1757 716 1791
rect 750 1757 762 1791
rect 704 1723 762 1757
rect 704 1689 716 1723
rect 750 1689 762 1723
rect 704 1655 762 1689
rect 704 1621 716 1655
rect 750 1621 762 1655
rect 704 1587 762 1621
rect 704 1553 716 1587
rect 750 1553 762 1587
rect 704 1519 762 1553
rect 704 1485 716 1519
rect 750 1485 762 1519
rect 704 1451 762 1485
rect 704 1417 716 1451
rect 750 1417 762 1451
rect 704 1383 762 1417
rect 704 1349 716 1383
rect 750 1349 762 1383
rect 704 1315 762 1349
rect 704 1281 716 1315
rect 750 1281 762 1315
rect 704 1247 762 1281
rect 704 1213 716 1247
rect 750 1213 762 1247
rect 704 1179 762 1213
rect 704 1145 716 1179
rect 750 1145 762 1179
rect 704 1111 762 1145
rect 704 1077 716 1111
rect 750 1077 762 1111
rect 704 1043 762 1077
rect 704 1009 716 1043
rect 750 1009 762 1043
rect 704 975 762 1009
rect 704 941 716 975
rect 750 941 762 975
rect 704 907 762 941
rect 704 873 716 907
rect 750 873 762 907
rect 704 839 762 873
rect 704 805 716 839
rect 750 805 762 839
rect 704 771 762 805
rect 704 737 716 771
rect 750 737 762 771
rect 704 703 762 737
rect 704 669 716 703
rect 750 669 762 703
rect 704 635 762 669
rect 704 601 716 635
rect 750 601 762 635
rect 704 567 762 601
rect 704 533 716 567
rect 750 533 762 567
rect 704 499 762 533
rect 704 465 716 499
rect 750 465 762 499
rect 704 431 762 465
rect 704 397 716 431
rect 750 397 762 431
rect 704 363 762 397
rect 704 329 716 363
rect 750 329 762 363
rect 704 295 762 329
rect 704 261 716 295
rect 750 261 762 295
rect 704 227 762 261
rect 704 193 716 227
rect 750 193 762 227
rect 704 159 762 193
rect 704 125 716 159
rect 750 125 762 159
rect 704 91 762 125
rect 704 57 716 91
rect 750 57 762 91
rect 704 26 762 57
rect 792 1995 850 2026
rect 792 1961 804 1995
rect 838 1961 850 1995
rect 792 1927 850 1961
rect 792 1893 804 1927
rect 838 1893 850 1927
rect 792 1859 850 1893
rect 792 1825 804 1859
rect 838 1825 850 1859
rect 792 1791 850 1825
rect 792 1757 804 1791
rect 838 1757 850 1791
rect 792 1723 850 1757
rect 792 1689 804 1723
rect 838 1689 850 1723
rect 792 1655 850 1689
rect 792 1621 804 1655
rect 838 1621 850 1655
rect 792 1587 850 1621
rect 792 1553 804 1587
rect 838 1553 850 1587
rect 792 1519 850 1553
rect 792 1485 804 1519
rect 838 1485 850 1519
rect 792 1451 850 1485
rect 792 1417 804 1451
rect 838 1417 850 1451
rect 792 1383 850 1417
rect 792 1349 804 1383
rect 838 1349 850 1383
rect 792 1315 850 1349
rect 792 1281 804 1315
rect 838 1281 850 1315
rect 792 1247 850 1281
rect 792 1213 804 1247
rect 838 1213 850 1247
rect 792 1179 850 1213
rect 792 1145 804 1179
rect 838 1145 850 1179
rect 792 1111 850 1145
rect 792 1077 804 1111
rect 838 1077 850 1111
rect 792 1043 850 1077
rect 792 1009 804 1043
rect 838 1009 850 1043
rect 792 975 850 1009
rect 792 941 804 975
rect 838 941 850 975
rect 792 907 850 941
rect 792 873 804 907
rect 838 873 850 907
rect 792 839 850 873
rect 792 805 804 839
rect 838 805 850 839
rect 792 771 850 805
rect 792 737 804 771
rect 838 737 850 771
rect 792 703 850 737
rect 792 669 804 703
rect 838 669 850 703
rect 792 635 850 669
rect 792 601 804 635
rect 838 601 850 635
rect 792 567 850 601
rect 792 533 804 567
rect 838 533 850 567
rect 792 499 850 533
rect 792 465 804 499
rect 838 465 850 499
rect 792 431 850 465
rect 792 397 804 431
rect 838 397 850 431
rect 792 363 850 397
rect 792 329 804 363
rect 838 329 850 363
rect 792 295 850 329
rect 792 261 804 295
rect 838 261 850 295
rect 792 227 850 261
rect 792 193 804 227
rect 838 193 850 227
rect 792 159 850 193
rect 792 125 804 159
rect 838 125 850 159
rect 792 91 850 125
rect 792 57 804 91
rect 838 57 850 91
rect 792 26 850 57
rect 880 1995 938 2026
rect 880 1961 892 1995
rect 926 1961 938 1995
rect 880 1927 938 1961
rect 880 1893 892 1927
rect 926 1893 938 1927
rect 880 1859 938 1893
rect 880 1825 892 1859
rect 926 1825 938 1859
rect 880 1791 938 1825
rect 880 1757 892 1791
rect 926 1757 938 1791
rect 880 1723 938 1757
rect 880 1689 892 1723
rect 926 1689 938 1723
rect 880 1655 938 1689
rect 880 1621 892 1655
rect 926 1621 938 1655
rect 880 1587 938 1621
rect 880 1553 892 1587
rect 926 1553 938 1587
rect 880 1519 938 1553
rect 880 1485 892 1519
rect 926 1485 938 1519
rect 880 1451 938 1485
rect 880 1417 892 1451
rect 926 1417 938 1451
rect 880 1383 938 1417
rect 880 1349 892 1383
rect 926 1349 938 1383
rect 880 1315 938 1349
rect 880 1281 892 1315
rect 926 1281 938 1315
rect 880 1247 938 1281
rect 880 1213 892 1247
rect 926 1213 938 1247
rect 880 1179 938 1213
rect 880 1145 892 1179
rect 926 1145 938 1179
rect 880 1111 938 1145
rect 880 1077 892 1111
rect 926 1077 938 1111
rect 880 1043 938 1077
rect 880 1009 892 1043
rect 926 1009 938 1043
rect 880 975 938 1009
rect 880 941 892 975
rect 926 941 938 975
rect 880 907 938 941
rect 880 873 892 907
rect 926 873 938 907
rect 880 839 938 873
rect 880 805 892 839
rect 926 805 938 839
rect 880 771 938 805
rect 880 737 892 771
rect 926 737 938 771
rect 880 703 938 737
rect 880 669 892 703
rect 926 669 938 703
rect 880 635 938 669
rect 880 601 892 635
rect 926 601 938 635
rect 880 567 938 601
rect 880 533 892 567
rect 926 533 938 567
rect 880 499 938 533
rect 880 465 892 499
rect 926 465 938 499
rect 880 431 938 465
rect 880 397 892 431
rect 926 397 938 431
rect 880 363 938 397
rect 880 329 892 363
rect 926 329 938 363
rect 880 295 938 329
rect 880 261 892 295
rect 926 261 938 295
rect 880 227 938 261
rect 880 193 892 227
rect 926 193 938 227
rect 880 159 938 193
rect 880 125 892 159
rect 926 125 938 159
rect 880 91 938 125
rect 880 57 892 91
rect 926 57 938 91
rect 880 26 938 57
rect 968 1995 1026 2026
rect 968 1961 980 1995
rect 1014 1961 1026 1995
rect 968 1927 1026 1961
rect 968 1893 980 1927
rect 1014 1893 1026 1927
rect 968 1859 1026 1893
rect 968 1825 980 1859
rect 1014 1825 1026 1859
rect 968 1791 1026 1825
rect 968 1757 980 1791
rect 1014 1757 1026 1791
rect 968 1723 1026 1757
rect 968 1689 980 1723
rect 1014 1689 1026 1723
rect 968 1655 1026 1689
rect 968 1621 980 1655
rect 1014 1621 1026 1655
rect 968 1587 1026 1621
rect 968 1553 980 1587
rect 1014 1553 1026 1587
rect 968 1519 1026 1553
rect 968 1485 980 1519
rect 1014 1485 1026 1519
rect 968 1451 1026 1485
rect 968 1417 980 1451
rect 1014 1417 1026 1451
rect 968 1383 1026 1417
rect 968 1349 980 1383
rect 1014 1349 1026 1383
rect 968 1315 1026 1349
rect 968 1281 980 1315
rect 1014 1281 1026 1315
rect 968 1247 1026 1281
rect 968 1213 980 1247
rect 1014 1213 1026 1247
rect 968 1179 1026 1213
rect 968 1145 980 1179
rect 1014 1145 1026 1179
rect 968 1111 1026 1145
rect 968 1077 980 1111
rect 1014 1077 1026 1111
rect 968 1043 1026 1077
rect 968 1009 980 1043
rect 1014 1009 1026 1043
rect 968 975 1026 1009
rect 968 941 980 975
rect 1014 941 1026 975
rect 968 907 1026 941
rect 968 873 980 907
rect 1014 873 1026 907
rect 968 839 1026 873
rect 968 805 980 839
rect 1014 805 1026 839
rect 968 771 1026 805
rect 968 737 980 771
rect 1014 737 1026 771
rect 968 703 1026 737
rect 968 669 980 703
rect 1014 669 1026 703
rect 968 635 1026 669
rect 968 601 980 635
rect 1014 601 1026 635
rect 968 567 1026 601
rect 968 533 980 567
rect 1014 533 1026 567
rect 968 499 1026 533
rect 968 465 980 499
rect 1014 465 1026 499
rect 968 431 1026 465
rect 968 397 980 431
rect 1014 397 1026 431
rect 968 363 1026 397
rect 968 329 980 363
rect 1014 329 1026 363
rect 968 295 1026 329
rect 968 261 980 295
rect 1014 261 1026 295
rect 968 227 1026 261
rect 968 193 980 227
rect 1014 193 1026 227
rect 968 159 1026 193
rect 968 125 980 159
rect 1014 125 1026 159
rect 968 91 1026 125
rect 968 57 980 91
rect 1014 57 1026 91
rect 968 26 1026 57
rect 1056 1995 1114 2026
rect 1056 1961 1068 1995
rect 1102 1961 1114 1995
rect 1056 1927 1114 1961
rect 1056 1893 1068 1927
rect 1102 1893 1114 1927
rect 1056 1859 1114 1893
rect 1056 1825 1068 1859
rect 1102 1825 1114 1859
rect 1056 1791 1114 1825
rect 1056 1757 1068 1791
rect 1102 1757 1114 1791
rect 1056 1723 1114 1757
rect 1056 1689 1068 1723
rect 1102 1689 1114 1723
rect 1056 1655 1114 1689
rect 1056 1621 1068 1655
rect 1102 1621 1114 1655
rect 1056 1587 1114 1621
rect 1056 1553 1068 1587
rect 1102 1553 1114 1587
rect 1056 1519 1114 1553
rect 1056 1485 1068 1519
rect 1102 1485 1114 1519
rect 1056 1451 1114 1485
rect 1056 1417 1068 1451
rect 1102 1417 1114 1451
rect 1056 1383 1114 1417
rect 1056 1349 1068 1383
rect 1102 1349 1114 1383
rect 1056 1315 1114 1349
rect 1056 1281 1068 1315
rect 1102 1281 1114 1315
rect 1056 1247 1114 1281
rect 1056 1213 1068 1247
rect 1102 1213 1114 1247
rect 1056 1179 1114 1213
rect 1056 1145 1068 1179
rect 1102 1145 1114 1179
rect 1056 1111 1114 1145
rect 1056 1077 1068 1111
rect 1102 1077 1114 1111
rect 1056 1043 1114 1077
rect 1056 1009 1068 1043
rect 1102 1009 1114 1043
rect 1056 975 1114 1009
rect 1056 941 1068 975
rect 1102 941 1114 975
rect 1056 907 1114 941
rect 1056 873 1068 907
rect 1102 873 1114 907
rect 1056 839 1114 873
rect 1056 805 1068 839
rect 1102 805 1114 839
rect 1056 771 1114 805
rect 1056 737 1068 771
rect 1102 737 1114 771
rect 1056 703 1114 737
rect 1056 669 1068 703
rect 1102 669 1114 703
rect 1056 635 1114 669
rect 1056 601 1068 635
rect 1102 601 1114 635
rect 1056 567 1114 601
rect 1056 533 1068 567
rect 1102 533 1114 567
rect 1056 499 1114 533
rect 1056 465 1068 499
rect 1102 465 1114 499
rect 1056 431 1114 465
rect 1056 397 1068 431
rect 1102 397 1114 431
rect 1056 363 1114 397
rect 1056 329 1068 363
rect 1102 329 1114 363
rect 1056 295 1114 329
rect 1056 261 1068 295
rect 1102 261 1114 295
rect 1056 227 1114 261
rect 1056 193 1068 227
rect 1102 193 1114 227
rect 1056 159 1114 193
rect 1056 125 1068 159
rect 1102 125 1114 159
rect 1056 91 1114 125
rect 1056 57 1068 91
rect 1102 57 1114 91
rect 1056 26 1114 57
rect 1144 1995 1202 2026
rect 1144 1961 1156 1995
rect 1190 1961 1202 1995
rect 1144 1927 1202 1961
rect 1144 1893 1156 1927
rect 1190 1893 1202 1927
rect 1144 1859 1202 1893
rect 1144 1825 1156 1859
rect 1190 1825 1202 1859
rect 1144 1791 1202 1825
rect 1144 1757 1156 1791
rect 1190 1757 1202 1791
rect 1144 1723 1202 1757
rect 1144 1689 1156 1723
rect 1190 1689 1202 1723
rect 1144 1655 1202 1689
rect 1144 1621 1156 1655
rect 1190 1621 1202 1655
rect 1144 1587 1202 1621
rect 1144 1553 1156 1587
rect 1190 1553 1202 1587
rect 1144 1519 1202 1553
rect 1144 1485 1156 1519
rect 1190 1485 1202 1519
rect 1144 1451 1202 1485
rect 1144 1417 1156 1451
rect 1190 1417 1202 1451
rect 1144 1383 1202 1417
rect 1144 1349 1156 1383
rect 1190 1349 1202 1383
rect 1144 1315 1202 1349
rect 1144 1281 1156 1315
rect 1190 1281 1202 1315
rect 1144 1247 1202 1281
rect 1144 1213 1156 1247
rect 1190 1213 1202 1247
rect 1144 1179 1202 1213
rect 1144 1145 1156 1179
rect 1190 1145 1202 1179
rect 1144 1111 1202 1145
rect 1144 1077 1156 1111
rect 1190 1077 1202 1111
rect 1144 1043 1202 1077
rect 1144 1009 1156 1043
rect 1190 1009 1202 1043
rect 1144 975 1202 1009
rect 1144 941 1156 975
rect 1190 941 1202 975
rect 1144 907 1202 941
rect 1144 873 1156 907
rect 1190 873 1202 907
rect 1144 839 1202 873
rect 1144 805 1156 839
rect 1190 805 1202 839
rect 1144 771 1202 805
rect 1144 737 1156 771
rect 1190 737 1202 771
rect 1144 703 1202 737
rect 1144 669 1156 703
rect 1190 669 1202 703
rect 1144 635 1202 669
rect 1144 601 1156 635
rect 1190 601 1202 635
rect 1144 567 1202 601
rect 1144 533 1156 567
rect 1190 533 1202 567
rect 1144 499 1202 533
rect 1144 465 1156 499
rect 1190 465 1202 499
rect 1144 431 1202 465
rect 1144 397 1156 431
rect 1190 397 1202 431
rect 1144 363 1202 397
rect 1144 329 1156 363
rect 1190 329 1202 363
rect 1144 295 1202 329
rect 1144 261 1156 295
rect 1190 261 1202 295
rect 1144 227 1202 261
rect 1144 193 1156 227
rect 1190 193 1202 227
rect 1144 159 1202 193
rect 1144 125 1156 159
rect 1190 125 1202 159
rect 1144 91 1202 125
rect 1144 57 1156 91
rect 1190 57 1202 91
rect 1144 26 1202 57
rect 1232 1995 1290 2026
rect 1232 1961 1244 1995
rect 1278 1961 1290 1995
rect 1232 1927 1290 1961
rect 1232 1893 1244 1927
rect 1278 1893 1290 1927
rect 1232 1859 1290 1893
rect 1232 1825 1244 1859
rect 1278 1825 1290 1859
rect 1232 1791 1290 1825
rect 1232 1757 1244 1791
rect 1278 1757 1290 1791
rect 1232 1723 1290 1757
rect 1232 1689 1244 1723
rect 1278 1689 1290 1723
rect 1232 1655 1290 1689
rect 1232 1621 1244 1655
rect 1278 1621 1290 1655
rect 1232 1587 1290 1621
rect 1232 1553 1244 1587
rect 1278 1553 1290 1587
rect 1232 1519 1290 1553
rect 1232 1485 1244 1519
rect 1278 1485 1290 1519
rect 1232 1451 1290 1485
rect 1232 1417 1244 1451
rect 1278 1417 1290 1451
rect 1232 1383 1290 1417
rect 1232 1349 1244 1383
rect 1278 1349 1290 1383
rect 1232 1315 1290 1349
rect 1232 1281 1244 1315
rect 1278 1281 1290 1315
rect 1232 1247 1290 1281
rect 1232 1213 1244 1247
rect 1278 1213 1290 1247
rect 1232 1179 1290 1213
rect 1232 1145 1244 1179
rect 1278 1145 1290 1179
rect 1232 1111 1290 1145
rect 1232 1077 1244 1111
rect 1278 1077 1290 1111
rect 1232 1043 1290 1077
rect 1232 1009 1244 1043
rect 1278 1009 1290 1043
rect 1232 975 1290 1009
rect 1232 941 1244 975
rect 1278 941 1290 975
rect 1232 907 1290 941
rect 1232 873 1244 907
rect 1278 873 1290 907
rect 1232 839 1290 873
rect 1232 805 1244 839
rect 1278 805 1290 839
rect 1232 771 1290 805
rect 1232 737 1244 771
rect 1278 737 1290 771
rect 1232 703 1290 737
rect 1232 669 1244 703
rect 1278 669 1290 703
rect 1232 635 1290 669
rect 1232 601 1244 635
rect 1278 601 1290 635
rect 1232 567 1290 601
rect 1232 533 1244 567
rect 1278 533 1290 567
rect 1232 499 1290 533
rect 1232 465 1244 499
rect 1278 465 1290 499
rect 1232 431 1290 465
rect 1232 397 1244 431
rect 1278 397 1290 431
rect 1232 363 1290 397
rect 1232 329 1244 363
rect 1278 329 1290 363
rect 1232 295 1290 329
rect 1232 261 1244 295
rect 1278 261 1290 295
rect 1232 227 1290 261
rect 1232 193 1244 227
rect 1278 193 1290 227
rect 1232 159 1290 193
rect 1232 125 1244 159
rect 1278 125 1290 159
rect 1232 91 1290 125
rect 1232 57 1244 91
rect 1278 57 1290 91
rect 1232 26 1290 57
rect 1320 1995 1378 2026
rect 1320 1961 1332 1995
rect 1366 1961 1378 1995
rect 1320 1927 1378 1961
rect 1320 1893 1332 1927
rect 1366 1893 1378 1927
rect 1320 1859 1378 1893
rect 1320 1825 1332 1859
rect 1366 1825 1378 1859
rect 1320 1791 1378 1825
rect 1320 1757 1332 1791
rect 1366 1757 1378 1791
rect 1320 1723 1378 1757
rect 1320 1689 1332 1723
rect 1366 1689 1378 1723
rect 1320 1655 1378 1689
rect 1320 1621 1332 1655
rect 1366 1621 1378 1655
rect 1320 1587 1378 1621
rect 1320 1553 1332 1587
rect 1366 1553 1378 1587
rect 1320 1519 1378 1553
rect 1320 1485 1332 1519
rect 1366 1485 1378 1519
rect 1320 1451 1378 1485
rect 1320 1417 1332 1451
rect 1366 1417 1378 1451
rect 1320 1383 1378 1417
rect 1320 1349 1332 1383
rect 1366 1349 1378 1383
rect 1320 1315 1378 1349
rect 1320 1281 1332 1315
rect 1366 1281 1378 1315
rect 1320 1247 1378 1281
rect 1320 1213 1332 1247
rect 1366 1213 1378 1247
rect 1320 1179 1378 1213
rect 1320 1145 1332 1179
rect 1366 1145 1378 1179
rect 1320 1111 1378 1145
rect 1320 1077 1332 1111
rect 1366 1077 1378 1111
rect 1320 1043 1378 1077
rect 1320 1009 1332 1043
rect 1366 1009 1378 1043
rect 1320 975 1378 1009
rect 1320 941 1332 975
rect 1366 941 1378 975
rect 1320 907 1378 941
rect 1320 873 1332 907
rect 1366 873 1378 907
rect 1320 839 1378 873
rect 1320 805 1332 839
rect 1366 805 1378 839
rect 1320 771 1378 805
rect 1320 737 1332 771
rect 1366 737 1378 771
rect 1320 703 1378 737
rect 1320 669 1332 703
rect 1366 669 1378 703
rect 1320 635 1378 669
rect 1320 601 1332 635
rect 1366 601 1378 635
rect 1320 567 1378 601
rect 1320 533 1332 567
rect 1366 533 1378 567
rect 1320 499 1378 533
rect 1320 465 1332 499
rect 1366 465 1378 499
rect 1320 431 1378 465
rect 1320 397 1332 431
rect 1366 397 1378 431
rect 1320 363 1378 397
rect 1320 329 1332 363
rect 1366 329 1378 363
rect 1320 295 1378 329
rect 1320 261 1332 295
rect 1366 261 1378 295
rect 1320 227 1378 261
rect 1320 193 1332 227
rect 1366 193 1378 227
rect 1320 159 1378 193
rect 1320 125 1332 159
rect 1366 125 1378 159
rect 1320 91 1378 125
rect 1320 57 1332 91
rect 1366 57 1378 91
rect 1320 26 1378 57
rect 1408 1995 1466 2026
rect 1408 1961 1420 1995
rect 1454 1961 1466 1995
rect 1408 1927 1466 1961
rect 1408 1893 1420 1927
rect 1454 1893 1466 1927
rect 1408 1859 1466 1893
rect 1408 1825 1420 1859
rect 1454 1825 1466 1859
rect 1408 1791 1466 1825
rect 1408 1757 1420 1791
rect 1454 1757 1466 1791
rect 1408 1723 1466 1757
rect 1408 1689 1420 1723
rect 1454 1689 1466 1723
rect 1408 1655 1466 1689
rect 1408 1621 1420 1655
rect 1454 1621 1466 1655
rect 1408 1587 1466 1621
rect 1408 1553 1420 1587
rect 1454 1553 1466 1587
rect 1408 1519 1466 1553
rect 1408 1485 1420 1519
rect 1454 1485 1466 1519
rect 1408 1451 1466 1485
rect 1408 1417 1420 1451
rect 1454 1417 1466 1451
rect 1408 1383 1466 1417
rect 1408 1349 1420 1383
rect 1454 1349 1466 1383
rect 1408 1315 1466 1349
rect 1408 1281 1420 1315
rect 1454 1281 1466 1315
rect 1408 1247 1466 1281
rect 1408 1213 1420 1247
rect 1454 1213 1466 1247
rect 1408 1179 1466 1213
rect 1408 1145 1420 1179
rect 1454 1145 1466 1179
rect 1408 1111 1466 1145
rect 1408 1077 1420 1111
rect 1454 1077 1466 1111
rect 1408 1043 1466 1077
rect 1408 1009 1420 1043
rect 1454 1009 1466 1043
rect 1408 975 1466 1009
rect 1408 941 1420 975
rect 1454 941 1466 975
rect 1408 907 1466 941
rect 1408 873 1420 907
rect 1454 873 1466 907
rect 1408 839 1466 873
rect 1408 805 1420 839
rect 1454 805 1466 839
rect 1408 771 1466 805
rect 1408 737 1420 771
rect 1454 737 1466 771
rect 1408 703 1466 737
rect 1408 669 1420 703
rect 1454 669 1466 703
rect 1408 635 1466 669
rect 1408 601 1420 635
rect 1454 601 1466 635
rect 1408 567 1466 601
rect 1408 533 1420 567
rect 1454 533 1466 567
rect 1408 499 1466 533
rect 1408 465 1420 499
rect 1454 465 1466 499
rect 1408 431 1466 465
rect 1408 397 1420 431
rect 1454 397 1466 431
rect 1408 363 1466 397
rect 1408 329 1420 363
rect 1454 329 1466 363
rect 1408 295 1466 329
rect 1408 261 1420 295
rect 1454 261 1466 295
rect 1408 227 1466 261
rect 1408 193 1420 227
rect 1454 193 1466 227
rect 1408 159 1466 193
rect 1408 125 1420 159
rect 1454 125 1466 159
rect 1408 91 1466 125
rect 1408 57 1420 91
rect 1454 57 1466 91
rect 1408 26 1466 57
rect 1496 1995 1554 2026
rect 1496 1961 1508 1995
rect 1542 1961 1554 1995
rect 1496 1927 1554 1961
rect 1496 1893 1508 1927
rect 1542 1893 1554 1927
rect 1496 1859 1554 1893
rect 1496 1825 1508 1859
rect 1542 1825 1554 1859
rect 1496 1791 1554 1825
rect 1496 1757 1508 1791
rect 1542 1757 1554 1791
rect 1496 1723 1554 1757
rect 1496 1689 1508 1723
rect 1542 1689 1554 1723
rect 1496 1655 1554 1689
rect 1496 1621 1508 1655
rect 1542 1621 1554 1655
rect 1496 1587 1554 1621
rect 1496 1553 1508 1587
rect 1542 1553 1554 1587
rect 1496 1519 1554 1553
rect 1496 1485 1508 1519
rect 1542 1485 1554 1519
rect 1496 1451 1554 1485
rect 1496 1417 1508 1451
rect 1542 1417 1554 1451
rect 1496 1383 1554 1417
rect 1496 1349 1508 1383
rect 1542 1349 1554 1383
rect 1496 1315 1554 1349
rect 1496 1281 1508 1315
rect 1542 1281 1554 1315
rect 1496 1247 1554 1281
rect 1496 1213 1508 1247
rect 1542 1213 1554 1247
rect 1496 1179 1554 1213
rect 1496 1145 1508 1179
rect 1542 1145 1554 1179
rect 1496 1111 1554 1145
rect 1496 1077 1508 1111
rect 1542 1077 1554 1111
rect 1496 1043 1554 1077
rect 1496 1009 1508 1043
rect 1542 1009 1554 1043
rect 1496 975 1554 1009
rect 1496 941 1508 975
rect 1542 941 1554 975
rect 1496 907 1554 941
rect 1496 873 1508 907
rect 1542 873 1554 907
rect 1496 839 1554 873
rect 1496 805 1508 839
rect 1542 805 1554 839
rect 1496 771 1554 805
rect 1496 737 1508 771
rect 1542 737 1554 771
rect 1496 703 1554 737
rect 1496 669 1508 703
rect 1542 669 1554 703
rect 1496 635 1554 669
rect 1496 601 1508 635
rect 1542 601 1554 635
rect 1496 567 1554 601
rect 1496 533 1508 567
rect 1542 533 1554 567
rect 1496 499 1554 533
rect 1496 465 1508 499
rect 1542 465 1554 499
rect 1496 431 1554 465
rect 1496 397 1508 431
rect 1542 397 1554 431
rect 1496 363 1554 397
rect 1496 329 1508 363
rect 1542 329 1554 363
rect 1496 295 1554 329
rect 1496 261 1508 295
rect 1542 261 1554 295
rect 1496 227 1554 261
rect 1496 193 1508 227
rect 1542 193 1554 227
rect 1496 159 1554 193
rect 1496 125 1508 159
rect 1542 125 1554 159
rect 1496 91 1554 125
rect 1496 57 1508 91
rect 1542 57 1554 91
rect 1496 26 1554 57
rect 1584 1995 1642 2026
rect 1584 1961 1596 1995
rect 1630 1961 1642 1995
rect 1584 1927 1642 1961
rect 1584 1893 1596 1927
rect 1630 1893 1642 1927
rect 1584 1859 1642 1893
rect 1584 1825 1596 1859
rect 1630 1825 1642 1859
rect 1584 1791 1642 1825
rect 1584 1757 1596 1791
rect 1630 1757 1642 1791
rect 1584 1723 1642 1757
rect 1584 1689 1596 1723
rect 1630 1689 1642 1723
rect 1584 1655 1642 1689
rect 1584 1621 1596 1655
rect 1630 1621 1642 1655
rect 1584 1587 1642 1621
rect 1584 1553 1596 1587
rect 1630 1553 1642 1587
rect 1584 1519 1642 1553
rect 1584 1485 1596 1519
rect 1630 1485 1642 1519
rect 1584 1451 1642 1485
rect 1584 1417 1596 1451
rect 1630 1417 1642 1451
rect 1584 1383 1642 1417
rect 1584 1349 1596 1383
rect 1630 1349 1642 1383
rect 1584 1315 1642 1349
rect 1584 1281 1596 1315
rect 1630 1281 1642 1315
rect 1584 1247 1642 1281
rect 1584 1213 1596 1247
rect 1630 1213 1642 1247
rect 1584 1179 1642 1213
rect 1584 1145 1596 1179
rect 1630 1145 1642 1179
rect 1584 1111 1642 1145
rect 1584 1077 1596 1111
rect 1630 1077 1642 1111
rect 1584 1043 1642 1077
rect 1584 1009 1596 1043
rect 1630 1009 1642 1043
rect 1584 975 1642 1009
rect 1584 941 1596 975
rect 1630 941 1642 975
rect 1584 907 1642 941
rect 1584 873 1596 907
rect 1630 873 1642 907
rect 1584 839 1642 873
rect 1584 805 1596 839
rect 1630 805 1642 839
rect 1584 771 1642 805
rect 1584 737 1596 771
rect 1630 737 1642 771
rect 1584 703 1642 737
rect 1584 669 1596 703
rect 1630 669 1642 703
rect 1584 635 1642 669
rect 1584 601 1596 635
rect 1630 601 1642 635
rect 1584 567 1642 601
rect 1584 533 1596 567
rect 1630 533 1642 567
rect 1584 499 1642 533
rect 1584 465 1596 499
rect 1630 465 1642 499
rect 1584 431 1642 465
rect 1584 397 1596 431
rect 1630 397 1642 431
rect 1584 363 1642 397
rect 1584 329 1596 363
rect 1630 329 1642 363
rect 1584 295 1642 329
rect 1584 261 1596 295
rect 1630 261 1642 295
rect 1584 227 1642 261
rect 1584 193 1596 227
rect 1630 193 1642 227
rect 1584 159 1642 193
rect 1584 125 1596 159
rect 1630 125 1642 159
rect 1584 91 1642 125
rect 1584 57 1596 91
rect 1630 57 1642 91
rect 1584 26 1642 57
rect 1672 1995 1730 2026
rect 1672 1961 1684 1995
rect 1718 1961 1730 1995
rect 1672 1927 1730 1961
rect 1672 1893 1684 1927
rect 1718 1893 1730 1927
rect 1672 1859 1730 1893
rect 1672 1825 1684 1859
rect 1718 1825 1730 1859
rect 1672 1791 1730 1825
rect 1672 1757 1684 1791
rect 1718 1757 1730 1791
rect 1672 1723 1730 1757
rect 1672 1689 1684 1723
rect 1718 1689 1730 1723
rect 1672 1655 1730 1689
rect 1672 1621 1684 1655
rect 1718 1621 1730 1655
rect 1672 1587 1730 1621
rect 1672 1553 1684 1587
rect 1718 1553 1730 1587
rect 1672 1519 1730 1553
rect 1672 1485 1684 1519
rect 1718 1485 1730 1519
rect 1672 1451 1730 1485
rect 1672 1417 1684 1451
rect 1718 1417 1730 1451
rect 1672 1383 1730 1417
rect 1672 1349 1684 1383
rect 1718 1349 1730 1383
rect 1672 1315 1730 1349
rect 1672 1281 1684 1315
rect 1718 1281 1730 1315
rect 1672 1247 1730 1281
rect 1672 1213 1684 1247
rect 1718 1213 1730 1247
rect 1672 1179 1730 1213
rect 1672 1145 1684 1179
rect 1718 1145 1730 1179
rect 1672 1111 1730 1145
rect 1672 1077 1684 1111
rect 1718 1077 1730 1111
rect 1672 1043 1730 1077
rect 1672 1009 1684 1043
rect 1718 1009 1730 1043
rect 1672 975 1730 1009
rect 1672 941 1684 975
rect 1718 941 1730 975
rect 1672 907 1730 941
rect 1672 873 1684 907
rect 1718 873 1730 907
rect 1672 839 1730 873
rect 1672 805 1684 839
rect 1718 805 1730 839
rect 1672 771 1730 805
rect 1672 737 1684 771
rect 1718 737 1730 771
rect 1672 703 1730 737
rect 1672 669 1684 703
rect 1718 669 1730 703
rect 1672 635 1730 669
rect 1672 601 1684 635
rect 1718 601 1730 635
rect 1672 567 1730 601
rect 1672 533 1684 567
rect 1718 533 1730 567
rect 1672 499 1730 533
rect 1672 465 1684 499
rect 1718 465 1730 499
rect 1672 431 1730 465
rect 1672 397 1684 431
rect 1718 397 1730 431
rect 1672 363 1730 397
rect 1672 329 1684 363
rect 1718 329 1730 363
rect 1672 295 1730 329
rect 1672 261 1684 295
rect 1718 261 1730 295
rect 1672 227 1730 261
rect 1672 193 1684 227
rect 1718 193 1730 227
rect 1672 159 1730 193
rect 1672 125 1684 159
rect 1718 125 1730 159
rect 1672 91 1730 125
rect 1672 57 1684 91
rect 1718 57 1730 91
rect 1672 26 1730 57
rect 1760 1995 1818 2026
rect 1760 1961 1772 1995
rect 1806 1961 1818 1995
rect 1760 1927 1818 1961
rect 1760 1893 1772 1927
rect 1806 1893 1818 1927
rect 1760 1859 1818 1893
rect 1760 1825 1772 1859
rect 1806 1825 1818 1859
rect 1760 1791 1818 1825
rect 1760 1757 1772 1791
rect 1806 1757 1818 1791
rect 1760 1723 1818 1757
rect 1760 1689 1772 1723
rect 1806 1689 1818 1723
rect 1760 1655 1818 1689
rect 1760 1621 1772 1655
rect 1806 1621 1818 1655
rect 1760 1587 1818 1621
rect 1760 1553 1772 1587
rect 1806 1553 1818 1587
rect 1760 1519 1818 1553
rect 1760 1485 1772 1519
rect 1806 1485 1818 1519
rect 1760 1451 1818 1485
rect 1760 1417 1772 1451
rect 1806 1417 1818 1451
rect 1760 1383 1818 1417
rect 1760 1349 1772 1383
rect 1806 1349 1818 1383
rect 1760 1315 1818 1349
rect 1760 1281 1772 1315
rect 1806 1281 1818 1315
rect 1760 1247 1818 1281
rect 1760 1213 1772 1247
rect 1806 1213 1818 1247
rect 1760 1179 1818 1213
rect 1760 1145 1772 1179
rect 1806 1145 1818 1179
rect 1760 1111 1818 1145
rect 1760 1077 1772 1111
rect 1806 1077 1818 1111
rect 1760 1043 1818 1077
rect 1760 1009 1772 1043
rect 1806 1009 1818 1043
rect 1760 975 1818 1009
rect 1760 941 1772 975
rect 1806 941 1818 975
rect 1760 907 1818 941
rect 1760 873 1772 907
rect 1806 873 1818 907
rect 1760 839 1818 873
rect 1760 805 1772 839
rect 1806 805 1818 839
rect 1760 771 1818 805
rect 1760 737 1772 771
rect 1806 737 1818 771
rect 1760 703 1818 737
rect 1760 669 1772 703
rect 1806 669 1818 703
rect 1760 635 1818 669
rect 1760 601 1772 635
rect 1806 601 1818 635
rect 1760 567 1818 601
rect 1760 533 1772 567
rect 1806 533 1818 567
rect 1760 499 1818 533
rect 1760 465 1772 499
rect 1806 465 1818 499
rect 1760 431 1818 465
rect 1760 397 1772 431
rect 1806 397 1818 431
rect 1760 363 1818 397
rect 1760 329 1772 363
rect 1806 329 1818 363
rect 1760 295 1818 329
rect 1760 261 1772 295
rect 1806 261 1818 295
rect 1760 227 1818 261
rect 1760 193 1772 227
rect 1806 193 1818 227
rect 1760 159 1818 193
rect 1760 125 1772 159
rect 1806 125 1818 159
rect 1760 91 1818 125
rect 1760 57 1772 91
rect 1806 57 1818 91
rect 1760 26 1818 57
rect 1848 1995 1906 2026
rect 1848 1961 1860 1995
rect 1894 1961 1906 1995
rect 1848 1927 1906 1961
rect 1848 1893 1860 1927
rect 1894 1893 1906 1927
rect 1848 1859 1906 1893
rect 1848 1825 1860 1859
rect 1894 1825 1906 1859
rect 1848 1791 1906 1825
rect 1848 1757 1860 1791
rect 1894 1757 1906 1791
rect 1848 1723 1906 1757
rect 1848 1689 1860 1723
rect 1894 1689 1906 1723
rect 1848 1655 1906 1689
rect 1848 1621 1860 1655
rect 1894 1621 1906 1655
rect 1848 1587 1906 1621
rect 1848 1553 1860 1587
rect 1894 1553 1906 1587
rect 1848 1519 1906 1553
rect 1848 1485 1860 1519
rect 1894 1485 1906 1519
rect 1848 1451 1906 1485
rect 1848 1417 1860 1451
rect 1894 1417 1906 1451
rect 1848 1383 1906 1417
rect 1848 1349 1860 1383
rect 1894 1349 1906 1383
rect 1848 1315 1906 1349
rect 1848 1281 1860 1315
rect 1894 1281 1906 1315
rect 1848 1247 1906 1281
rect 1848 1213 1860 1247
rect 1894 1213 1906 1247
rect 1848 1179 1906 1213
rect 1848 1145 1860 1179
rect 1894 1145 1906 1179
rect 1848 1111 1906 1145
rect 1848 1077 1860 1111
rect 1894 1077 1906 1111
rect 1848 1043 1906 1077
rect 1848 1009 1860 1043
rect 1894 1009 1906 1043
rect 1848 975 1906 1009
rect 1848 941 1860 975
rect 1894 941 1906 975
rect 1848 907 1906 941
rect 1848 873 1860 907
rect 1894 873 1906 907
rect 1848 839 1906 873
rect 1848 805 1860 839
rect 1894 805 1906 839
rect 1848 771 1906 805
rect 1848 737 1860 771
rect 1894 737 1906 771
rect 1848 703 1906 737
rect 1848 669 1860 703
rect 1894 669 1906 703
rect 1848 635 1906 669
rect 1848 601 1860 635
rect 1894 601 1906 635
rect 1848 567 1906 601
rect 1848 533 1860 567
rect 1894 533 1906 567
rect 1848 499 1906 533
rect 1848 465 1860 499
rect 1894 465 1906 499
rect 1848 431 1906 465
rect 1848 397 1860 431
rect 1894 397 1906 431
rect 1848 363 1906 397
rect 1848 329 1860 363
rect 1894 329 1906 363
rect 1848 295 1906 329
rect 1848 261 1860 295
rect 1894 261 1906 295
rect 1848 227 1906 261
rect 1848 193 1860 227
rect 1894 193 1906 227
rect 1848 159 1906 193
rect 1848 125 1860 159
rect 1894 125 1906 159
rect 1848 91 1906 125
rect 1848 57 1860 91
rect 1894 57 1906 91
rect 1848 26 1906 57
rect 1936 1995 1994 2026
rect 1936 1961 1948 1995
rect 1982 1961 1994 1995
rect 1936 1927 1994 1961
rect 1936 1893 1948 1927
rect 1982 1893 1994 1927
rect 1936 1859 1994 1893
rect 1936 1825 1948 1859
rect 1982 1825 1994 1859
rect 1936 1791 1994 1825
rect 1936 1757 1948 1791
rect 1982 1757 1994 1791
rect 1936 1723 1994 1757
rect 1936 1689 1948 1723
rect 1982 1689 1994 1723
rect 1936 1655 1994 1689
rect 1936 1621 1948 1655
rect 1982 1621 1994 1655
rect 1936 1587 1994 1621
rect 1936 1553 1948 1587
rect 1982 1553 1994 1587
rect 1936 1519 1994 1553
rect 1936 1485 1948 1519
rect 1982 1485 1994 1519
rect 1936 1451 1994 1485
rect 1936 1417 1948 1451
rect 1982 1417 1994 1451
rect 1936 1383 1994 1417
rect 1936 1349 1948 1383
rect 1982 1349 1994 1383
rect 1936 1315 1994 1349
rect 1936 1281 1948 1315
rect 1982 1281 1994 1315
rect 1936 1247 1994 1281
rect 1936 1213 1948 1247
rect 1982 1213 1994 1247
rect 1936 1179 1994 1213
rect 1936 1145 1948 1179
rect 1982 1145 1994 1179
rect 1936 1111 1994 1145
rect 1936 1077 1948 1111
rect 1982 1077 1994 1111
rect 1936 1043 1994 1077
rect 1936 1009 1948 1043
rect 1982 1009 1994 1043
rect 1936 975 1994 1009
rect 1936 941 1948 975
rect 1982 941 1994 975
rect 1936 907 1994 941
rect 1936 873 1948 907
rect 1982 873 1994 907
rect 1936 839 1994 873
rect 1936 805 1948 839
rect 1982 805 1994 839
rect 1936 771 1994 805
rect 1936 737 1948 771
rect 1982 737 1994 771
rect 1936 703 1994 737
rect 1936 669 1948 703
rect 1982 669 1994 703
rect 1936 635 1994 669
rect 1936 601 1948 635
rect 1982 601 1994 635
rect 1936 567 1994 601
rect 1936 533 1948 567
rect 1982 533 1994 567
rect 1936 499 1994 533
rect 1936 465 1948 499
rect 1982 465 1994 499
rect 1936 431 1994 465
rect 1936 397 1948 431
rect 1982 397 1994 431
rect 1936 363 1994 397
rect 1936 329 1948 363
rect 1982 329 1994 363
rect 1936 295 1994 329
rect 1936 261 1948 295
rect 1982 261 1994 295
rect 1936 227 1994 261
rect 1936 193 1948 227
rect 1982 193 1994 227
rect 1936 159 1994 193
rect 1936 125 1948 159
rect 1982 125 1994 159
rect 1936 91 1994 125
rect 1936 57 1948 91
rect 1982 57 1994 91
rect 1936 26 1994 57
rect 2024 1995 2082 2026
rect 2024 1961 2036 1995
rect 2070 1961 2082 1995
rect 2024 1927 2082 1961
rect 2024 1893 2036 1927
rect 2070 1893 2082 1927
rect 2024 1859 2082 1893
rect 2024 1825 2036 1859
rect 2070 1825 2082 1859
rect 2024 1791 2082 1825
rect 2024 1757 2036 1791
rect 2070 1757 2082 1791
rect 2024 1723 2082 1757
rect 2024 1689 2036 1723
rect 2070 1689 2082 1723
rect 2024 1655 2082 1689
rect 2024 1621 2036 1655
rect 2070 1621 2082 1655
rect 2024 1587 2082 1621
rect 2024 1553 2036 1587
rect 2070 1553 2082 1587
rect 2024 1519 2082 1553
rect 2024 1485 2036 1519
rect 2070 1485 2082 1519
rect 2024 1451 2082 1485
rect 2024 1417 2036 1451
rect 2070 1417 2082 1451
rect 2024 1383 2082 1417
rect 2024 1349 2036 1383
rect 2070 1349 2082 1383
rect 2024 1315 2082 1349
rect 2024 1281 2036 1315
rect 2070 1281 2082 1315
rect 2024 1247 2082 1281
rect 2024 1213 2036 1247
rect 2070 1213 2082 1247
rect 2024 1179 2082 1213
rect 2024 1145 2036 1179
rect 2070 1145 2082 1179
rect 2024 1111 2082 1145
rect 2024 1077 2036 1111
rect 2070 1077 2082 1111
rect 2024 1043 2082 1077
rect 2024 1009 2036 1043
rect 2070 1009 2082 1043
rect 2024 975 2082 1009
rect 2024 941 2036 975
rect 2070 941 2082 975
rect 2024 907 2082 941
rect 2024 873 2036 907
rect 2070 873 2082 907
rect 2024 839 2082 873
rect 2024 805 2036 839
rect 2070 805 2082 839
rect 2024 771 2082 805
rect 2024 737 2036 771
rect 2070 737 2082 771
rect 2024 703 2082 737
rect 2024 669 2036 703
rect 2070 669 2082 703
rect 2024 635 2082 669
rect 2024 601 2036 635
rect 2070 601 2082 635
rect 2024 567 2082 601
rect 2024 533 2036 567
rect 2070 533 2082 567
rect 2024 499 2082 533
rect 2024 465 2036 499
rect 2070 465 2082 499
rect 2024 431 2082 465
rect 2024 397 2036 431
rect 2070 397 2082 431
rect 2024 363 2082 397
rect 2024 329 2036 363
rect 2070 329 2082 363
rect 2024 295 2082 329
rect 2024 261 2036 295
rect 2070 261 2082 295
rect 2024 227 2082 261
rect 2024 193 2036 227
rect 2070 193 2082 227
rect 2024 159 2082 193
rect 2024 125 2036 159
rect 2070 125 2082 159
rect 2024 91 2082 125
rect 2024 57 2036 91
rect 2070 57 2082 91
rect 2024 26 2082 57
rect 2112 1995 2170 2026
rect 2112 1961 2124 1995
rect 2158 1961 2170 1995
rect 2112 1927 2170 1961
rect 2112 1893 2124 1927
rect 2158 1893 2170 1927
rect 2112 1859 2170 1893
rect 2112 1825 2124 1859
rect 2158 1825 2170 1859
rect 2112 1791 2170 1825
rect 2112 1757 2124 1791
rect 2158 1757 2170 1791
rect 2112 1723 2170 1757
rect 2112 1689 2124 1723
rect 2158 1689 2170 1723
rect 2112 1655 2170 1689
rect 2112 1621 2124 1655
rect 2158 1621 2170 1655
rect 2112 1587 2170 1621
rect 2112 1553 2124 1587
rect 2158 1553 2170 1587
rect 2112 1519 2170 1553
rect 2112 1485 2124 1519
rect 2158 1485 2170 1519
rect 2112 1451 2170 1485
rect 2112 1417 2124 1451
rect 2158 1417 2170 1451
rect 2112 1383 2170 1417
rect 2112 1349 2124 1383
rect 2158 1349 2170 1383
rect 2112 1315 2170 1349
rect 2112 1281 2124 1315
rect 2158 1281 2170 1315
rect 2112 1247 2170 1281
rect 2112 1213 2124 1247
rect 2158 1213 2170 1247
rect 2112 1179 2170 1213
rect 2112 1145 2124 1179
rect 2158 1145 2170 1179
rect 2112 1111 2170 1145
rect 2112 1077 2124 1111
rect 2158 1077 2170 1111
rect 2112 1043 2170 1077
rect 2112 1009 2124 1043
rect 2158 1009 2170 1043
rect 2112 975 2170 1009
rect 2112 941 2124 975
rect 2158 941 2170 975
rect 2112 907 2170 941
rect 2112 873 2124 907
rect 2158 873 2170 907
rect 2112 839 2170 873
rect 2112 805 2124 839
rect 2158 805 2170 839
rect 2112 771 2170 805
rect 2112 737 2124 771
rect 2158 737 2170 771
rect 2112 703 2170 737
rect 2112 669 2124 703
rect 2158 669 2170 703
rect 2112 635 2170 669
rect 2112 601 2124 635
rect 2158 601 2170 635
rect 2112 567 2170 601
rect 2112 533 2124 567
rect 2158 533 2170 567
rect 2112 499 2170 533
rect 2112 465 2124 499
rect 2158 465 2170 499
rect 2112 431 2170 465
rect 2112 397 2124 431
rect 2158 397 2170 431
rect 2112 363 2170 397
rect 2112 329 2124 363
rect 2158 329 2170 363
rect 2112 295 2170 329
rect 2112 261 2124 295
rect 2158 261 2170 295
rect 2112 227 2170 261
rect 2112 193 2124 227
rect 2158 193 2170 227
rect 2112 159 2170 193
rect 2112 125 2124 159
rect 2158 125 2170 159
rect 2112 91 2170 125
rect 2112 57 2124 91
rect 2158 57 2170 91
rect 2112 26 2170 57
rect 2200 1995 2258 2026
rect 2200 1961 2212 1995
rect 2246 1961 2258 1995
rect 2200 1927 2258 1961
rect 2200 1893 2212 1927
rect 2246 1893 2258 1927
rect 2200 1859 2258 1893
rect 2200 1825 2212 1859
rect 2246 1825 2258 1859
rect 2200 1791 2258 1825
rect 2200 1757 2212 1791
rect 2246 1757 2258 1791
rect 2200 1723 2258 1757
rect 2200 1689 2212 1723
rect 2246 1689 2258 1723
rect 2200 1655 2258 1689
rect 2200 1621 2212 1655
rect 2246 1621 2258 1655
rect 2200 1587 2258 1621
rect 2200 1553 2212 1587
rect 2246 1553 2258 1587
rect 2200 1519 2258 1553
rect 2200 1485 2212 1519
rect 2246 1485 2258 1519
rect 2200 1451 2258 1485
rect 2200 1417 2212 1451
rect 2246 1417 2258 1451
rect 2200 1383 2258 1417
rect 2200 1349 2212 1383
rect 2246 1349 2258 1383
rect 2200 1315 2258 1349
rect 2200 1281 2212 1315
rect 2246 1281 2258 1315
rect 2200 1247 2258 1281
rect 2200 1213 2212 1247
rect 2246 1213 2258 1247
rect 2200 1179 2258 1213
rect 2200 1145 2212 1179
rect 2246 1145 2258 1179
rect 2200 1111 2258 1145
rect 2200 1077 2212 1111
rect 2246 1077 2258 1111
rect 2200 1043 2258 1077
rect 2200 1009 2212 1043
rect 2246 1009 2258 1043
rect 2200 975 2258 1009
rect 2200 941 2212 975
rect 2246 941 2258 975
rect 2200 907 2258 941
rect 2200 873 2212 907
rect 2246 873 2258 907
rect 2200 839 2258 873
rect 2200 805 2212 839
rect 2246 805 2258 839
rect 2200 771 2258 805
rect 2200 737 2212 771
rect 2246 737 2258 771
rect 2200 703 2258 737
rect 2200 669 2212 703
rect 2246 669 2258 703
rect 2200 635 2258 669
rect 2200 601 2212 635
rect 2246 601 2258 635
rect 2200 567 2258 601
rect 2200 533 2212 567
rect 2246 533 2258 567
rect 2200 499 2258 533
rect 2200 465 2212 499
rect 2246 465 2258 499
rect 2200 431 2258 465
rect 2200 397 2212 431
rect 2246 397 2258 431
rect 2200 363 2258 397
rect 2200 329 2212 363
rect 2246 329 2258 363
rect 2200 295 2258 329
rect 2200 261 2212 295
rect 2246 261 2258 295
rect 2200 227 2258 261
rect 2200 193 2212 227
rect 2246 193 2258 227
rect 2200 159 2258 193
rect 2200 125 2212 159
rect 2246 125 2258 159
rect 2200 91 2258 125
rect 2200 57 2212 91
rect 2246 57 2258 91
rect 2200 26 2258 57
rect 2288 1995 2346 2026
rect 2288 1961 2300 1995
rect 2334 1961 2346 1995
rect 2288 1927 2346 1961
rect 2288 1893 2300 1927
rect 2334 1893 2346 1927
rect 2288 1859 2346 1893
rect 2288 1825 2300 1859
rect 2334 1825 2346 1859
rect 2288 1791 2346 1825
rect 2288 1757 2300 1791
rect 2334 1757 2346 1791
rect 2288 1723 2346 1757
rect 2288 1689 2300 1723
rect 2334 1689 2346 1723
rect 2288 1655 2346 1689
rect 2288 1621 2300 1655
rect 2334 1621 2346 1655
rect 2288 1587 2346 1621
rect 2288 1553 2300 1587
rect 2334 1553 2346 1587
rect 2288 1519 2346 1553
rect 2288 1485 2300 1519
rect 2334 1485 2346 1519
rect 2288 1451 2346 1485
rect 2288 1417 2300 1451
rect 2334 1417 2346 1451
rect 2288 1383 2346 1417
rect 2288 1349 2300 1383
rect 2334 1349 2346 1383
rect 2288 1315 2346 1349
rect 2288 1281 2300 1315
rect 2334 1281 2346 1315
rect 2288 1247 2346 1281
rect 2288 1213 2300 1247
rect 2334 1213 2346 1247
rect 2288 1179 2346 1213
rect 2288 1145 2300 1179
rect 2334 1145 2346 1179
rect 2288 1111 2346 1145
rect 2288 1077 2300 1111
rect 2334 1077 2346 1111
rect 2288 1043 2346 1077
rect 2288 1009 2300 1043
rect 2334 1009 2346 1043
rect 2288 975 2346 1009
rect 2288 941 2300 975
rect 2334 941 2346 975
rect 2288 907 2346 941
rect 2288 873 2300 907
rect 2334 873 2346 907
rect 2288 839 2346 873
rect 2288 805 2300 839
rect 2334 805 2346 839
rect 2288 771 2346 805
rect 2288 737 2300 771
rect 2334 737 2346 771
rect 2288 703 2346 737
rect 2288 669 2300 703
rect 2334 669 2346 703
rect 2288 635 2346 669
rect 2288 601 2300 635
rect 2334 601 2346 635
rect 2288 567 2346 601
rect 2288 533 2300 567
rect 2334 533 2346 567
rect 2288 499 2346 533
rect 2288 465 2300 499
rect 2334 465 2346 499
rect 2288 431 2346 465
rect 2288 397 2300 431
rect 2334 397 2346 431
rect 2288 363 2346 397
rect 2288 329 2300 363
rect 2334 329 2346 363
rect 2288 295 2346 329
rect 2288 261 2300 295
rect 2334 261 2346 295
rect 2288 227 2346 261
rect 2288 193 2300 227
rect 2334 193 2346 227
rect 2288 159 2346 193
rect 2288 125 2300 159
rect 2334 125 2346 159
rect 2288 91 2346 125
rect 2288 57 2300 91
rect 2334 57 2346 91
rect 2288 26 2346 57
rect 2376 1995 2434 2026
rect 2376 1961 2388 1995
rect 2422 1961 2434 1995
rect 2376 1927 2434 1961
rect 2376 1893 2388 1927
rect 2422 1893 2434 1927
rect 2376 1859 2434 1893
rect 2376 1825 2388 1859
rect 2422 1825 2434 1859
rect 2376 1791 2434 1825
rect 2376 1757 2388 1791
rect 2422 1757 2434 1791
rect 2376 1723 2434 1757
rect 2376 1689 2388 1723
rect 2422 1689 2434 1723
rect 2376 1655 2434 1689
rect 2376 1621 2388 1655
rect 2422 1621 2434 1655
rect 2376 1587 2434 1621
rect 2376 1553 2388 1587
rect 2422 1553 2434 1587
rect 2376 1519 2434 1553
rect 2376 1485 2388 1519
rect 2422 1485 2434 1519
rect 2376 1451 2434 1485
rect 2376 1417 2388 1451
rect 2422 1417 2434 1451
rect 2376 1383 2434 1417
rect 2376 1349 2388 1383
rect 2422 1349 2434 1383
rect 2376 1315 2434 1349
rect 2376 1281 2388 1315
rect 2422 1281 2434 1315
rect 2376 1247 2434 1281
rect 2376 1213 2388 1247
rect 2422 1213 2434 1247
rect 2376 1179 2434 1213
rect 2376 1145 2388 1179
rect 2422 1145 2434 1179
rect 2376 1111 2434 1145
rect 2376 1077 2388 1111
rect 2422 1077 2434 1111
rect 2376 1043 2434 1077
rect 2376 1009 2388 1043
rect 2422 1009 2434 1043
rect 2376 975 2434 1009
rect 2376 941 2388 975
rect 2422 941 2434 975
rect 2376 907 2434 941
rect 2376 873 2388 907
rect 2422 873 2434 907
rect 2376 839 2434 873
rect 2376 805 2388 839
rect 2422 805 2434 839
rect 2376 771 2434 805
rect 2376 737 2388 771
rect 2422 737 2434 771
rect 2376 703 2434 737
rect 2376 669 2388 703
rect 2422 669 2434 703
rect 2376 635 2434 669
rect 2376 601 2388 635
rect 2422 601 2434 635
rect 2376 567 2434 601
rect 2376 533 2388 567
rect 2422 533 2434 567
rect 2376 499 2434 533
rect 2376 465 2388 499
rect 2422 465 2434 499
rect 2376 431 2434 465
rect 2376 397 2388 431
rect 2422 397 2434 431
rect 2376 363 2434 397
rect 2376 329 2388 363
rect 2422 329 2434 363
rect 2376 295 2434 329
rect 2376 261 2388 295
rect 2422 261 2434 295
rect 2376 227 2434 261
rect 2376 193 2388 227
rect 2422 193 2434 227
rect 2376 159 2434 193
rect 2376 125 2388 159
rect 2422 125 2434 159
rect 2376 91 2434 125
rect 2376 57 2388 91
rect 2422 57 2434 91
rect 2376 26 2434 57
rect 2464 1995 2522 2026
rect 2464 1961 2476 1995
rect 2510 1961 2522 1995
rect 2464 1927 2522 1961
rect 2464 1893 2476 1927
rect 2510 1893 2522 1927
rect 2464 1859 2522 1893
rect 2464 1825 2476 1859
rect 2510 1825 2522 1859
rect 2464 1791 2522 1825
rect 2464 1757 2476 1791
rect 2510 1757 2522 1791
rect 2464 1723 2522 1757
rect 2464 1689 2476 1723
rect 2510 1689 2522 1723
rect 2464 1655 2522 1689
rect 2464 1621 2476 1655
rect 2510 1621 2522 1655
rect 2464 1587 2522 1621
rect 2464 1553 2476 1587
rect 2510 1553 2522 1587
rect 2464 1519 2522 1553
rect 2464 1485 2476 1519
rect 2510 1485 2522 1519
rect 2464 1451 2522 1485
rect 2464 1417 2476 1451
rect 2510 1417 2522 1451
rect 2464 1383 2522 1417
rect 2464 1349 2476 1383
rect 2510 1349 2522 1383
rect 2464 1315 2522 1349
rect 2464 1281 2476 1315
rect 2510 1281 2522 1315
rect 2464 1247 2522 1281
rect 2464 1213 2476 1247
rect 2510 1213 2522 1247
rect 2464 1179 2522 1213
rect 2464 1145 2476 1179
rect 2510 1145 2522 1179
rect 2464 1111 2522 1145
rect 2464 1077 2476 1111
rect 2510 1077 2522 1111
rect 2464 1043 2522 1077
rect 2464 1009 2476 1043
rect 2510 1009 2522 1043
rect 2464 975 2522 1009
rect 2464 941 2476 975
rect 2510 941 2522 975
rect 2464 907 2522 941
rect 2464 873 2476 907
rect 2510 873 2522 907
rect 2464 839 2522 873
rect 2464 805 2476 839
rect 2510 805 2522 839
rect 2464 771 2522 805
rect 2464 737 2476 771
rect 2510 737 2522 771
rect 2464 703 2522 737
rect 2464 669 2476 703
rect 2510 669 2522 703
rect 2464 635 2522 669
rect 2464 601 2476 635
rect 2510 601 2522 635
rect 2464 567 2522 601
rect 2464 533 2476 567
rect 2510 533 2522 567
rect 2464 499 2522 533
rect 2464 465 2476 499
rect 2510 465 2522 499
rect 2464 431 2522 465
rect 2464 397 2476 431
rect 2510 397 2522 431
rect 2464 363 2522 397
rect 2464 329 2476 363
rect 2510 329 2522 363
rect 2464 295 2522 329
rect 2464 261 2476 295
rect 2510 261 2522 295
rect 2464 227 2522 261
rect 2464 193 2476 227
rect 2510 193 2522 227
rect 2464 159 2522 193
rect 2464 125 2476 159
rect 2510 125 2522 159
rect 2464 91 2522 125
rect 2464 57 2476 91
rect 2510 57 2522 91
rect 2464 26 2522 57
rect 2552 1995 2610 2026
rect 2552 1961 2564 1995
rect 2598 1961 2610 1995
rect 2552 1927 2610 1961
rect 2552 1893 2564 1927
rect 2598 1893 2610 1927
rect 2552 1859 2610 1893
rect 2552 1825 2564 1859
rect 2598 1825 2610 1859
rect 2552 1791 2610 1825
rect 2552 1757 2564 1791
rect 2598 1757 2610 1791
rect 2552 1723 2610 1757
rect 2552 1689 2564 1723
rect 2598 1689 2610 1723
rect 2552 1655 2610 1689
rect 2552 1621 2564 1655
rect 2598 1621 2610 1655
rect 2552 1587 2610 1621
rect 2552 1553 2564 1587
rect 2598 1553 2610 1587
rect 2552 1519 2610 1553
rect 2552 1485 2564 1519
rect 2598 1485 2610 1519
rect 2552 1451 2610 1485
rect 2552 1417 2564 1451
rect 2598 1417 2610 1451
rect 2552 1383 2610 1417
rect 2552 1349 2564 1383
rect 2598 1349 2610 1383
rect 2552 1315 2610 1349
rect 2552 1281 2564 1315
rect 2598 1281 2610 1315
rect 2552 1247 2610 1281
rect 2552 1213 2564 1247
rect 2598 1213 2610 1247
rect 2552 1179 2610 1213
rect 2552 1145 2564 1179
rect 2598 1145 2610 1179
rect 2552 1111 2610 1145
rect 2552 1077 2564 1111
rect 2598 1077 2610 1111
rect 2552 1043 2610 1077
rect 2552 1009 2564 1043
rect 2598 1009 2610 1043
rect 2552 975 2610 1009
rect 2552 941 2564 975
rect 2598 941 2610 975
rect 2552 907 2610 941
rect 2552 873 2564 907
rect 2598 873 2610 907
rect 2552 839 2610 873
rect 2552 805 2564 839
rect 2598 805 2610 839
rect 2552 771 2610 805
rect 2552 737 2564 771
rect 2598 737 2610 771
rect 2552 703 2610 737
rect 2552 669 2564 703
rect 2598 669 2610 703
rect 2552 635 2610 669
rect 2552 601 2564 635
rect 2598 601 2610 635
rect 2552 567 2610 601
rect 2552 533 2564 567
rect 2598 533 2610 567
rect 2552 499 2610 533
rect 2552 465 2564 499
rect 2598 465 2610 499
rect 2552 431 2610 465
rect 2552 397 2564 431
rect 2598 397 2610 431
rect 2552 363 2610 397
rect 2552 329 2564 363
rect 2598 329 2610 363
rect 2552 295 2610 329
rect 2552 261 2564 295
rect 2598 261 2610 295
rect 2552 227 2610 261
rect 2552 193 2564 227
rect 2598 193 2610 227
rect 2552 159 2610 193
rect 2552 125 2564 159
rect 2598 125 2610 159
rect 2552 91 2610 125
rect 2552 57 2564 91
rect 2598 57 2610 91
rect 2552 26 2610 57
rect 2640 1995 2698 2026
rect 2640 1961 2652 1995
rect 2686 1961 2698 1995
rect 2640 1927 2698 1961
rect 2640 1893 2652 1927
rect 2686 1893 2698 1927
rect 2640 1859 2698 1893
rect 2640 1825 2652 1859
rect 2686 1825 2698 1859
rect 2640 1791 2698 1825
rect 2640 1757 2652 1791
rect 2686 1757 2698 1791
rect 2640 1723 2698 1757
rect 2640 1689 2652 1723
rect 2686 1689 2698 1723
rect 2640 1655 2698 1689
rect 2640 1621 2652 1655
rect 2686 1621 2698 1655
rect 2640 1587 2698 1621
rect 2640 1553 2652 1587
rect 2686 1553 2698 1587
rect 2640 1519 2698 1553
rect 2640 1485 2652 1519
rect 2686 1485 2698 1519
rect 2640 1451 2698 1485
rect 2640 1417 2652 1451
rect 2686 1417 2698 1451
rect 2640 1383 2698 1417
rect 2640 1349 2652 1383
rect 2686 1349 2698 1383
rect 2640 1315 2698 1349
rect 2640 1281 2652 1315
rect 2686 1281 2698 1315
rect 2640 1247 2698 1281
rect 2640 1213 2652 1247
rect 2686 1213 2698 1247
rect 2640 1179 2698 1213
rect 2640 1145 2652 1179
rect 2686 1145 2698 1179
rect 2640 1111 2698 1145
rect 2640 1077 2652 1111
rect 2686 1077 2698 1111
rect 2640 1043 2698 1077
rect 2640 1009 2652 1043
rect 2686 1009 2698 1043
rect 2640 975 2698 1009
rect 2640 941 2652 975
rect 2686 941 2698 975
rect 2640 907 2698 941
rect 2640 873 2652 907
rect 2686 873 2698 907
rect 2640 839 2698 873
rect 2640 805 2652 839
rect 2686 805 2698 839
rect 2640 771 2698 805
rect 2640 737 2652 771
rect 2686 737 2698 771
rect 2640 703 2698 737
rect 2640 669 2652 703
rect 2686 669 2698 703
rect 2640 635 2698 669
rect 2640 601 2652 635
rect 2686 601 2698 635
rect 2640 567 2698 601
rect 2640 533 2652 567
rect 2686 533 2698 567
rect 2640 499 2698 533
rect 2640 465 2652 499
rect 2686 465 2698 499
rect 2640 431 2698 465
rect 2640 397 2652 431
rect 2686 397 2698 431
rect 2640 363 2698 397
rect 2640 329 2652 363
rect 2686 329 2698 363
rect 2640 295 2698 329
rect 2640 261 2652 295
rect 2686 261 2698 295
rect 2640 227 2698 261
rect 2640 193 2652 227
rect 2686 193 2698 227
rect 2640 159 2698 193
rect 2640 125 2652 159
rect 2686 125 2698 159
rect 2640 91 2698 125
rect 2640 57 2652 91
rect 2686 57 2698 91
rect 2640 26 2698 57
<< ndiffc >>
rect 12 1961 46 1995
rect 12 1893 46 1927
rect 12 1825 46 1859
rect 12 1757 46 1791
rect 12 1689 46 1723
rect 12 1621 46 1655
rect 12 1553 46 1587
rect 12 1485 46 1519
rect 12 1417 46 1451
rect 12 1349 46 1383
rect 12 1281 46 1315
rect 12 1213 46 1247
rect 12 1145 46 1179
rect 12 1077 46 1111
rect 12 1009 46 1043
rect 12 941 46 975
rect 12 873 46 907
rect 12 805 46 839
rect 12 737 46 771
rect 12 669 46 703
rect 12 601 46 635
rect 12 533 46 567
rect 12 465 46 499
rect 12 397 46 431
rect 12 329 46 363
rect 12 261 46 295
rect 12 193 46 227
rect 12 125 46 159
rect 12 57 46 91
rect 100 1961 134 1995
rect 100 1893 134 1927
rect 100 1825 134 1859
rect 100 1757 134 1791
rect 100 1689 134 1723
rect 100 1621 134 1655
rect 100 1553 134 1587
rect 100 1485 134 1519
rect 100 1417 134 1451
rect 100 1349 134 1383
rect 100 1281 134 1315
rect 100 1213 134 1247
rect 100 1145 134 1179
rect 100 1077 134 1111
rect 100 1009 134 1043
rect 100 941 134 975
rect 100 873 134 907
rect 100 805 134 839
rect 100 737 134 771
rect 100 669 134 703
rect 100 601 134 635
rect 100 533 134 567
rect 100 465 134 499
rect 100 397 134 431
rect 100 329 134 363
rect 100 261 134 295
rect 100 193 134 227
rect 100 125 134 159
rect 100 57 134 91
rect 188 1961 222 1995
rect 188 1893 222 1927
rect 188 1825 222 1859
rect 188 1757 222 1791
rect 188 1689 222 1723
rect 188 1621 222 1655
rect 188 1553 222 1587
rect 188 1485 222 1519
rect 188 1417 222 1451
rect 188 1349 222 1383
rect 188 1281 222 1315
rect 188 1213 222 1247
rect 188 1145 222 1179
rect 188 1077 222 1111
rect 188 1009 222 1043
rect 188 941 222 975
rect 188 873 222 907
rect 188 805 222 839
rect 188 737 222 771
rect 188 669 222 703
rect 188 601 222 635
rect 188 533 222 567
rect 188 465 222 499
rect 188 397 222 431
rect 188 329 222 363
rect 188 261 222 295
rect 188 193 222 227
rect 188 125 222 159
rect 188 57 222 91
rect 276 1961 310 1995
rect 276 1893 310 1927
rect 276 1825 310 1859
rect 276 1757 310 1791
rect 276 1689 310 1723
rect 276 1621 310 1655
rect 276 1553 310 1587
rect 276 1485 310 1519
rect 276 1417 310 1451
rect 276 1349 310 1383
rect 276 1281 310 1315
rect 276 1213 310 1247
rect 276 1145 310 1179
rect 276 1077 310 1111
rect 276 1009 310 1043
rect 276 941 310 975
rect 276 873 310 907
rect 276 805 310 839
rect 276 737 310 771
rect 276 669 310 703
rect 276 601 310 635
rect 276 533 310 567
rect 276 465 310 499
rect 276 397 310 431
rect 276 329 310 363
rect 276 261 310 295
rect 276 193 310 227
rect 276 125 310 159
rect 276 57 310 91
rect 364 1961 398 1995
rect 364 1893 398 1927
rect 364 1825 398 1859
rect 364 1757 398 1791
rect 364 1689 398 1723
rect 364 1621 398 1655
rect 364 1553 398 1587
rect 364 1485 398 1519
rect 364 1417 398 1451
rect 364 1349 398 1383
rect 364 1281 398 1315
rect 364 1213 398 1247
rect 364 1145 398 1179
rect 364 1077 398 1111
rect 364 1009 398 1043
rect 364 941 398 975
rect 364 873 398 907
rect 364 805 398 839
rect 364 737 398 771
rect 364 669 398 703
rect 364 601 398 635
rect 364 533 398 567
rect 364 465 398 499
rect 364 397 398 431
rect 364 329 398 363
rect 364 261 398 295
rect 364 193 398 227
rect 364 125 398 159
rect 364 57 398 91
rect 452 1961 486 1995
rect 452 1893 486 1927
rect 452 1825 486 1859
rect 452 1757 486 1791
rect 452 1689 486 1723
rect 452 1621 486 1655
rect 452 1553 486 1587
rect 452 1485 486 1519
rect 452 1417 486 1451
rect 452 1349 486 1383
rect 452 1281 486 1315
rect 452 1213 486 1247
rect 452 1145 486 1179
rect 452 1077 486 1111
rect 452 1009 486 1043
rect 452 941 486 975
rect 452 873 486 907
rect 452 805 486 839
rect 452 737 486 771
rect 452 669 486 703
rect 452 601 486 635
rect 452 533 486 567
rect 452 465 486 499
rect 452 397 486 431
rect 452 329 486 363
rect 452 261 486 295
rect 452 193 486 227
rect 452 125 486 159
rect 452 57 486 91
rect 540 1961 574 1995
rect 540 1893 574 1927
rect 540 1825 574 1859
rect 540 1757 574 1791
rect 540 1689 574 1723
rect 540 1621 574 1655
rect 540 1553 574 1587
rect 540 1485 574 1519
rect 540 1417 574 1451
rect 540 1349 574 1383
rect 540 1281 574 1315
rect 540 1213 574 1247
rect 540 1145 574 1179
rect 540 1077 574 1111
rect 540 1009 574 1043
rect 540 941 574 975
rect 540 873 574 907
rect 540 805 574 839
rect 540 737 574 771
rect 540 669 574 703
rect 540 601 574 635
rect 540 533 574 567
rect 540 465 574 499
rect 540 397 574 431
rect 540 329 574 363
rect 540 261 574 295
rect 540 193 574 227
rect 540 125 574 159
rect 540 57 574 91
rect 628 1961 662 1995
rect 628 1893 662 1927
rect 628 1825 662 1859
rect 628 1757 662 1791
rect 628 1689 662 1723
rect 628 1621 662 1655
rect 628 1553 662 1587
rect 628 1485 662 1519
rect 628 1417 662 1451
rect 628 1349 662 1383
rect 628 1281 662 1315
rect 628 1213 662 1247
rect 628 1145 662 1179
rect 628 1077 662 1111
rect 628 1009 662 1043
rect 628 941 662 975
rect 628 873 662 907
rect 628 805 662 839
rect 628 737 662 771
rect 628 669 662 703
rect 628 601 662 635
rect 628 533 662 567
rect 628 465 662 499
rect 628 397 662 431
rect 628 329 662 363
rect 628 261 662 295
rect 628 193 662 227
rect 628 125 662 159
rect 628 57 662 91
rect 716 1961 750 1995
rect 716 1893 750 1927
rect 716 1825 750 1859
rect 716 1757 750 1791
rect 716 1689 750 1723
rect 716 1621 750 1655
rect 716 1553 750 1587
rect 716 1485 750 1519
rect 716 1417 750 1451
rect 716 1349 750 1383
rect 716 1281 750 1315
rect 716 1213 750 1247
rect 716 1145 750 1179
rect 716 1077 750 1111
rect 716 1009 750 1043
rect 716 941 750 975
rect 716 873 750 907
rect 716 805 750 839
rect 716 737 750 771
rect 716 669 750 703
rect 716 601 750 635
rect 716 533 750 567
rect 716 465 750 499
rect 716 397 750 431
rect 716 329 750 363
rect 716 261 750 295
rect 716 193 750 227
rect 716 125 750 159
rect 716 57 750 91
rect 804 1961 838 1995
rect 804 1893 838 1927
rect 804 1825 838 1859
rect 804 1757 838 1791
rect 804 1689 838 1723
rect 804 1621 838 1655
rect 804 1553 838 1587
rect 804 1485 838 1519
rect 804 1417 838 1451
rect 804 1349 838 1383
rect 804 1281 838 1315
rect 804 1213 838 1247
rect 804 1145 838 1179
rect 804 1077 838 1111
rect 804 1009 838 1043
rect 804 941 838 975
rect 804 873 838 907
rect 804 805 838 839
rect 804 737 838 771
rect 804 669 838 703
rect 804 601 838 635
rect 804 533 838 567
rect 804 465 838 499
rect 804 397 838 431
rect 804 329 838 363
rect 804 261 838 295
rect 804 193 838 227
rect 804 125 838 159
rect 804 57 838 91
rect 892 1961 926 1995
rect 892 1893 926 1927
rect 892 1825 926 1859
rect 892 1757 926 1791
rect 892 1689 926 1723
rect 892 1621 926 1655
rect 892 1553 926 1587
rect 892 1485 926 1519
rect 892 1417 926 1451
rect 892 1349 926 1383
rect 892 1281 926 1315
rect 892 1213 926 1247
rect 892 1145 926 1179
rect 892 1077 926 1111
rect 892 1009 926 1043
rect 892 941 926 975
rect 892 873 926 907
rect 892 805 926 839
rect 892 737 926 771
rect 892 669 926 703
rect 892 601 926 635
rect 892 533 926 567
rect 892 465 926 499
rect 892 397 926 431
rect 892 329 926 363
rect 892 261 926 295
rect 892 193 926 227
rect 892 125 926 159
rect 892 57 926 91
rect 980 1961 1014 1995
rect 980 1893 1014 1927
rect 980 1825 1014 1859
rect 980 1757 1014 1791
rect 980 1689 1014 1723
rect 980 1621 1014 1655
rect 980 1553 1014 1587
rect 980 1485 1014 1519
rect 980 1417 1014 1451
rect 980 1349 1014 1383
rect 980 1281 1014 1315
rect 980 1213 1014 1247
rect 980 1145 1014 1179
rect 980 1077 1014 1111
rect 980 1009 1014 1043
rect 980 941 1014 975
rect 980 873 1014 907
rect 980 805 1014 839
rect 980 737 1014 771
rect 980 669 1014 703
rect 980 601 1014 635
rect 980 533 1014 567
rect 980 465 1014 499
rect 980 397 1014 431
rect 980 329 1014 363
rect 980 261 1014 295
rect 980 193 1014 227
rect 980 125 1014 159
rect 980 57 1014 91
rect 1068 1961 1102 1995
rect 1068 1893 1102 1927
rect 1068 1825 1102 1859
rect 1068 1757 1102 1791
rect 1068 1689 1102 1723
rect 1068 1621 1102 1655
rect 1068 1553 1102 1587
rect 1068 1485 1102 1519
rect 1068 1417 1102 1451
rect 1068 1349 1102 1383
rect 1068 1281 1102 1315
rect 1068 1213 1102 1247
rect 1068 1145 1102 1179
rect 1068 1077 1102 1111
rect 1068 1009 1102 1043
rect 1068 941 1102 975
rect 1068 873 1102 907
rect 1068 805 1102 839
rect 1068 737 1102 771
rect 1068 669 1102 703
rect 1068 601 1102 635
rect 1068 533 1102 567
rect 1068 465 1102 499
rect 1068 397 1102 431
rect 1068 329 1102 363
rect 1068 261 1102 295
rect 1068 193 1102 227
rect 1068 125 1102 159
rect 1068 57 1102 91
rect 1156 1961 1190 1995
rect 1156 1893 1190 1927
rect 1156 1825 1190 1859
rect 1156 1757 1190 1791
rect 1156 1689 1190 1723
rect 1156 1621 1190 1655
rect 1156 1553 1190 1587
rect 1156 1485 1190 1519
rect 1156 1417 1190 1451
rect 1156 1349 1190 1383
rect 1156 1281 1190 1315
rect 1156 1213 1190 1247
rect 1156 1145 1190 1179
rect 1156 1077 1190 1111
rect 1156 1009 1190 1043
rect 1156 941 1190 975
rect 1156 873 1190 907
rect 1156 805 1190 839
rect 1156 737 1190 771
rect 1156 669 1190 703
rect 1156 601 1190 635
rect 1156 533 1190 567
rect 1156 465 1190 499
rect 1156 397 1190 431
rect 1156 329 1190 363
rect 1156 261 1190 295
rect 1156 193 1190 227
rect 1156 125 1190 159
rect 1156 57 1190 91
rect 1244 1961 1278 1995
rect 1244 1893 1278 1927
rect 1244 1825 1278 1859
rect 1244 1757 1278 1791
rect 1244 1689 1278 1723
rect 1244 1621 1278 1655
rect 1244 1553 1278 1587
rect 1244 1485 1278 1519
rect 1244 1417 1278 1451
rect 1244 1349 1278 1383
rect 1244 1281 1278 1315
rect 1244 1213 1278 1247
rect 1244 1145 1278 1179
rect 1244 1077 1278 1111
rect 1244 1009 1278 1043
rect 1244 941 1278 975
rect 1244 873 1278 907
rect 1244 805 1278 839
rect 1244 737 1278 771
rect 1244 669 1278 703
rect 1244 601 1278 635
rect 1244 533 1278 567
rect 1244 465 1278 499
rect 1244 397 1278 431
rect 1244 329 1278 363
rect 1244 261 1278 295
rect 1244 193 1278 227
rect 1244 125 1278 159
rect 1244 57 1278 91
rect 1332 1961 1366 1995
rect 1332 1893 1366 1927
rect 1332 1825 1366 1859
rect 1332 1757 1366 1791
rect 1332 1689 1366 1723
rect 1332 1621 1366 1655
rect 1332 1553 1366 1587
rect 1332 1485 1366 1519
rect 1332 1417 1366 1451
rect 1332 1349 1366 1383
rect 1332 1281 1366 1315
rect 1332 1213 1366 1247
rect 1332 1145 1366 1179
rect 1332 1077 1366 1111
rect 1332 1009 1366 1043
rect 1332 941 1366 975
rect 1332 873 1366 907
rect 1332 805 1366 839
rect 1332 737 1366 771
rect 1332 669 1366 703
rect 1332 601 1366 635
rect 1332 533 1366 567
rect 1332 465 1366 499
rect 1332 397 1366 431
rect 1332 329 1366 363
rect 1332 261 1366 295
rect 1332 193 1366 227
rect 1332 125 1366 159
rect 1332 57 1366 91
rect 1420 1961 1454 1995
rect 1420 1893 1454 1927
rect 1420 1825 1454 1859
rect 1420 1757 1454 1791
rect 1420 1689 1454 1723
rect 1420 1621 1454 1655
rect 1420 1553 1454 1587
rect 1420 1485 1454 1519
rect 1420 1417 1454 1451
rect 1420 1349 1454 1383
rect 1420 1281 1454 1315
rect 1420 1213 1454 1247
rect 1420 1145 1454 1179
rect 1420 1077 1454 1111
rect 1420 1009 1454 1043
rect 1420 941 1454 975
rect 1420 873 1454 907
rect 1420 805 1454 839
rect 1420 737 1454 771
rect 1420 669 1454 703
rect 1420 601 1454 635
rect 1420 533 1454 567
rect 1420 465 1454 499
rect 1420 397 1454 431
rect 1420 329 1454 363
rect 1420 261 1454 295
rect 1420 193 1454 227
rect 1420 125 1454 159
rect 1420 57 1454 91
rect 1508 1961 1542 1995
rect 1508 1893 1542 1927
rect 1508 1825 1542 1859
rect 1508 1757 1542 1791
rect 1508 1689 1542 1723
rect 1508 1621 1542 1655
rect 1508 1553 1542 1587
rect 1508 1485 1542 1519
rect 1508 1417 1542 1451
rect 1508 1349 1542 1383
rect 1508 1281 1542 1315
rect 1508 1213 1542 1247
rect 1508 1145 1542 1179
rect 1508 1077 1542 1111
rect 1508 1009 1542 1043
rect 1508 941 1542 975
rect 1508 873 1542 907
rect 1508 805 1542 839
rect 1508 737 1542 771
rect 1508 669 1542 703
rect 1508 601 1542 635
rect 1508 533 1542 567
rect 1508 465 1542 499
rect 1508 397 1542 431
rect 1508 329 1542 363
rect 1508 261 1542 295
rect 1508 193 1542 227
rect 1508 125 1542 159
rect 1508 57 1542 91
rect 1596 1961 1630 1995
rect 1596 1893 1630 1927
rect 1596 1825 1630 1859
rect 1596 1757 1630 1791
rect 1596 1689 1630 1723
rect 1596 1621 1630 1655
rect 1596 1553 1630 1587
rect 1596 1485 1630 1519
rect 1596 1417 1630 1451
rect 1596 1349 1630 1383
rect 1596 1281 1630 1315
rect 1596 1213 1630 1247
rect 1596 1145 1630 1179
rect 1596 1077 1630 1111
rect 1596 1009 1630 1043
rect 1596 941 1630 975
rect 1596 873 1630 907
rect 1596 805 1630 839
rect 1596 737 1630 771
rect 1596 669 1630 703
rect 1596 601 1630 635
rect 1596 533 1630 567
rect 1596 465 1630 499
rect 1596 397 1630 431
rect 1596 329 1630 363
rect 1596 261 1630 295
rect 1596 193 1630 227
rect 1596 125 1630 159
rect 1596 57 1630 91
rect 1684 1961 1718 1995
rect 1684 1893 1718 1927
rect 1684 1825 1718 1859
rect 1684 1757 1718 1791
rect 1684 1689 1718 1723
rect 1684 1621 1718 1655
rect 1684 1553 1718 1587
rect 1684 1485 1718 1519
rect 1684 1417 1718 1451
rect 1684 1349 1718 1383
rect 1684 1281 1718 1315
rect 1684 1213 1718 1247
rect 1684 1145 1718 1179
rect 1684 1077 1718 1111
rect 1684 1009 1718 1043
rect 1684 941 1718 975
rect 1684 873 1718 907
rect 1684 805 1718 839
rect 1684 737 1718 771
rect 1684 669 1718 703
rect 1684 601 1718 635
rect 1684 533 1718 567
rect 1684 465 1718 499
rect 1684 397 1718 431
rect 1684 329 1718 363
rect 1684 261 1718 295
rect 1684 193 1718 227
rect 1684 125 1718 159
rect 1684 57 1718 91
rect 1772 1961 1806 1995
rect 1772 1893 1806 1927
rect 1772 1825 1806 1859
rect 1772 1757 1806 1791
rect 1772 1689 1806 1723
rect 1772 1621 1806 1655
rect 1772 1553 1806 1587
rect 1772 1485 1806 1519
rect 1772 1417 1806 1451
rect 1772 1349 1806 1383
rect 1772 1281 1806 1315
rect 1772 1213 1806 1247
rect 1772 1145 1806 1179
rect 1772 1077 1806 1111
rect 1772 1009 1806 1043
rect 1772 941 1806 975
rect 1772 873 1806 907
rect 1772 805 1806 839
rect 1772 737 1806 771
rect 1772 669 1806 703
rect 1772 601 1806 635
rect 1772 533 1806 567
rect 1772 465 1806 499
rect 1772 397 1806 431
rect 1772 329 1806 363
rect 1772 261 1806 295
rect 1772 193 1806 227
rect 1772 125 1806 159
rect 1772 57 1806 91
rect 1860 1961 1894 1995
rect 1860 1893 1894 1927
rect 1860 1825 1894 1859
rect 1860 1757 1894 1791
rect 1860 1689 1894 1723
rect 1860 1621 1894 1655
rect 1860 1553 1894 1587
rect 1860 1485 1894 1519
rect 1860 1417 1894 1451
rect 1860 1349 1894 1383
rect 1860 1281 1894 1315
rect 1860 1213 1894 1247
rect 1860 1145 1894 1179
rect 1860 1077 1894 1111
rect 1860 1009 1894 1043
rect 1860 941 1894 975
rect 1860 873 1894 907
rect 1860 805 1894 839
rect 1860 737 1894 771
rect 1860 669 1894 703
rect 1860 601 1894 635
rect 1860 533 1894 567
rect 1860 465 1894 499
rect 1860 397 1894 431
rect 1860 329 1894 363
rect 1860 261 1894 295
rect 1860 193 1894 227
rect 1860 125 1894 159
rect 1860 57 1894 91
rect 1948 1961 1982 1995
rect 1948 1893 1982 1927
rect 1948 1825 1982 1859
rect 1948 1757 1982 1791
rect 1948 1689 1982 1723
rect 1948 1621 1982 1655
rect 1948 1553 1982 1587
rect 1948 1485 1982 1519
rect 1948 1417 1982 1451
rect 1948 1349 1982 1383
rect 1948 1281 1982 1315
rect 1948 1213 1982 1247
rect 1948 1145 1982 1179
rect 1948 1077 1982 1111
rect 1948 1009 1982 1043
rect 1948 941 1982 975
rect 1948 873 1982 907
rect 1948 805 1982 839
rect 1948 737 1982 771
rect 1948 669 1982 703
rect 1948 601 1982 635
rect 1948 533 1982 567
rect 1948 465 1982 499
rect 1948 397 1982 431
rect 1948 329 1982 363
rect 1948 261 1982 295
rect 1948 193 1982 227
rect 1948 125 1982 159
rect 1948 57 1982 91
rect 2036 1961 2070 1995
rect 2036 1893 2070 1927
rect 2036 1825 2070 1859
rect 2036 1757 2070 1791
rect 2036 1689 2070 1723
rect 2036 1621 2070 1655
rect 2036 1553 2070 1587
rect 2036 1485 2070 1519
rect 2036 1417 2070 1451
rect 2036 1349 2070 1383
rect 2036 1281 2070 1315
rect 2036 1213 2070 1247
rect 2036 1145 2070 1179
rect 2036 1077 2070 1111
rect 2036 1009 2070 1043
rect 2036 941 2070 975
rect 2036 873 2070 907
rect 2036 805 2070 839
rect 2036 737 2070 771
rect 2036 669 2070 703
rect 2036 601 2070 635
rect 2036 533 2070 567
rect 2036 465 2070 499
rect 2036 397 2070 431
rect 2036 329 2070 363
rect 2036 261 2070 295
rect 2036 193 2070 227
rect 2036 125 2070 159
rect 2036 57 2070 91
rect 2124 1961 2158 1995
rect 2124 1893 2158 1927
rect 2124 1825 2158 1859
rect 2124 1757 2158 1791
rect 2124 1689 2158 1723
rect 2124 1621 2158 1655
rect 2124 1553 2158 1587
rect 2124 1485 2158 1519
rect 2124 1417 2158 1451
rect 2124 1349 2158 1383
rect 2124 1281 2158 1315
rect 2124 1213 2158 1247
rect 2124 1145 2158 1179
rect 2124 1077 2158 1111
rect 2124 1009 2158 1043
rect 2124 941 2158 975
rect 2124 873 2158 907
rect 2124 805 2158 839
rect 2124 737 2158 771
rect 2124 669 2158 703
rect 2124 601 2158 635
rect 2124 533 2158 567
rect 2124 465 2158 499
rect 2124 397 2158 431
rect 2124 329 2158 363
rect 2124 261 2158 295
rect 2124 193 2158 227
rect 2124 125 2158 159
rect 2124 57 2158 91
rect 2212 1961 2246 1995
rect 2212 1893 2246 1927
rect 2212 1825 2246 1859
rect 2212 1757 2246 1791
rect 2212 1689 2246 1723
rect 2212 1621 2246 1655
rect 2212 1553 2246 1587
rect 2212 1485 2246 1519
rect 2212 1417 2246 1451
rect 2212 1349 2246 1383
rect 2212 1281 2246 1315
rect 2212 1213 2246 1247
rect 2212 1145 2246 1179
rect 2212 1077 2246 1111
rect 2212 1009 2246 1043
rect 2212 941 2246 975
rect 2212 873 2246 907
rect 2212 805 2246 839
rect 2212 737 2246 771
rect 2212 669 2246 703
rect 2212 601 2246 635
rect 2212 533 2246 567
rect 2212 465 2246 499
rect 2212 397 2246 431
rect 2212 329 2246 363
rect 2212 261 2246 295
rect 2212 193 2246 227
rect 2212 125 2246 159
rect 2212 57 2246 91
rect 2300 1961 2334 1995
rect 2300 1893 2334 1927
rect 2300 1825 2334 1859
rect 2300 1757 2334 1791
rect 2300 1689 2334 1723
rect 2300 1621 2334 1655
rect 2300 1553 2334 1587
rect 2300 1485 2334 1519
rect 2300 1417 2334 1451
rect 2300 1349 2334 1383
rect 2300 1281 2334 1315
rect 2300 1213 2334 1247
rect 2300 1145 2334 1179
rect 2300 1077 2334 1111
rect 2300 1009 2334 1043
rect 2300 941 2334 975
rect 2300 873 2334 907
rect 2300 805 2334 839
rect 2300 737 2334 771
rect 2300 669 2334 703
rect 2300 601 2334 635
rect 2300 533 2334 567
rect 2300 465 2334 499
rect 2300 397 2334 431
rect 2300 329 2334 363
rect 2300 261 2334 295
rect 2300 193 2334 227
rect 2300 125 2334 159
rect 2300 57 2334 91
rect 2388 1961 2422 1995
rect 2388 1893 2422 1927
rect 2388 1825 2422 1859
rect 2388 1757 2422 1791
rect 2388 1689 2422 1723
rect 2388 1621 2422 1655
rect 2388 1553 2422 1587
rect 2388 1485 2422 1519
rect 2388 1417 2422 1451
rect 2388 1349 2422 1383
rect 2388 1281 2422 1315
rect 2388 1213 2422 1247
rect 2388 1145 2422 1179
rect 2388 1077 2422 1111
rect 2388 1009 2422 1043
rect 2388 941 2422 975
rect 2388 873 2422 907
rect 2388 805 2422 839
rect 2388 737 2422 771
rect 2388 669 2422 703
rect 2388 601 2422 635
rect 2388 533 2422 567
rect 2388 465 2422 499
rect 2388 397 2422 431
rect 2388 329 2422 363
rect 2388 261 2422 295
rect 2388 193 2422 227
rect 2388 125 2422 159
rect 2388 57 2422 91
rect 2476 1961 2510 1995
rect 2476 1893 2510 1927
rect 2476 1825 2510 1859
rect 2476 1757 2510 1791
rect 2476 1689 2510 1723
rect 2476 1621 2510 1655
rect 2476 1553 2510 1587
rect 2476 1485 2510 1519
rect 2476 1417 2510 1451
rect 2476 1349 2510 1383
rect 2476 1281 2510 1315
rect 2476 1213 2510 1247
rect 2476 1145 2510 1179
rect 2476 1077 2510 1111
rect 2476 1009 2510 1043
rect 2476 941 2510 975
rect 2476 873 2510 907
rect 2476 805 2510 839
rect 2476 737 2510 771
rect 2476 669 2510 703
rect 2476 601 2510 635
rect 2476 533 2510 567
rect 2476 465 2510 499
rect 2476 397 2510 431
rect 2476 329 2510 363
rect 2476 261 2510 295
rect 2476 193 2510 227
rect 2476 125 2510 159
rect 2476 57 2510 91
rect 2564 1961 2598 1995
rect 2564 1893 2598 1927
rect 2564 1825 2598 1859
rect 2564 1757 2598 1791
rect 2564 1689 2598 1723
rect 2564 1621 2598 1655
rect 2564 1553 2598 1587
rect 2564 1485 2598 1519
rect 2564 1417 2598 1451
rect 2564 1349 2598 1383
rect 2564 1281 2598 1315
rect 2564 1213 2598 1247
rect 2564 1145 2598 1179
rect 2564 1077 2598 1111
rect 2564 1009 2598 1043
rect 2564 941 2598 975
rect 2564 873 2598 907
rect 2564 805 2598 839
rect 2564 737 2598 771
rect 2564 669 2598 703
rect 2564 601 2598 635
rect 2564 533 2598 567
rect 2564 465 2598 499
rect 2564 397 2598 431
rect 2564 329 2598 363
rect 2564 261 2598 295
rect 2564 193 2598 227
rect 2564 125 2598 159
rect 2564 57 2598 91
rect 2652 1961 2686 1995
rect 2652 1893 2686 1927
rect 2652 1825 2686 1859
rect 2652 1757 2686 1791
rect 2652 1689 2686 1723
rect 2652 1621 2686 1655
rect 2652 1553 2686 1587
rect 2652 1485 2686 1519
rect 2652 1417 2686 1451
rect 2652 1349 2686 1383
rect 2652 1281 2686 1315
rect 2652 1213 2686 1247
rect 2652 1145 2686 1179
rect 2652 1077 2686 1111
rect 2652 1009 2686 1043
rect 2652 941 2686 975
rect 2652 873 2686 907
rect 2652 805 2686 839
rect 2652 737 2686 771
rect 2652 669 2686 703
rect 2652 601 2686 635
rect 2652 533 2686 567
rect 2652 465 2686 499
rect 2652 397 2686 431
rect 2652 329 2686 363
rect 2652 261 2686 295
rect 2652 193 2686 227
rect 2652 125 2686 159
rect 2652 57 2686 91
<< psubdiff >>
rect -399 2775 3195 2808
rect -399 2605 14 2775
rect 2768 2605 3195 2775
rect -399 2573 3195 2605
rect -399 1995 -178 2573
rect -399 57 -374 1995
rect -204 57 -178 1995
rect -399 -392 -178 57
rect 2974 1981 3195 2573
rect 2974 43 2999 1981
rect 3169 43 3195 1981
rect 2974 -392 3195 43
rect -399 -425 3195 -392
rect -399 -595 -85 -425
rect 2669 -557 3195 -425
rect 2669 -595 3194 -557
rect -399 -627 3194 -595
<< psubdiffcont >>
rect 14 2605 2768 2775
rect -374 57 -204 1995
rect 2999 43 3169 1981
rect -85 -595 2669 -425
<< poly >>
rect 58 2026 88 2052
rect 146 2026 176 2052
rect 234 2026 264 2052
rect 322 2026 352 2052
rect 410 2026 440 2052
rect 498 2026 528 2052
rect 586 2026 616 2052
rect 674 2026 704 2052
rect 762 2026 792 2052
rect 850 2026 880 2052
rect 938 2026 968 2052
rect 1026 2026 1056 2052
rect 1114 2026 1144 2052
rect 1202 2026 1232 2052
rect 1290 2026 1320 2052
rect 1378 2026 1408 2052
rect 1466 2026 1496 2052
rect 1554 2026 1584 2052
rect 1642 2026 1672 2052
rect 1730 2026 1760 2052
rect 1818 2026 1848 2052
rect 1906 2026 1936 2052
rect 1994 2026 2024 2052
rect 2082 2026 2112 2052
rect 2170 2026 2200 2052
rect 2258 2026 2288 2052
rect 2346 2026 2376 2052
rect 2434 2026 2464 2052
rect 2522 2026 2552 2052
rect 2610 2026 2640 2052
rect 58 22 88 26
rect 146 0 176 26
rect 58 -29 176 0
rect 58 -63 100 -29
rect 134 -63 176 -29
rect 58 -92 176 -63
rect 234 0 264 26
rect 322 0 352 26
rect 234 -29 352 0
rect 234 -63 276 -29
rect 310 -63 352 -29
rect 234 -92 352 -63
rect 410 0 440 26
rect 498 0 528 26
rect 410 -29 528 0
rect 410 -63 452 -29
rect 486 -63 528 -29
rect 410 -92 528 -63
rect 586 0 616 26
rect 674 0 704 26
rect 586 -29 704 0
rect 586 -63 628 -29
rect 662 -63 704 -29
rect 586 -92 704 -63
rect 762 0 792 26
rect 850 0 880 26
rect 762 -193 880 0
rect 938 0 968 26
rect 1026 0 1056 26
rect 938 -29 1056 0
rect 938 -63 980 -29
rect 1014 -63 1056 -29
rect 938 -92 1056 -63
rect 1114 0 1144 26
rect 1202 0 1232 26
rect 762 -227 804 -193
rect 838 -227 880 -193
rect 762 -256 880 -227
rect 1114 -193 1232 0
rect 1290 0 1320 26
rect 1378 0 1408 26
rect 1290 -29 1408 0
rect 1290 -63 1332 -29
rect 1366 -63 1408 -29
rect 1290 -92 1408 -63
rect 1466 0 1496 26
rect 1554 0 1584 26
rect 1114 -227 1156 -193
rect 1190 -227 1232 -193
rect 1114 -256 1232 -227
rect 1466 -193 1584 0
rect 1642 0 1672 26
rect 1730 0 1760 26
rect 1642 -29 1760 0
rect 1642 -63 1684 -29
rect 1718 -63 1760 -29
rect 1642 -92 1760 -63
rect 1818 0 1848 26
rect 1906 0 1936 26
rect 1466 -227 1508 -193
rect 1542 -227 1584 -193
rect 1466 -256 1584 -227
rect 1818 -193 1936 0
rect 1994 0 2024 26
rect 2082 0 2112 26
rect 1994 -29 2112 0
rect 1994 -63 2036 -29
rect 2070 -63 2112 -29
rect 1994 -92 2112 -63
rect 2170 0 2200 26
rect 2258 0 2288 26
rect 1818 -227 1860 -193
rect 1894 -227 1936 -193
rect 1818 -256 1936 -227
rect 2170 -193 2288 0
rect 2346 0 2376 26
rect 2434 0 2464 26
rect 2346 -29 2464 0
rect 2346 -63 2388 -29
rect 2422 -63 2464 -29
rect 2346 -92 2464 -63
rect 2522 0 2552 26
rect 2610 0 2640 26
rect 2522 -29 2640 0
rect 2522 -63 2564 -29
rect 2598 -63 2640 -29
rect 2522 -92 2640 -63
rect 2170 -227 2212 -193
rect 2246 -227 2288 -193
rect 2170 -256 2288 -227
<< polycont >>
rect 100 -63 134 -29
rect 276 -63 310 -29
rect 452 -63 486 -29
rect 628 -63 662 -29
rect 980 -63 1014 -29
rect 804 -227 838 -193
rect 1332 -63 1366 -29
rect 1156 -227 1190 -193
rect 1684 -63 1718 -29
rect 1508 -227 1542 -193
rect 2036 -63 2070 -29
rect 1860 -227 1894 -193
rect 2388 -63 2422 -29
rect 2564 -63 2598 -29
rect 2212 -227 2246 -193
<< locali >>
rect -399 2775 3195 2808
rect -399 2605 14 2775
rect 2768 2605 3195 2775
rect -399 2573 3195 2605
rect -399 1995 -178 2573
rect 609 2378 681 2396
rect 609 2344 628 2378
rect 662 2344 681 2378
rect 609 2326 681 2344
rect 961 2378 1033 2396
rect 961 2344 980 2378
rect 1014 2344 1033 2378
rect 961 2326 1033 2344
rect 1313 2378 1385 2396
rect 1313 2344 1332 2378
rect 1366 2344 1385 2378
rect 1313 2326 1385 2344
rect 1665 2378 1737 2396
rect 1665 2344 1684 2378
rect 1718 2344 1737 2378
rect 1665 2326 1737 2344
rect 2017 2378 2089 2396
rect 2017 2344 2036 2378
rect 2070 2344 2089 2378
rect 2017 2326 2089 2344
rect 81 2273 153 2291
rect 81 2239 100 2273
rect 134 2239 153 2273
rect 81 2221 153 2239
rect 257 2273 329 2291
rect 257 2239 276 2273
rect 310 2239 329 2273
rect 257 2221 329 2239
rect 433 2273 505 2291
rect 433 2239 452 2273
rect 486 2239 505 2273
rect 433 2221 505 2239
rect -7 2169 65 2187
rect -7 2135 12 2169
rect 46 2135 65 2169
rect -7 2117 65 2135
rect -399 57 -374 1995
rect -204 57 -178 1995
rect -399 -392 -178 57
rect 12 1995 46 2117
rect 12 1927 46 1945
rect 12 1859 46 1873
rect 12 1791 46 1801
rect 12 1723 46 1729
rect 12 1655 46 1657
rect 12 1619 46 1621
rect 12 1547 46 1553
rect 12 1475 46 1485
rect 12 1403 46 1417
rect 12 1331 46 1349
rect 12 1259 46 1281
rect 12 1187 46 1213
rect 12 1115 46 1145
rect 12 1043 46 1077
rect 12 975 46 1009
rect 12 907 46 937
rect 12 839 46 865
rect 12 771 46 793
rect 12 703 46 721
rect 12 635 46 649
rect 12 567 46 577
rect 12 499 46 505
rect 12 431 46 433
rect 12 395 46 397
rect 12 323 46 329
rect 12 251 46 261
rect 12 179 46 193
rect 12 107 46 125
rect 12 22 46 57
rect 100 1995 134 2221
rect 169 2169 241 2187
rect 169 2135 188 2169
rect 222 2135 241 2169
rect 169 2117 241 2135
rect 100 1927 134 1945
rect 100 1859 134 1873
rect 100 1791 134 1801
rect 100 1723 134 1729
rect 100 1655 134 1657
rect 100 1619 134 1621
rect 100 1547 134 1553
rect 100 1475 134 1485
rect 100 1403 134 1417
rect 100 1331 134 1349
rect 100 1259 134 1281
rect 100 1187 134 1213
rect 100 1115 134 1145
rect 100 1043 134 1077
rect 100 975 134 1009
rect 100 907 134 937
rect 100 839 134 865
rect 100 771 134 793
rect 100 703 134 721
rect 100 635 134 649
rect 100 567 134 577
rect 100 499 134 505
rect 100 431 134 433
rect 100 395 134 397
rect 100 323 134 329
rect 100 251 134 261
rect 100 179 134 193
rect 100 107 134 125
rect 100 22 134 57
rect 188 1995 222 2117
rect 188 1927 222 1945
rect 188 1859 222 1873
rect 188 1791 222 1801
rect 188 1723 222 1729
rect 188 1655 222 1657
rect 188 1619 222 1621
rect 188 1547 222 1553
rect 188 1475 222 1485
rect 188 1403 222 1417
rect 188 1331 222 1349
rect 188 1259 222 1281
rect 188 1187 222 1213
rect 188 1115 222 1145
rect 188 1043 222 1077
rect 188 975 222 1009
rect 188 907 222 937
rect 188 839 222 865
rect 188 771 222 793
rect 188 703 222 721
rect 188 635 222 649
rect 188 567 222 577
rect 188 499 222 505
rect 188 431 222 433
rect 188 395 222 397
rect 188 323 222 329
rect 188 251 222 261
rect 188 179 222 193
rect 188 107 222 125
rect 188 22 222 57
rect 276 1995 310 2221
rect 345 2169 417 2187
rect 345 2135 364 2169
rect 398 2135 417 2169
rect 345 2117 417 2135
rect 276 1927 310 1945
rect 276 1859 310 1873
rect 276 1791 310 1801
rect 276 1723 310 1729
rect 276 1655 310 1657
rect 276 1619 310 1621
rect 276 1547 310 1553
rect 276 1475 310 1485
rect 276 1403 310 1417
rect 276 1331 310 1349
rect 276 1259 310 1281
rect 276 1187 310 1213
rect 276 1115 310 1145
rect 276 1043 310 1077
rect 276 975 310 1009
rect 276 907 310 937
rect 276 839 310 865
rect 276 771 310 793
rect 276 703 310 721
rect 276 635 310 649
rect 276 567 310 577
rect 276 499 310 505
rect 276 431 310 433
rect 276 395 310 397
rect 276 323 310 329
rect 276 251 310 261
rect 276 179 310 193
rect 276 107 310 125
rect 276 22 310 57
rect 364 1995 398 2117
rect 364 1927 398 1945
rect 364 1859 398 1873
rect 364 1791 398 1801
rect 364 1723 398 1729
rect 364 1655 398 1657
rect 364 1619 398 1621
rect 364 1547 398 1553
rect 364 1475 398 1485
rect 364 1403 398 1417
rect 364 1331 398 1349
rect 364 1259 398 1281
rect 364 1187 398 1213
rect 364 1115 398 1145
rect 364 1043 398 1077
rect 364 975 398 1009
rect 364 907 398 937
rect 364 839 398 865
rect 364 771 398 793
rect 364 703 398 721
rect 364 635 398 649
rect 364 567 398 577
rect 364 499 398 505
rect 364 431 398 433
rect 364 395 398 397
rect 364 323 398 329
rect 364 251 398 261
rect 364 179 398 193
rect 364 107 398 125
rect 364 22 398 57
rect 452 1995 486 2221
rect 521 2169 593 2187
rect 521 2135 540 2169
rect 574 2135 593 2169
rect 521 2117 593 2135
rect 452 1927 486 1945
rect 452 1859 486 1873
rect 452 1791 486 1801
rect 452 1723 486 1729
rect 452 1655 486 1657
rect 452 1619 486 1621
rect 452 1547 486 1553
rect 452 1475 486 1485
rect 452 1403 486 1417
rect 452 1331 486 1349
rect 452 1259 486 1281
rect 452 1187 486 1213
rect 452 1115 486 1145
rect 452 1043 486 1077
rect 452 975 486 1009
rect 452 907 486 937
rect 452 839 486 865
rect 452 771 486 793
rect 452 703 486 721
rect 452 635 486 649
rect 452 567 486 577
rect 452 499 486 505
rect 452 431 486 433
rect 452 395 486 397
rect 452 323 486 329
rect 452 251 486 261
rect 452 179 486 193
rect 452 107 486 125
rect 452 22 486 57
rect 540 1995 574 2117
rect 540 1927 574 1945
rect 540 1859 574 1873
rect 540 1791 574 1801
rect 540 1723 574 1729
rect 540 1655 574 1657
rect 540 1619 574 1621
rect 540 1547 574 1553
rect 540 1475 574 1485
rect 540 1403 574 1417
rect 540 1331 574 1349
rect 540 1259 574 1281
rect 540 1187 574 1213
rect 540 1115 574 1145
rect 540 1043 574 1077
rect 540 975 574 1009
rect 540 907 574 937
rect 540 839 574 865
rect 540 771 574 793
rect 540 703 574 721
rect 540 635 574 649
rect 540 567 574 577
rect 540 499 574 505
rect 540 431 574 433
rect 540 395 574 397
rect 540 323 574 329
rect 540 251 574 261
rect 540 179 574 193
rect 540 107 574 125
rect 540 22 574 57
rect 628 1995 662 2326
rect 785 2273 857 2291
rect 785 2239 804 2273
rect 838 2239 857 2273
rect 785 2221 857 2239
rect 697 2169 769 2187
rect 697 2135 716 2169
rect 750 2135 769 2169
rect 697 2117 769 2135
rect 628 1927 662 1945
rect 628 1859 662 1873
rect 628 1791 662 1801
rect 628 1723 662 1729
rect 628 1655 662 1657
rect 628 1619 662 1621
rect 628 1547 662 1553
rect 628 1475 662 1485
rect 628 1403 662 1417
rect 628 1331 662 1349
rect 628 1259 662 1281
rect 628 1187 662 1213
rect 628 1115 662 1145
rect 628 1043 662 1077
rect 628 975 662 1009
rect 628 907 662 937
rect 628 839 662 865
rect 628 771 662 793
rect 628 703 662 721
rect 628 635 662 649
rect 628 567 662 577
rect 628 499 662 505
rect 628 431 662 433
rect 628 395 662 397
rect 628 323 662 329
rect 628 251 662 261
rect 628 179 662 193
rect 628 107 662 125
rect 628 22 662 57
rect 716 1995 750 2117
rect 716 1927 750 1945
rect 716 1859 750 1873
rect 716 1791 750 1801
rect 716 1723 750 1729
rect 716 1655 750 1657
rect 716 1619 750 1621
rect 716 1547 750 1553
rect 716 1475 750 1485
rect 716 1403 750 1417
rect 716 1331 750 1349
rect 716 1259 750 1281
rect 716 1187 750 1213
rect 716 1115 750 1145
rect 716 1043 750 1077
rect 716 975 750 1009
rect 716 907 750 937
rect 716 839 750 865
rect 716 771 750 793
rect 716 703 750 721
rect 716 635 750 649
rect 716 567 750 577
rect 716 499 750 505
rect 716 431 750 433
rect 716 395 750 397
rect 716 323 750 329
rect 716 251 750 261
rect 716 179 750 193
rect 716 107 750 125
rect 716 22 750 57
rect 804 1995 838 2221
rect 873 2169 945 2187
rect 873 2135 892 2169
rect 926 2135 945 2169
rect 873 2117 945 2135
rect 804 1927 838 1945
rect 804 1859 838 1873
rect 804 1791 838 1801
rect 804 1723 838 1729
rect 804 1655 838 1657
rect 804 1619 838 1621
rect 804 1547 838 1553
rect 804 1475 838 1485
rect 804 1403 838 1417
rect 804 1331 838 1349
rect 804 1259 838 1281
rect 804 1187 838 1213
rect 804 1115 838 1145
rect 804 1043 838 1077
rect 804 975 838 1009
rect 804 907 838 937
rect 804 839 838 865
rect 804 771 838 793
rect 804 703 838 721
rect 804 635 838 649
rect 804 567 838 577
rect 804 499 838 505
rect 804 431 838 433
rect 804 395 838 397
rect 804 323 838 329
rect 804 251 838 261
rect 804 179 838 193
rect 804 107 838 125
rect 804 22 838 57
rect 892 1995 926 2117
rect 892 1927 926 1945
rect 892 1859 926 1873
rect 892 1791 926 1801
rect 892 1723 926 1729
rect 892 1655 926 1657
rect 892 1619 926 1621
rect 892 1547 926 1553
rect 892 1475 926 1485
rect 892 1403 926 1417
rect 892 1331 926 1349
rect 892 1259 926 1281
rect 892 1187 926 1213
rect 892 1115 926 1145
rect 892 1043 926 1077
rect 892 975 926 1009
rect 892 907 926 937
rect 892 839 926 865
rect 892 771 926 793
rect 892 703 926 721
rect 892 635 926 649
rect 892 567 926 577
rect 892 499 926 505
rect 892 431 926 433
rect 892 395 926 397
rect 892 323 926 329
rect 892 251 926 261
rect 892 179 926 193
rect 892 107 926 125
rect 892 22 926 57
rect 980 1995 1014 2326
rect 1137 2273 1209 2291
rect 1137 2239 1156 2273
rect 1190 2239 1209 2273
rect 1137 2221 1209 2239
rect 1049 2169 1121 2187
rect 1049 2135 1068 2169
rect 1102 2135 1121 2169
rect 1049 2117 1121 2135
rect 980 1927 1014 1945
rect 980 1859 1014 1873
rect 980 1791 1014 1801
rect 980 1723 1014 1729
rect 980 1655 1014 1657
rect 980 1619 1014 1621
rect 980 1547 1014 1553
rect 980 1475 1014 1485
rect 980 1403 1014 1417
rect 980 1331 1014 1349
rect 980 1259 1014 1281
rect 980 1187 1014 1213
rect 980 1115 1014 1145
rect 980 1043 1014 1077
rect 980 975 1014 1009
rect 980 907 1014 937
rect 980 839 1014 865
rect 980 771 1014 793
rect 980 703 1014 721
rect 980 635 1014 649
rect 980 567 1014 577
rect 980 499 1014 505
rect 980 431 1014 433
rect 980 395 1014 397
rect 980 323 1014 329
rect 980 251 1014 261
rect 980 179 1014 193
rect 980 107 1014 125
rect 980 22 1014 57
rect 1068 1995 1102 2117
rect 1068 1927 1102 1945
rect 1068 1859 1102 1873
rect 1068 1791 1102 1801
rect 1068 1723 1102 1729
rect 1068 1655 1102 1657
rect 1068 1619 1102 1621
rect 1068 1547 1102 1553
rect 1068 1475 1102 1485
rect 1068 1403 1102 1417
rect 1068 1331 1102 1349
rect 1068 1259 1102 1281
rect 1068 1187 1102 1213
rect 1068 1115 1102 1145
rect 1068 1043 1102 1077
rect 1068 975 1102 1009
rect 1068 907 1102 937
rect 1068 839 1102 865
rect 1068 771 1102 793
rect 1068 703 1102 721
rect 1068 635 1102 649
rect 1068 567 1102 577
rect 1068 499 1102 505
rect 1068 431 1102 433
rect 1068 395 1102 397
rect 1068 323 1102 329
rect 1068 251 1102 261
rect 1068 179 1102 193
rect 1068 107 1102 125
rect 1068 22 1102 57
rect 1156 1995 1190 2221
rect 1225 2169 1297 2187
rect 1225 2135 1244 2169
rect 1278 2135 1297 2169
rect 1225 2117 1297 2135
rect 1156 1927 1190 1945
rect 1156 1859 1190 1873
rect 1156 1791 1190 1801
rect 1156 1723 1190 1729
rect 1156 1655 1190 1657
rect 1156 1619 1190 1621
rect 1156 1547 1190 1553
rect 1156 1475 1190 1485
rect 1156 1403 1190 1417
rect 1156 1331 1190 1349
rect 1156 1259 1190 1281
rect 1156 1187 1190 1213
rect 1156 1115 1190 1145
rect 1156 1043 1190 1077
rect 1156 975 1190 1009
rect 1156 907 1190 937
rect 1156 839 1190 865
rect 1156 771 1190 793
rect 1156 703 1190 721
rect 1156 635 1190 649
rect 1156 567 1190 577
rect 1156 499 1190 505
rect 1156 431 1190 433
rect 1156 395 1190 397
rect 1156 323 1190 329
rect 1156 251 1190 261
rect 1156 179 1190 193
rect 1156 107 1190 125
rect 1156 22 1190 57
rect 1244 1995 1278 2117
rect 1244 1927 1278 1945
rect 1244 1859 1278 1873
rect 1244 1791 1278 1801
rect 1244 1723 1278 1729
rect 1244 1655 1278 1657
rect 1244 1619 1278 1621
rect 1244 1547 1278 1553
rect 1244 1475 1278 1485
rect 1244 1403 1278 1417
rect 1244 1331 1278 1349
rect 1244 1259 1278 1281
rect 1244 1187 1278 1213
rect 1244 1115 1278 1145
rect 1244 1043 1278 1077
rect 1244 975 1278 1009
rect 1244 907 1278 937
rect 1244 839 1278 865
rect 1244 771 1278 793
rect 1244 703 1278 721
rect 1244 635 1278 649
rect 1244 567 1278 577
rect 1244 499 1278 505
rect 1244 431 1278 433
rect 1244 395 1278 397
rect 1244 323 1278 329
rect 1244 251 1278 261
rect 1244 179 1278 193
rect 1244 107 1278 125
rect 1244 22 1278 57
rect 1332 1995 1366 2326
rect 1489 2273 1561 2291
rect 1489 2239 1508 2273
rect 1542 2239 1561 2273
rect 1489 2221 1561 2239
rect 1401 2169 1473 2187
rect 1401 2135 1420 2169
rect 1454 2135 1473 2169
rect 1401 2117 1473 2135
rect 1332 1927 1366 1945
rect 1332 1859 1366 1873
rect 1332 1791 1366 1801
rect 1332 1723 1366 1729
rect 1332 1655 1366 1657
rect 1332 1619 1366 1621
rect 1332 1547 1366 1553
rect 1332 1475 1366 1485
rect 1332 1403 1366 1417
rect 1332 1331 1366 1349
rect 1332 1259 1366 1281
rect 1332 1187 1366 1213
rect 1332 1115 1366 1145
rect 1332 1043 1366 1077
rect 1332 975 1366 1009
rect 1332 907 1366 937
rect 1332 839 1366 865
rect 1332 771 1366 793
rect 1332 703 1366 721
rect 1332 635 1366 649
rect 1332 567 1366 577
rect 1332 499 1366 505
rect 1332 431 1366 433
rect 1332 395 1366 397
rect 1332 323 1366 329
rect 1332 251 1366 261
rect 1332 179 1366 193
rect 1332 107 1366 125
rect 1332 22 1366 57
rect 1420 1995 1454 2117
rect 1420 1927 1454 1945
rect 1420 1859 1454 1873
rect 1420 1791 1454 1801
rect 1420 1723 1454 1729
rect 1420 1655 1454 1657
rect 1420 1619 1454 1621
rect 1420 1547 1454 1553
rect 1420 1475 1454 1485
rect 1420 1403 1454 1417
rect 1420 1331 1454 1349
rect 1420 1259 1454 1281
rect 1420 1187 1454 1213
rect 1420 1115 1454 1145
rect 1420 1043 1454 1077
rect 1420 975 1454 1009
rect 1420 907 1454 937
rect 1420 839 1454 865
rect 1420 771 1454 793
rect 1420 703 1454 721
rect 1420 635 1454 649
rect 1420 567 1454 577
rect 1420 499 1454 505
rect 1420 431 1454 433
rect 1420 395 1454 397
rect 1420 323 1454 329
rect 1420 251 1454 261
rect 1420 179 1454 193
rect 1420 107 1454 125
rect 1420 22 1454 57
rect 1508 1995 1542 2221
rect 1577 2169 1649 2187
rect 1577 2135 1596 2169
rect 1630 2135 1649 2169
rect 1577 2117 1649 2135
rect 1508 1927 1542 1945
rect 1508 1859 1542 1873
rect 1508 1791 1542 1801
rect 1508 1723 1542 1729
rect 1508 1655 1542 1657
rect 1508 1619 1542 1621
rect 1508 1547 1542 1553
rect 1508 1475 1542 1485
rect 1508 1403 1542 1417
rect 1508 1331 1542 1349
rect 1508 1259 1542 1281
rect 1508 1187 1542 1213
rect 1508 1115 1542 1145
rect 1508 1043 1542 1077
rect 1508 975 1542 1009
rect 1508 907 1542 937
rect 1508 839 1542 865
rect 1508 771 1542 793
rect 1508 703 1542 721
rect 1508 635 1542 649
rect 1508 567 1542 577
rect 1508 499 1542 505
rect 1508 431 1542 433
rect 1508 395 1542 397
rect 1508 323 1542 329
rect 1508 251 1542 261
rect 1508 179 1542 193
rect 1508 107 1542 125
rect 1508 22 1542 57
rect 1596 1995 1630 2117
rect 1596 1927 1630 1945
rect 1596 1859 1630 1873
rect 1596 1791 1630 1801
rect 1596 1723 1630 1729
rect 1596 1655 1630 1657
rect 1596 1619 1630 1621
rect 1596 1547 1630 1553
rect 1596 1475 1630 1485
rect 1596 1403 1630 1417
rect 1596 1331 1630 1349
rect 1596 1259 1630 1281
rect 1596 1187 1630 1213
rect 1596 1115 1630 1145
rect 1596 1043 1630 1077
rect 1596 975 1630 1009
rect 1596 907 1630 937
rect 1596 839 1630 865
rect 1596 771 1630 793
rect 1596 703 1630 721
rect 1596 635 1630 649
rect 1596 567 1630 577
rect 1596 499 1630 505
rect 1596 431 1630 433
rect 1596 395 1630 397
rect 1596 323 1630 329
rect 1596 251 1630 261
rect 1596 179 1630 193
rect 1596 107 1630 125
rect 1596 22 1630 57
rect 1684 1995 1718 2326
rect 1841 2273 1913 2291
rect 1841 2239 1860 2273
rect 1894 2239 1913 2273
rect 1841 2221 1913 2239
rect 1753 2169 1825 2187
rect 1753 2135 1772 2169
rect 1806 2135 1825 2169
rect 1753 2117 1825 2135
rect 1684 1927 1718 1945
rect 1684 1859 1718 1873
rect 1684 1791 1718 1801
rect 1684 1723 1718 1729
rect 1684 1655 1718 1657
rect 1684 1619 1718 1621
rect 1684 1547 1718 1553
rect 1684 1475 1718 1485
rect 1684 1403 1718 1417
rect 1684 1331 1718 1349
rect 1684 1259 1718 1281
rect 1684 1187 1718 1213
rect 1684 1115 1718 1145
rect 1684 1043 1718 1077
rect 1684 975 1718 1009
rect 1684 907 1718 937
rect 1684 839 1718 865
rect 1684 771 1718 793
rect 1684 703 1718 721
rect 1684 635 1718 649
rect 1684 567 1718 577
rect 1684 499 1718 505
rect 1684 431 1718 433
rect 1684 395 1718 397
rect 1684 323 1718 329
rect 1684 251 1718 261
rect 1684 179 1718 193
rect 1684 107 1718 125
rect 1684 22 1718 57
rect 1772 1995 1806 2117
rect 1772 1927 1806 1945
rect 1772 1859 1806 1873
rect 1772 1791 1806 1801
rect 1772 1723 1806 1729
rect 1772 1655 1806 1657
rect 1772 1619 1806 1621
rect 1772 1547 1806 1553
rect 1772 1475 1806 1485
rect 1772 1403 1806 1417
rect 1772 1331 1806 1349
rect 1772 1259 1806 1281
rect 1772 1187 1806 1213
rect 1772 1115 1806 1145
rect 1772 1043 1806 1077
rect 1772 975 1806 1009
rect 1772 907 1806 937
rect 1772 839 1806 865
rect 1772 771 1806 793
rect 1772 703 1806 721
rect 1772 635 1806 649
rect 1772 567 1806 577
rect 1772 499 1806 505
rect 1772 431 1806 433
rect 1772 395 1806 397
rect 1772 323 1806 329
rect 1772 251 1806 261
rect 1772 179 1806 193
rect 1772 107 1806 125
rect 1772 22 1806 57
rect 1860 1995 1894 2221
rect 1929 2169 2001 2187
rect 1929 2135 1948 2169
rect 1982 2135 2001 2169
rect 1929 2117 2001 2135
rect 1860 1927 1894 1945
rect 1860 1859 1894 1873
rect 1860 1791 1894 1801
rect 1860 1723 1894 1729
rect 1860 1655 1894 1657
rect 1860 1619 1894 1621
rect 1860 1547 1894 1553
rect 1860 1475 1894 1485
rect 1860 1403 1894 1417
rect 1860 1331 1894 1349
rect 1860 1259 1894 1281
rect 1860 1187 1894 1213
rect 1860 1115 1894 1145
rect 1860 1043 1894 1077
rect 1860 975 1894 1009
rect 1860 907 1894 937
rect 1860 839 1894 865
rect 1860 771 1894 793
rect 1860 703 1894 721
rect 1860 635 1894 649
rect 1860 567 1894 577
rect 1860 499 1894 505
rect 1860 431 1894 433
rect 1860 395 1894 397
rect 1860 323 1894 329
rect 1860 251 1894 261
rect 1860 179 1894 193
rect 1860 107 1894 125
rect 1860 22 1894 57
rect 1948 1995 1982 2117
rect 1948 1927 1982 1945
rect 1948 1859 1982 1873
rect 1948 1791 1982 1801
rect 1948 1723 1982 1729
rect 1948 1655 1982 1657
rect 1948 1619 1982 1621
rect 1948 1547 1982 1553
rect 1948 1475 1982 1485
rect 1948 1403 1982 1417
rect 1948 1331 1982 1349
rect 1948 1259 1982 1281
rect 1948 1187 1982 1213
rect 1948 1115 1982 1145
rect 1948 1043 1982 1077
rect 1948 975 1982 1009
rect 1948 907 1982 937
rect 1948 839 1982 865
rect 1948 771 1982 793
rect 1948 703 1982 721
rect 1948 635 1982 649
rect 1948 567 1982 577
rect 1948 499 1982 505
rect 1948 431 1982 433
rect 1948 395 1982 397
rect 1948 323 1982 329
rect 1948 251 1982 261
rect 1948 179 1982 193
rect 1948 107 1982 125
rect 1948 22 1982 57
rect 2036 1995 2070 2326
rect 2193 2273 2265 2291
rect 2193 2239 2212 2273
rect 2246 2239 2265 2273
rect 2193 2221 2265 2239
rect 2369 2273 2441 2291
rect 2369 2239 2388 2273
rect 2422 2239 2441 2273
rect 2369 2221 2441 2239
rect 2545 2273 2617 2291
rect 2545 2239 2564 2273
rect 2598 2239 2617 2273
rect 2545 2221 2617 2239
rect 2105 2169 2177 2187
rect 2105 2135 2124 2169
rect 2158 2135 2177 2169
rect 2105 2117 2177 2135
rect 2036 1927 2070 1945
rect 2036 1859 2070 1873
rect 2036 1791 2070 1801
rect 2036 1723 2070 1729
rect 2036 1655 2070 1657
rect 2036 1619 2070 1621
rect 2036 1547 2070 1553
rect 2036 1475 2070 1485
rect 2036 1403 2070 1417
rect 2036 1331 2070 1349
rect 2036 1259 2070 1281
rect 2036 1187 2070 1213
rect 2036 1115 2070 1145
rect 2036 1043 2070 1077
rect 2036 975 2070 1009
rect 2036 907 2070 937
rect 2036 839 2070 865
rect 2036 771 2070 793
rect 2036 703 2070 721
rect 2036 635 2070 649
rect 2036 567 2070 577
rect 2036 499 2070 505
rect 2036 431 2070 433
rect 2036 395 2070 397
rect 2036 323 2070 329
rect 2036 251 2070 261
rect 2036 179 2070 193
rect 2036 107 2070 125
rect 2036 22 2070 57
rect 2124 1995 2158 2117
rect 2124 1927 2158 1945
rect 2124 1859 2158 1873
rect 2124 1791 2158 1801
rect 2124 1723 2158 1729
rect 2124 1655 2158 1657
rect 2124 1619 2158 1621
rect 2124 1547 2158 1553
rect 2124 1475 2158 1485
rect 2124 1403 2158 1417
rect 2124 1331 2158 1349
rect 2124 1259 2158 1281
rect 2124 1187 2158 1213
rect 2124 1115 2158 1145
rect 2124 1043 2158 1077
rect 2124 975 2158 1009
rect 2124 907 2158 937
rect 2124 839 2158 865
rect 2124 771 2158 793
rect 2124 703 2158 721
rect 2124 635 2158 649
rect 2124 567 2158 577
rect 2124 499 2158 505
rect 2124 431 2158 433
rect 2124 395 2158 397
rect 2124 323 2158 329
rect 2124 251 2158 261
rect 2124 179 2158 193
rect 2124 107 2158 125
rect 2124 22 2158 57
rect 2212 1995 2246 2221
rect 2281 2169 2353 2187
rect 2281 2135 2300 2169
rect 2334 2135 2353 2169
rect 2281 2117 2353 2135
rect 2212 1927 2246 1945
rect 2212 1859 2246 1873
rect 2212 1791 2246 1801
rect 2212 1723 2246 1729
rect 2212 1655 2246 1657
rect 2212 1619 2246 1621
rect 2212 1547 2246 1553
rect 2212 1475 2246 1485
rect 2212 1403 2246 1417
rect 2212 1331 2246 1349
rect 2212 1259 2246 1281
rect 2212 1187 2246 1213
rect 2212 1115 2246 1145
rect 2212 1043 2246 1077
rect 2212 975 2246 1009
rect 2212 907 2246 937
rect 2212 839 2246 865
rect 2212 771 2246 793
rect 2212 703 2246 721
rect 2212 635 2246 649
rect 2212 567 2246 577
rect 2212 499 2246 505
rect 2212 431 2246 433
rect 2212 395 2246 397
rect 2212 323 2246 329
rect 2212 251 2246 261
rect 2212 179 2246 193
rect 2212 107 2246 125
rect 2212 22 2246 57
rect 2300 1995 2334 2117
rect 2300 1927 2334 1945
rect 2300 1859 2334 1873
rect 2300 1791 2334 1801
rect 2300 1723 2334 1729
rect 2300 1655 2334 1657
rect 2300 1619 2334 1621
rect 2300 1547 2334 1553
rect 2300 1475 2334 1485
rect 2300 1403 2334 1417
rect 2300 1331 2334 1349
rect 2300 1259 2334 1281
rect 2300 1187 2334 1213
rect 2300 1115 2334 1145
rect 2300 1043 2334 1077
rect 2300 975 2334 1009
rect 2300 907 2334 937
rect 2300 839 2334 865
rect 2300 771 2334 793
rect 2300 703 2334 721
rect 2300 635 2334 649
rect 2300 567 2334 577
rect 2300 499 2334 505
rect 2300 431 2334 433
rect 2300 395 2334 397
rect 2300 323 2334 329
rect 2300 251 2334 261
rect 2300 179 2334 193
rect 2300 107 2334 125
rect 2300 22 2334 57
rect 2388 1995 2422 2221
rect 2457 2169 2529 2187
rect 2457 2135 2476 2169
rect 2510 2135 2529 2169
rect 2457 2117 2529 2135
rect 2388 1927 2422 1945
rect 2388 1859 2422 1873
rect 2388 1791 2422 1801
rect 2388 1723 2422 1729
rect 2388 1655 2422 1657
rect 2388 1619 2422 1621
rect 2388 1547 2422 1553
rect 2388 1475 2422 1485
rect 2388 1403 2422 1417
rect 2388 1331 2422 1349
rect 2388 1259 2422 1281
rect 2388 1187 2422 1213
rect 2388 1115 2422 1145
rect 2388 1043 2422 1077
rect 2388 975 2422 1009
rect 2388 907 2422 937
rect 2388 839 2422 865
rect 2388 771 2422 793
rect 2388 703 2422 721
rect 2388 635 2422 649
rect 2388 567 2422 577
rect 2388 499 2422 505
rect 2388 431 2422 433
rect 2388 395 2422 397
rect 2388 323 2422 329
rect 2388 251 2422 261
rect 2388 179 2422 193
rect 2388 107 2422 125
rect 2388 22 2422 57
rect 2476 1995 2510 2117
rect 2476 1927 2510 1945
rect 2476 1859 2510 1873
rect 2476 1791 2510 1801
rect 2476 1723 2510 1729
rect 2476 1655 2510 1657
rect 2476 1619 2510 1621
rect 2476 1547 2510 1553
rect 2476 1475 2510 1485
rect 2476 1403 2510 1417
rect 2476 1331 2510 1349
rect 2476 1259 2510 1281
rect 2476 1187 2510 1213
rect 2476 1115 2510 1145
rect 2476 1043 2510 1077
rect 2476 975 2510 1009
rect 2476 907 2510 937
rect 2476 839 2510 865
rect 2476 771 2510 793
rect 2476 703 2510 721
rect 2476 635 2510 649
rect 2476 567 2510 577
rect 2476 499 2510 505
rect 2476 431 2510 433
rect 2476 395 2510 397
rect 2476 323 2510 329
rect 2476 251 2510 261
rect 2476 179 2510 193
rect 2476 107 2510 125
rect 2476 22 2510 57
rect 2564 1995 2598 2221
rect 2633 2169 2705 2187
rect 2633 2135 2652 2169
rect 2686 2135 2705 2169
rect 2633 2117 2705 2135
rect 2564 1927 2598 1945
rect 2564 1859 2598 1873
rect 2564 1791 2598 1801
rect 2564 1723 2598 1729
rect 2564 1655 2598 1657
rect 2564 1619 2598 1621
rect 2564 1547 2598 1553
rect 2564 1475 2598 1485
rect 2564 1403 2598 1417
rect 2564 1331 2598 1349
rect 2564 1259 2598 1281
rect 2564 1187 2598 1213
rect 2564 1115 2598 1145
rect 2564 1043 2598 1077
rect 2564 975 2598 1009
rect 2564 907 2598 937
rect 2564 839 2598 865
rect 2564 771 2598 793
rect 2564 703 2598 721
rect 2564 635 2598 649
rect 2564 567 2598 577
rect 2564 499 2598 505
rect 2564 431 2598 433
rect 2564 395 2598 397
rect 2564 323 2598 329
rect 2564 251 2598 261
rect 2564 179 2598 193
rect 2564 107 2598 125
rect 2564 22 2598 57
rect 2652 1995 2686 2117
rect 2652 1927 2686 1945
rect 2652 1859 2686 1873
rect 2652 1791 2686 1801
rect 2652 1723 2686 1729
rect 2652 1655 2686 1657
rect 2652 1619 2686 1621
rect 2652 1547 2686 1553
rect 2652 1475 2686 1485
rect 2652 1403 2686 1417
rect 2652 1331 2686 1349
rect 2652 1259 2686 1281
rect 2652 1187 2686 1213
rect 2652 1115 2686 1145
rect 2652 1043 2686 1077
rect 2652 975 2686 1009
rect 2652 907 2686 937
rect 2652 839 2686 865
rect 2652 771 2686 793
rect 2652 703 2686 721
rect 2652 635 2686 649
rect 2652 567 2686 577
rect 2652 499 2686 505
rect 2652 431 2686 433
rect 2652 395 2686 397
rect 2652 323 2686 329
rect 2652 251 2686 261
rect 2652 179 2686 193
rect 2652 107 2686 125
rect 2652 22 2686 57
rect 2974 1981 3195 2573
rect 2974 43 2999 1981
rect 3169 43 3195 1981
rect 48 -29 528 -14
rect 48 -63 100 -29
rect 134 -63 276 -29
rect 310 -63 452 -29
rect 486 -63 528 -29
rect 48 -211 528 -63
rect 586 -29 704 -14
rect 586 -92 628 -29
rect 662 -92 704 -29
rect 586 -135 704 -92
rect 938 -29 1056 -14
rect 938 -92 980 -29
rect 1014 -92 1056 -29
rect 938 -135 1056 -92
rect 1290 -29 1408 -14
rect 1290 -92 1332 -29
rect 1366 -92 1408 -29
rect 1290 -135 1408 -92
rect 1642 -29 1760 -14
rect 1642 -92 1684 -29
rect 1718 -92 1760 -29
rect 1642 -135 1760 -92
rect 1994 -29 2112 -14
rect 1994 -92 2036 -29
rect 2070 -92 2112 -29
rect 1994 -135 2112 -92
rect 2346 -29 2464 -14
rect 2346 -92 2388 -29
rect 2422 -92 2464 -29
rect 2346 -135 2464 -92
rect 2522 -29 2640 -14
rect 2522 -92 2564 -29
rect 2598 -92 2640 -29
rect 2522 -135 2640 -92
rect 48 -245 96 -211
rect 130 -245 168 -211
rect 202 -245 240 -211
rect 274 -245 312 -211
rect 346 -245 384 -211
rect 418 -245 456 -211
rect 490 -245 528 -211
rect 48 -302 528 -245
rect 762 -193 880 -178
rect 762 -256 804 -193
rect 838 -256 880 -193
rect 762 -299 880 -256
rect 1114 -193 1232 -178
rect 1114 -256 1156 -193
rect 1190 -256 1232 -193
rect 1114 -299 1232 -256
rect 1466 -193 1584 -178
rect 1466 -256 1508 -193
rect 1542 -256 1584 -193
rect 1466 -299 1584 -256
rect 1818 -193 1936 -178
rect 1818 -256 1860 -193
rect 1894 -256 1936 -193
rect 1818 -299 1936 -256
rect 2170 -193 2288 -178
rect 2170 -256 2212 -193
rect 2246 -256 2288 -193
rect 2170 -299 2288 -256
rect 2974 -392 3195 43
rect -399 -425 3195 -392
rect -399 -595 -85 -425
rect 2669 -557 3195 -425
rect 2669 -595 3194 -557
rect -399 -627 3194 -595
<< viali >>
rect 628 2344 662 2378
rect 980 2344 1014 2378
rect 1332 2344 1366 2378
rect 1684 2344 1718 2378
rect 2036 2344 2070 2378
rect 100 2239 134 2273
rect 276 2239 310 2273
rect 452 2239 486 2273
rect 12 2135 46 2169
rect 12 1961 46 1979
rect 12 1945 46 1961
rect 12 1893 46 1907
rect 12 1873 46 1893
rect 12 1825 46 1835
rect 12 1801 46 1825
rect 12 1757 46 1763
rect 12 1729 46 1757
rect 12 1689 46 1691
rect 12 1657 46 1689
rect 12 1587 46 1619
rect 12 1585 46 1587
rect 12 1519 46 1547
rect 12 1513 46 1519
rect 12 1451 46 1475
rect 12 1441 46 1451
rect 12 1383 46 1403
rect 12 1369 46 1383
rect 12 1315 46 1331
rect 12 1297 46 1315
rect 12 1247 46 1259
rect 12 1225 46 1247
rect 12 1179 46 1187
rect 12 1153 46 1179
rect 12 1111 46 1115
rect 12 1081 46 1111
rect 12 1009 46 1043
rect 12 941 46 971
rect 12 937 46 941
rect 12 873 46 899
rect 12 865 46 873
rect 12 805 46 827
rect 12 793 46 805
rect 12 737 46 755
rect 12 721 46 737
rect 12 669 46 683
rect 12 649 46 669
rect 12 601 46 611
rect 12 577 46 601
rect 12 533 46 539
rect 12 505 46 533
rect 12 465 46 467
rect 12 433 46 465
rect 12 363 46 395
rect 12 361 46 363
rect 12 295 46 323
rect 12 289 46 295
rect 12 227 46 251
rect 12 217 46 227
rect 12 159 46 179
rect 12 145 46 159
rect 12 91 46 107
rect 12 73 46 91
rect 188 2135 222 2169
rect 100 1961 134 1979
rect 100 1945 134 1961
rect 100 1893 134 1907
rect 100 1873 134 1893
rect 100 1825 134 1835
rect 100 1801 134 1825
rect 100 1757 134 1763
rect 100 1729 134 1757
rect 100 1689 134 1691
rect 100 1657 134 1689
rect 100 1587 134 1619
rect 100 1585 134 1587
rect 100 1519 134 1547
rect 100 1513 134 1519
rect 100 1451 134 1475
rect 100 1441 134 1451
rect 100 1383 134 1403
rect 100 1369 134 1383
rect 100 1315 134 1331
rect 100 1297 134 1315
rect 100 1247 134 1259
rect 100 1225 134 1247
rect 100 1179 134 1187
rect 100 1153 134 1179
rect 100 1111 134 1115
rect 100 1081 134 1111
rect 100 1009 134 1043
rect 100 941 134 971
rect 100 937 134 941
rect 100 873 134 899
rect 100 865 134 873
rect 100 805 134 827
rect 100 793 134 805
rect 100 737 134 755
rect 100 721 134 737
rect 100 669 134 683
rect 100 649 134 669
rect 100 601 134 611
rect 100 577 134 601
rect 100 533 134 539
rect 100 505 134 533
rect 100 465 134 467
rect 100 433 134 465
rect 100 363 134 395
rect 100 361 134 363
rect 100 295 134 323
rect 100 289 134 295
rect 100 227 134 251
rect 100 217 134 227
rect 100 159 134 179
rect 100 145 134 159
rect 100 91 134 107
rect 100 73 134 91
rect 188 1961 222 1979
rect 188 1945 222 1961
rect 188 1893 222 1907
rect 188 1873 222 1893
rect 188 1825 222 1835
rect 188 1801 222 1825
rect 188 1757 222 1763
rect 188 1729 222 1757
rect 188 1689 222 1691
rect 188 1657 222 1689
rect 188 1587 222 1619
rect 188 1585 222 1587
rect 188 1519 222 1547
rect 188 1513 222 1519
rect 188 1451 222 1475
rect 188 1441 222 1451
rect 188 1383 222 1403
rect 188 1369 222 1383
rect 188 1315 222 1331
rect 188 1297 222 1315
rect 188 1247 222 1259
rect 188 1225 222 1247
rect 188 1179 222 1187
rect 188 1153 222 1179
rect 188 1111 222 1115
rect 188 1081 222 1111
rect 188 1009 222 1043
rect 188 941 222 971
rect 188 937 222 941
rect 188 873 222 899
rect 188 865 222 873
rect 188 805 222 827
rect 188 793 222 805
rect 188 737 222 755
rect 188 721 222 737
rect 188 669 222 683
rect 188 649 222 669
rect 188 601 222 611
rect 188 577 222 601
rect 188 533 222 539
rect 188 505 222 533
rect 188 465 222 467
rect 188 433 222 465
rect 188 363 222 395
rect 188 361 222 363
rect 188 295 222 323
rect 188 289 222 295
rect 188 227 222 251
rect 188 217 222 227
rect 188 159 222 179
rect 188 145 222 159
rect 188 91 222 107
rect 188 73 222 91
rect 364 2135 398 2169
rect 276 1961 310 1979
rect 276 1945 310 1961
rect 276 1893 310 1907
rect 276 1873 310 1893
rect 276 1825 310 1835
rect 276 1801 310 1825
rect 276 1757 310 1763
rect 276 1729 310 1757
rect 276 1689 310 1691
rect 276 1657 310 1689
rect 276 1587 310 1619
rect 276 1585 310 1587
rect 276 1519 310 1547
rect 276 1513 310 1519
rect 276 1451 310 1475
rect 276 1441 310 1451
rect 276 1383 310 1403
rect 276 1369 310 1383
rect 276 1315 310 1331
rect 276 1297 310 1315
rect 276 1247 310 1259
rect 276 1225 310 1247
rect 276 1179 310 1187
rect 276 1153 310 1179
rect 276 1111 310 1115
rect 276 1081 310 1111
rect 276 1009 310 1043
rect 276 941 310 971
rect 276 937 310 941
rect 276 873 310 899
rect 276 865 310 873
rect 276 805 310 827
rect 276 793 310 805
rect 276 737 310 755
rect 276 721 310 737
rect 276 669 310 683
rect 276 649 310 669
rect 276 601 310 611
rect 276 577 310 601
rect 276 533 310 539
rect 276 505 310 533
rect 276 465 310 467
rect 276 433 310 465
rect 276 363 310 395
rect 276 361 310 363
rect 276 295 310 323
rect 276 289 310 295
rect 276 227 310 251
rect 276 217 310 227
rect 276 159 310 179
rect 276 145 310 159
rect 276 91 310 107
rect 276 73 310 91
rect 364 1961 398 1979
rect 364 1945 398 1961
rect 364 1893 398 1907
rect 364 1873 398 1893
rect 364 1825 398 1835
rect 364 1801 398 1825
rect 364 1757 398 1763
rect 364 1729 398 1757
rect 364 1689 398 1691
rect 364 1657 398 1689
rect 364 1587 398 1619
rect 364 1585 398 1587
rect 364 1519 398 1547
rect 364 1513 398 1519
rect 364 1451 398 1475
rect 364 1441 398 1451
rect 364 1383 398 1403
rect 364 1369 398 1383
rect 364 1315 398 1331
rect 364 1297 398 1315
rect 364 1247 398 1259
rect 364 1225 398 1247
rect 364 1179 398 1187
rect 364 1153 398 1179
rect 364 1111 398 1115
rect 364 1081 398 1111
rect 364 1009 398 1043
rect 364 941 398 971
rect 364 937 398 941
rect 364 873 398 899
rect 364 865 398 873
rect 364 805 398 827
rect 364 793 398 805
rect 364 737 398 755
rect 364 721 398 737
rect 364 669 398 683
rect 364 649 398 669
rect 364 601 398 611
rect 364 577 398 601
rect 364 533 398 539
rect 364 505 398 533
rect 364 465 398 467
rect 364 433 398 465
rect 364 363 398 395
rect 364 361 398 363
rect 364 295 398 323
rect 364 289 398 295
rect 364 227 398 251
rect 364 217 398 227
rect 364 159 398 179
rect 364 145 398 159
rect 364 91 398 107
rect 364 73 398 91
rect 540 2135 574 2169
rect 452 1961 486 1979
rect 452 1945 486 1961
rect 452 1893 486 1907
rect 452 1873 486 1893
rect 452 1825 486 1835
rect 452 1801 486 1825
rect 452 1757 486 1763
rect 452 1729 486 1757
rect 452 1689 486 1691
rect 452 1657 486 1689
rect 452 1587 486 1619
rect 452 1585 486 1587
rect 452 1519 486 1547
rect 452 1513 486 1519
rect 452 1451 486 1475
rect 452 1441 486 1451
rect 452 1383 486 1403
rect 452 1369 486 1383
rect 452 1315 486 1331
rect 452 1297 486 1315
rect 452 1247 486 1259
rect 452 1225 486 1247
rect 452 1179 486 1187
rect 452 1153 486 1179
rect 452 1111 486 1115
rect 452 1081 486 1111
rect 452 1009 486 1043
rect 452 941 486 971
rect 452 937 486 941
rect 452 873 486 899
rect 452 865 486 873
rect 452 805 486 827
rect 452 793 486 805
rect 452 737 486 755
rect 452 721 486 737
rect 452 669 486 683
rect 452 649 486 669
rect 452 601 486 611
rect 452 577 486 601
rect 452 533 486 539
rect 452 505 486 533
rect 452 465 486 467
rect 452 433 486 465
rect 452 363 486 395
rect 452 361 486 363
rect 452 295 486 323
rect 452 289 486 295
rect 452 227 486 251
rect 452 217 486 227
rect 452 159 486 179
rect 452 145 486 159
rect 452 91 486 107
rect 452 73 486 91
rect 540 1961 574 1979
rect 540 1945 574 1961
rect 540 1893 574 1907
rect 540 1873 574 1893
rect 540 1825 574 1835
rect 540 1801 574 1825
rect 540 1757 574 1763
rect 540 1729 574 1757
rect 540 1689 574 1691
rect 540 1657 574 1689
rect 540 1587 574 1619
rect 540 1585 574 1587
rect 540 1519 574 1547
rect 540 1513 574 1519
rect 540 1451 574 1475
rect 540 1441 574 1451
rect 540 1383 574 1403
rect 540 1369 574 1383
rect 540 1315 574 1331
rect 540 1297 574 1315
rect 540 1247 574 1259
rect 540 1225 574 1247
rect 540 1179 574 1187
rect 540 1153 574 1179
rect 540 1111 574 1115
rect 540 1081 574 1111
rect 540 1009 574 1043
rect 540 941 574 971
rect 540 937 574 941
rect 540 873 574 899
rect 540 865 574 873
rect 540 805 574 827
rect 540 793 574 805
rect 540 737 574 755
rect 540 721 574 737
rect 540 669 574 683
rect 540 649 574 669
rect 540 601 574 611
rect 540 577 574 601
rect 540 533 574 539
rect 540 505 574 533
rect 540 465 574 467
rect 540 433 574 465
rect 540 363 574 395
rect 540 361 574 363
rect 540 295 574 323
rect 540 289 574 295
rect 540 227 574 251
rect 540 217 574 227
rect 540 159 574 179
rect 540 145 574 159
rect 540 91 574 107
rect 540 73 574 91
rect 804 2239 838 2273
rect 716 2135 750 2169
rect 628 1961 662 1979
rect 628 1945 662 1961
rect 628 1893 662 1907
rect 628 1873 662 1893
rect 628 1825 662 1835
rect 628 1801 662 1825
rect 628 1757 662 1763
rect 628 1729 662 1757
rect 628 1689 662 1691
rect 628 1657 662 1689
rect 628 1587 662 1619
rect 628 1585 662 1587
rect 628 1519 662 1547
rect 628 1513 662 1519
rect 628 1451 662 1475
rect 628 1441 662 1451
rect 628 1383 662 1403
rect 628 1369 662 1383
rect 628 1315 662 1331
rect 628 1297 662 1315
rect 628 1247 662 1259
rect 628 1225 662 1247
rect 628 1179 662 1187
rect 628 1153 662 1179
rect 628 1111 662 1115
rect 628 1081 662 1111
rect 628 1009 662 1043
rect 628 941 662 971
rect 628 937 662 941
rect 628 873 662 899
rect 628 865 662 873
rect 628 805 662 827
rect 628 793 662 805
rect 628 737 662 755
rect 628 721 662 737
rect 628 669 662 683
rect 628 649 662 669
rect 628 601 662 611
rect 628 577 662 601
rect 628 533 662 539
rect 628 505 662 533
rect 628 465 662 467
rect 628 433 662 465
rect 628 363 662 395
rect 628 361 662 363
rect 628 295 662 323
rect 628 289 662 295
rect 628 227 662 251
rect 628 217 662 227
rect 628 159 662 179
rect 628 145 662 159
rect 628 91 662 107
rect 628 73 662 91
rect 716 1961 750 1979
rect 716 1945 750 1961
rect 716 1893 750 1907
rect 716 1873 750 1893
rect 716 1825 750 1835
rect 716 1801 750 1825
rect 716 1757 750 1763
rect 716 1729 750 1757
rect 716 1689 750 1691
rect 716 1657 750 1689
rect 716 1587 750 1619
rect 716 1585 750 1587
rect 716 1519 750 1547
rect 716 1513 750 1519
rect 716 1451 750 1475
rect 716 1441 750 1451
rect 716 1383 750 1403
rect 716 1369 750 1383
rect 716 1315 750 1331
rect 716 1297 750 1315
rect 716 1247 750 1259
rect 716 1225 750 1247
rect 716 1179 750 1187
rect 716 1153 750 1179
rect 716 1111 750 1115
rect 716 1081 750 1111
rect 716 1009 750 1043
rect 716 941 750 971
rect 716 937 750 941
rect 716 873 750 899
rect 716 865 750 873
rect 716 805 750 827
rect 716 793 750 805
rect 716 737 750 755
rect 716 721 750 737
rect 716 669 750 683
rect 716 649 750 669
rect 716 601 750 611
rect 716 577 750 601
rect 716 533 750 539
rect 716 505 750 533
rect 716 465 750 467
rect 716 433 750 465
rect 716 363 750 395
rect 716 361 750 363
rect 716 295 750 323
rect 716 289 750 295
rect 716 227 750 251
rect 716 217 750 227
rect 716 159 750 179
rect 716 145 750 159
rect 716 91 750 107
rect 716 73 750 91
rect 892 2135 926 2169
rect 804 1961 838 1979
rect 804 1945 838 1961
rect 804 1893 838 1907
rect 804 1873 838 1893
rect 804 1825 838 1835
rect 804 1801 838 1825
rect 804 1757 838 1763
rect 804 1729 838 1757
rect 804 1689 838 1691
rect 804 1657 838 1689
rect 804 1587 838 1619
rect 804 1585 838 1587
rect 804 1519 838 1547
rect 804 1513 838 1519
rect 804 1451 838 1475
rect 804 1441 838 1451
rect 804 1383 838 1403
rect 804 1369 838 1383
rect 804 1315 838 1331
rect 804 1297 838 1315
rect 804 1247 838 1259
rect 804 1225 838 1247
rect 804 1179 838 1187
rect 804 1153 838 1179
rect 804 1111 838 1115
rect 804 1081 838 1111
rect 804 1009 838 1043
rect 804 941 838 971
rect 804 937 838 941
rect 804 873 838 899
rect 804 865 838 873
rect 804 805 838 827
rect 804 793 838 805
rect 804 737 838 755
rect 804 721 838 737
rect 804 669 838 683
rect 804 649 838 669
rect 804 601 838 611
rect 804 577 838 601
rect 804 533 838 539
rect 804 505 838 533
rect 804 465 838 467
rect 804 433 838 465
rect 804 363 838 395
rect 804 361 838 363
rect 804 295 838 323
rect 804 289 838 295
rect 804 227 838 251
rect 804 217 838 227
rect 804 159 838 179
rect 804 145 838 159
rect 804 91 838 107
rect 804 73 838 91
rect 892 1961 926 1979
rect 892 1945 926 1961
rect 892 1893 926 1907
rect 892 1873 926 1893
rect 892 1825 926 1835
rect 892 1801 926 1825
rect 892 1757 926 1763
rect 892 1729 926 1757
rect 892 1689 926 1691
rect 892 1657 926 1689
rect 892 1587 926 1619
rect 892 1585 926 1587
rect 892 1519 926 1547
rect 892 1513 926 1519
rect 892 1451 926 1475
rect 892 1441 926 1451
rect 892 1383 926 1403
rect 892 1369 926 1383
rect 892 1315 926 1331
rect 892 1297 926 1315
rect 892 1247 926 1259
rect 892 1225 926 1247
rect 892 1179 926 1187
rect 892 1153 926 1179
rect 892 1111 926 1115
rect 892 1081 926 1111
rect 892 1009 926 1043
rect 892 941 926 971
rect 892 937 926 941
rect 892 873 926 899
rect 892 865 926 873
rect 892 805 926 827
rect 892 793 926 805
rect 892 737 926 755
rect 892 721 926 737
rect 892 669 926 683
rect 892 649 926 669
rect 892 601 926 611
rect 892 577 926 601
rect 892 533 926 539
rect 892 505 926 533
rect 892 465 926 467
rect 892 433 926 465
rect 892 363 926 395
rect 892 361 926 363
rect 892 295 926 323
rect 892 289 926 295
rect 892 227 926 251
rect 892 217 926 227
rect 892 159 926 179
rect 892 145 926 159
rect 892 91 926 107
rect 892 73 926 91
rect 1156 2239 1190 2273
rect 1068 2135 1102 2169
rect 980 1961 1014 1979
rect 980 1945 1014 1961
rect 980 1893 1014 1907
rect 980 1873 1014 1893
rect 980 1825 1014 1835
rect 980 1801 1014 1825
rect 980 1757 1014 1763
rect 980 1729 1014 1757
rect 980 1689 1014 1691
rect 980 1657 1014 1689
rect 980 1587 1014 1619
rect 980 1585 1014 1587
rect 980 1519 1014 1547
rect 980 1513 1014 1519
rect 980 1451 1014 1475
rect 980 1441 1014 1451
rect 980 1383 1014 1403
rect 980 1369 1014 1383
rect 980 1315 1014 1331
rect 980 1297 1014 1315
rect 980 1247 1014 1259
rect 980 1225 1014 1247
rect 980 1179 1014 1187
rect 980 1153 1014 1179
rect 980 1111 1014 1115
rect 980 1081 1014 1111
rect 980 1009 1014 1043
rect 980 941 1014 971
rect 980 937 1014 941
rect 980 873 1014 899
rect 980 865 1014 873
rect 980 805 1014 827
rect 980 793 1014 805
rect 980 737 1014 755
rect 980 721 1014 737
rect 980 669 1014 683
rect 980 649 1014 669
rect 980 601 1014 611
rect 980 577 1014 601
rect 980 533 1014 539
rect 980 505 1014 533
rect 980 465 1014 467
rect 980 433 1014 465
rect 980 363 1014 395
rect 980 361 1014 363
rect 980 295 1014 323
rect 980 289 1014 295
rect 980 227 1014 251
rect 980 217 1014 227
rect 980 159 1014 179
rect 980 145 1014 159
rect 980 91 1014 107
rect 980 73 1014 91
rect 1068 1961 1102 1979
rect 1068 1945 1102 1961
rect 1068 1893 1102 1907
rect 1068 1873 1102 1893
rect 1068 1825 1102 1835
rect 1068 1801 1102 1825
rect 1068 1757 1102 1763
rect 1068 1729 1102 1757
rect 1068 1689 1102 1691
rect 1068 1657 1102 1689
rect 1068 1587 1102 1619
rect 1068 1585 1102 1587
rect 1068 1519 1102 1547
rect 1068 1513 1102 1519
rect 1068 1451 1102 1475
rect 1068 1441 1102 1451
rect 1068 1383 1102 1403
rect 1068 1369 1102 1383
rect 1068 1315 1102 1331
rect 1068 1297 1102 1315
rect 1068 1247 1102 1259
rect 1068 1225 1102 1247
rect 1068 1179 1102 1187
rect 1068 1153 1102 1179
rect 1068 1111 1102 1115
rect 1068 1081 1102 1111
rect 1068 1009 1102 1043
rect 1068 941 1102 971
rect 1068 937 1102 941
rect 1068 873 1102 899
rect 1068 865 1102 873
rect 1068 805 1102 827
rect 1068 793 1102 805
rect 1068 737 1102 755
rect 1068 721 1102 737
rect 1068 669 1102 683
rect 1068 649 1102 669
rect 1068 601 1102 611
rect 1068 577 1102 601
rect 1068 533 1102 539
rect 1068 505 1102 533
rect 1068 465 1102 467
rect 1068 433 1102 465
rect 1068 363 1102 395
rect 1068 361 1102 363
rect 1068 295 1102 323
rect 1068 289 1102 295
rect 1068 227 1102 251
rect 1068 217 1102 227
rect 1068 159 1102 179
rect 1068 145 1102 159
rect 1068 91 1102 107
rect 1068 73 1102 91
rect 1244 2135 1278 2169
rect 1156 1961 1190 1979
rect 1156 1945 1190 1961
rect 1156 1893 1190 1907
rect 1156 1873 1190 1893
rect 1156 1825 1190 1835
rect 1156 1801 1190 1825
rect 1156 1757 1190 1763
rect 1156 1729 1190 1757
rect 1156 1689 1190 1691
rect 1156 1657 1190 1689
rect 1156 1587 1190 1619
rect 1156 1585 1190 1587
rect 1156 1519 1190 1547
rect 1156 1513 1190 1519
rect 1156 1451 1190 1475
rect 1156 1441 1190 1451
rect 1156 1383 1190 1403
rect 1156 1369 1190 1383
rect 1156 1315 1190 1331
rect 1156 1297 1190 1315
rect 1156 1247 1190 1259
rect 1156 1225 1190 1247
rect 1156 1179 1190 1187
rect 1156 1153 1190 1179
rect 1156 1111 1190 1115
rect 1156 1081 1190 1111
rect 1156 1009 1190 1043
rect 1156 941 1190 971
rect 1156 937 1190 941
rect 1156 873 1190 899
rect 1156 865 1190 873
rect 1156 805 1190 827
rect 1156 793 1190 805
rect 1156 737 1190 755
rect 1156 721 1190 737
rect 1156 669 1190 683
rect 1156 649 1190 669
rect 1156 601 1190 611
rect 1156 577 1190 601
rect 1156 533 1190 539
rect 1156 505 1190 533
rect 1156 465 1190 467
rect 1156 433 1190 465
rect 1156 363 1190 395
rect 1156 361 1190 363
rect 1156 295 1190 323
rect 1156 289 1190 295
rect 1156 227 1190 251
rect 1156 217 1190 227
rect 1156 159 1190 179
rect 1156 145 1190 159
rect 1156 91 1190 107
rect 1156 73 1190 91
rect 1244 1961 1278 1979
rect 1244 1945 1278 1961
rect 1244 1893 1278 1907
rect 1244 1873 1278 1893
rect 1244 1825 1278 1835
rect 1244 1801 1278 1825
rect 1244 1757 1278 1763
rect 1244 1729 1278 1757
rect 1244 1689 1278 1691
rect 1244 1657 1278 1689
rect 1244 1587 1278 1619
rect 1244 1585 1278 1587
rect 1244 1519 1278 1547
rect 1244 1513 1278 1519
rect 1244 1451 1278 1475
rect 1244 1441 1278 1451
rect 1244 1383 1278 1403
rect 1244 1369 1278 1383
rect 1244 1315 1278 1331
rect 1244 1297 1278 1315
rect 1244 1247 1278 1259
rect 1244 1225 1278 1247
rect 1244 1179 1278 1187
rect 1244 1153 1278 1179
rect 1244 1111 1278 1115
rect 1244 1081 1278 1111
rect 1244 1009 1278 1043
rect 1244 941 1278 971
rect 1244 937 1278 941
rect 1244 873 1278 899
rect 1244 865 1278 873
rect 1244 805 1278 827
rect 1244 793 1278 805
rect 1244 737 1278 755
rect 1244 721 1278 737
rect 1244 669 1278 683
rect 1244 649 1278 669
rect 1244 601 1278 611
rect 1244 577 1278 601
rect 1244 533 1278 539
rect 1244 505 1278 533
rect 1244 465 1278 467
rect 1244 433 1278 465
rect 1244 363 1278 395
rect 1244 361 1278 363
rect 1244 295 1278 323
rect 1244 289 1278 295
rect 1244 227 1278 251
rect 1244 217 1278 227
rect 1244 159 1278 179
rect 1244 145 1278 159
rect 1244 91 1278 107
rect 1244 73 1278 91
rect 1508 2239 1542 2273
rect 1420 2135 1454 2169
rect 1332 1961 1366 1979
rect 1332 1945 1366 1961
rect 1332 1893 1366 1907
rect 1332 1873 1366 1893
rect 1332 1825 1366 1835
rect 1332 1801 1366 1825
rect 1332 1757 1366 1763
rect 1332 1729 1366 1757
rect 1332 1689 1366 1691
rect 1332 1657 1366 1689
rect 1332 1587 1366 1619
rect 1332 1585 1366 1587
rect 1332 1519 1366 1547
rect 1332 1513 1366 1519
rect 1332 1451 1366 1475
rect 1332 1441 1366 1451
rect 1332 1383 1366 1403
rect 1332 1369 1366 1383
rect 1332 1315 1366 1331
rect 1332 1297 1366 1315
rect 1332 1247 1366 1259
rect 1332 1225 1366 1247
rect 1332 1179 1366 1187
rect 1332 1153 1366 1179
rect 1332 1111 1366 1115
rect 1332 1081 1366 1111
rect 1332 1009 1366 1043
rect 1332 941 1366 971
rect 1332 937 1366 941
rect 1332 873 1366 899
rect 1332 865 1366 873
rect 1332 805 1366 827
rect 1332 793 1366 805
rect 1332 737 1366 755
rect 1332 721 1366 737
rect 1332 669 1366 683
rect 1332 649 1366 669
rect 1332 601 1366 611
rect 1332 577 1366 601
rect 1332 533 1366 539
rect 1332 505 1366 533
rect 1332 465 1366 467
rect 1332 433 1366 465
rect 1332 363 1366 395
rect 1332 361 1366 363
rect 1332 295 1366 323
rect 1332 289 1366 295
rect 1332 227 1366 251
rect 1332 217 1366 227
rect 1332 159 1366 179
rect 1332 145 1366 159
rect 1332 91 1366 107
rect 1332 73 1366 91
rect 1420 1961 1454 1979
rect 1420 1945 1454 1961
rect 1420 1893 1454 1907
rect 1420 1873 1454 1893
rect 1420 1825 1454 1835
rect 1420 1801 1454 1825
rect 1420 1757 1454 1763
rect 1420 1729 1454 1757
rect 1420 1689 1454 1691
rect 1420 1657 1454 1689
rect 1420 1587 1454 1619
rect 1420 1585 1454 1587
rect 1420 1519 1454 1547
rect 1420 1513 1454 1519
rect 1420 1451 1454 1475
rect 1420 1441 1454 1451
rect 1420 1383 1454 1403
rect 1420 1369 1454 1383
rect 1420 1315 1454 1331
rect 1420 1297 1454 1315
rect 1420 1247 1454 1259
rect 1420 1225 1454 1247
rect 1420 1179 1454 1187
rect 1420 1153 1454 1179
rect 1420 1111 1454 1115
rect 1420 1081 1454 1111
rect 1420 1009 1454 1043
rect 1420 941 1454 971
rect 1420 937 1454 941
rect 1420 873 1454 899
rect 1420 865 1454 873
rect 1420 805 1454 827
rect 1420 793 1454 805
rect 1420 737 1454 755
rect 1420 721 1454 737
rect 1420 669 1454 683
rect 1420 649 1454 669
rect 1420 601 1454 611
rect 1420 577 1454 601
rect 1420 533 1454 539
rect 1420 505 1454 533
rect 1420 465 1454 467
rect 1420 433 1454 465
rect 1420 363 1454 395
rect 1420 361 1454 363
rect 1420 295 1454 323
rect 1420 289 1454 295
rect 1420 227 1454 251
rect 1420 217 1454 227
rect 1420 159 1454 179
rect 1420 145 1454 159
rect 1420 91 1454 107
rect 1420 73 1454 91
rect 1596 2135 1630 2169
rect 1508 1961 1542 1979
rect 1508 1945 1542 1961
rect 1508 1893 1542 1907
rect 1508 1873 1542 1893
rect 1508 1825 1542 1835
rect 1508 1801 1542 1825
rect 1508 1757 1542 1763
rect 1508 1729 1542 1757
rect 1508 1689 1542 1691
rect 1508 1657 1542 1689
rect 1508 1587 1542 1619
rect 1508 1585 1542 1587
rect 1508 1519 1542 1547
rect 1508 1513 1542 1519
rect 1508 1451 1542 1475
rect 1508 1441 1542 1451
rect 1508 1383 1542 1403
rect 1508 1369 1542 1383
rect 1508 1315 1542 1331
rect 1508 1297 1542 1315
rect 1508 1247 1542 1259
rect 1508 1225 1542 1247
rect 1508 1179 1542 1187
rect 1508 1153 1542 1179
rect 1508 1111 1542 1115
rect 1508 1081 1542 1111
rect 1508 1009 1542 1043
rect 1508 941 1542 971
rect 1508 937 1542 941
rect 1508 873 1542 899
rect 1508 865 1542 873
rect 1508 805 1542 827
rect 1508 793 1542 805
rect 1508 737 1542 755
rect 1508 721 1542 737
rect 1508 669 1542 683
rect 1508 649 1542 669
rect 1508 601 1542 611
rect 1508 577 1542 601
rect 1508 533 1542 539
rect 1508 505 1542 533
rect 1508 465 1542 467
rect 1508 433 1542 465
rect 1508 363 1542 395
rect 1508 361 1542 363
rect 1508 295 1542 323
rect 1508 289 1542 295
rect 1508 227 1542 251
rect 1508 217 1542 227
rect 1508 159 1542 179
rect 1508 145 1542 159
rect 1508 91 1542 107
rect 1508 73 1542 91
rect 1596 1961 1630 1979
rect 1596 1945 1630 1961
rect 1596 1893 1630 1907
rect 1596 1873 1630 1893
rect 1596 1825 1630 1835
rect 1596 1801 1630 1825
rect 1596 1757 1630 1763
rect 1596 1729 1630 1757
rect 1596 1689 1630 1691
rect 1596 1657 1630 1689
rect 1596 1587 1630 1619
rect 1596 1585 1630 1587
rect 1596 1519 1630 1547
rect 1596 1513 1630 1519
rect 1596 1451 1630 1475
rect 1596 1441 1630 1451
rect 1596 1383 1630 1403
rect 1596 1369 1630 1383
rect 1596 1315 1630 1331
rect 1596 1297 1630 1315
rect 1596 1247 1630 1259
rect 1596 1225 1630 1247
rect 1596 1179 1630 1187
rect 1596 1153 1630 1179
rect 1596 1111 1630 1115
rect 1596 1081 1630 1111
rect 1596 1009 1630 1043
rect 1596 941 1630 971
rect 1596 937 1630 941
rect 1596 873 1630 899
rect 1596 865 1630 873
rect 1596 805 1630 827
rect 1596 793 1630 805
rect 1596 737 1630 755
rect 1596 721 1630 737
rect 1596 669 1630 683
rect 1596 649 1630 669
rect 1596 601 1630 611
rect 1596 577 1630 601
rect 1596 533 1630 539
rect 1596 505 1630 533
rect 1596 465 1630 467
rect 1596 433 1630 465
rect 1596 363 1630 395
rect 1596 361 1630 363
rect 1596 295 1630 323
rect 1596 289 1630 295
rect 1596 227 1630 251
rect 1596 217 1630 227
rect 1596 159 1630 179
rect 1596 145 1630 159
rect 1596 91 1630 107
rect 1596 73 1630 91
rect 1860 2239 1894 2273
rect 1772 2135 1806 2169
rect 1684 1961 1718 1979
rect 1684 1945 1718 1961
rect 1684 1893 1718 1907
rect 1684 1873 1718 1893
rect 1684 1825 1718 1835
rect 1684 1801 1718 1825
rect 1684 1757 1718 1763
rect 1684 1729 1718 1757
rect 1684 1689 1718 1691
rect 1684 1657 1718 1689
rect 1684 1587 1718 1619
rect 1684 1585 1718 1587
rect 1684 1519 1718 1547
rect 1684 1513 1718 1519
rect 1684 1451 1718 1475
rect 1684 1441 1718 1451
rect 1684 1383 1718 1403
rect 1684 1369 1718 1383
rect 1684 1315 1718 1331
rect 1684 1297 1718 1315
rect 1684 1247 1718 1259
rect 1684 1225 1718 1247
rect 1684 1179 1718 1187
rect 1684 1153 1718 1179
rect 1684 1111 1718 1115
rect 1684 1081 1718 1111
rect 1684 1009 1718 1043
rect 1684 941 1718 971
rect 1684 937 1718 941
rect 1684 873 1718 899
rect 1684 865 1718 873
rect 1684 805 1718 827
rect 1684 793 1718 805
rect 1684 737 1718 755
rect 1684 721 1718 737
rect 1684 669 1718 683
rect 1684 649 1718 669
rect 1684 601 1718 611
rect 1684 577 1718 601
rect 1684 533 1718 539
rect 1684 505 1718 533
rect 1684 465 1718 467
rect 1684 433 1718 465
rect 1684 363 1718 395
rect 1684 361 1718 363
rect 1684 295 1718 323
rect 1684 289 1718 295
rect 1684 227 1718 251
rect 1684 217 1718 227
rect 1684 159 1718 179
rect 1684 145 1718 159
rect 1684 91 1718 107
rect 1684 73 1718 91
rect 1772 1961 1806 1979
rect 1772 1945 1806 1961
rect 1772 1893 1806 1907
rect 1772 1873 1806 1893
rect 1772 1825 1806 1835
rect 1772 1801 1806 1825
rect 1772 1757 1806 1763
rect 1772 1729 1806 1757
rect 1772 1689 1806 1691
rect 1772 1657 1806 1689
rect 1772 1587 1806 1619
rect 1772 1585 1806 1587
rect 1772 1519 1806 1547
rect 1772 1513 1806 1519
rect 1772 1451 1806 1475
rect 1772 1441 1806 1451
rect 1772 1383 1806 1403
rect 1772 1369 1806 1383
rect 1772 1315 1806 1331
rect 1772 1297 1806 1315
rect 1772 1247 1806 1259
rect 1772 1225 1806 1247
rect 1772 1179 1806 1187
rect 1772 1153 1806 1179
rect 1772 1111 1806 1115
rect 1772 1081 1806 1111
rect 1772 1009 1806 1043
rect 1772 941 1806 971
rect 1772 937 1806 941
rect 1772 873 1806 899
rect 1772 865 1806 873
rect 1772 805 1806 827
rect 1772 793 1806 805
rect 1772 737 1806 755
rect 1772 721 1806 737
rect 1772 669 1806 683
rect 1772 649 1806 669
rect 1772 601 1806 611
rect 1772 577 1806 601
rect 1772 533 1806 539
rect 1772 505 1806 533
rect 1772 465 1806 467
rect 1772 433 1806 465
rect 1772 363 1806 395
rect 1772 361 1806 363
rect 1772 295 1806 323
rect 1772 289 1806 295
rect 1772 227 1806 251
rect 1772 217 1806 227
rect 1772 159 1806 179
rect 1772 145 1806 159
rect 1772 91 1806 107
rect 1772 73 1806 91
rect 1948 2135 1982 2169
rect 1860 1961 1894 1979
rect 1860 1945 1894 1961
rect 1860 1893 1894 1907
rect 1860 1873 1894 1893
rect 1860 1825 1894 1835
rect 1860 1801 1894 1825
rect 1860 1757 1894 1763
rect 1860 1729 1894 1757
rect 1860 1689 1894 1691
rect 1860 1657 1894 1689
rect 1860 1587 1894 1619
rect 1860 1585 1894 1587
rect 1860 1519 1894 1547
rect 1860 1513 1894 1519
rect 1860 1451 1894 1475
rect 1860 1441 1894 1451
rect 1860 1383 1894 1403
rect 1860 1369 1894 1383
rect 1860 1315 1894 1331
rect 1860 1297 1894 1315
rect 1860 1247 1894 1259
rect 1860 1225 1894 1247
rect 1860 1179 1894 1187
rect 1860 1153 1894 1179
rect 1860 1111 1894 1115
rect 1860 1081 1894 1111
rect 1860 1009 1894 1043
rect 1860 941 1894 971
rect 1860 937 1894 941
rect 1860 873 1894 899
rect 1860 865 1894 873
rect 1860 805 1894 827
rect 1860 793 1894 805
rect 1860 737 1894 755
rect 1860 721 1894 737
rect 1860 669 1894 683
rect 1860 649 1894 669
rect 1860 601 1894 611
rect 1860 577 1894 601
rect 1860 533 1894 539
rect 1860 505 1894 533
rect 1860 465 1894 467
rect 1860 433 1894 465
rect 1860 363 1894 395
rect 1860 361 1894 363
rect 1860 295 1894 323
rect 1860 289 1894 295
rect 1860 227 1894 251
rect 1860 217 1894 227
rect 1860 159 1894 179
rect 1860 145 1894 159
rect 1860 91 1894 107
rect 1860 73 1894 91
rect 1948 1961 1982 1979
rect 1948 1945 1982 1961
rect 1948 1893 1982 1907
rect 1948 1873 1982 1893
rect 1948 1825 1982 1835
rect 1948 1801 1982 1825
rect 1948 1757 1982 1763
rect 1948 1729 1982 1757
rect 1948 1689 1982 1691
rect 1948 1657 1982 1689
rect 1948 1587 1982 1619
rect 1948 1585 1982 1587
rect 1948 1519 1982 1547
rect 1948 1513 1982 1519
rect 1948 1451 1982 1475
rect 1948 1441 1982 1451
rect 1948 1383 1982 1403
rect 1948 1369 1982 1383
rect 1948 1315 1982 1331
rect 1948 1297 1982 1315
rect 1948 1247 1982 1259
rect 1948 1225 1982 1247
rect 1948 1179 1982 1187
rect 1948 1153 1982 1179
rect 1948 1111 1982 1115
rect 1948 1081 1982 1111
rect 1948 1009 1982 1043
rect 1948 941 1982 971
rect 1948 937 1982 941
rect 1948 873 1982 899
rect 1948 865 1982 873
rect 1948 805 1982 827
rect 1948 793 1982 805
rect 1948 737 1982 755
rect 1948 721 1982 737
rect 1948 669 1982 683
rect 1948 649 1982 669
rect 1948 601 1982 611
rect 1948 577 1982 601
rect 1948 533 1982 539
rect 1948 505 1982 533
rect 1948 465 1982 467
rect 1948 433 1982 465
rect 1948 363 1982 395
rect 1948 361 1982 363
rect 1948 295 1982 323
rect 1948 289 1982 295
rect 1948 227 1982 251
rect 1948 217 1982 227
rect 1948 159 1982 179
rect 1948 145 1982 159
rect 1948 91 1982 107
rect 1948 73 1982 91
rect 2212 2239 2246 2273
rect 2388 2239 2422 2273
rect 2564 2239 2598 2273
rect 2124 2135 2158 2169
rect 2036 1961 2070 1979
rect 2036 1945 2070 1961
rect 2036 1893 2070 1907
rect 2036 1873 2070 1893
rect 2036 1825 2070 1835
rect 2036 1801 2070 1825
rect 2036 1757 2070 1763
rect 2036 1729 2070 1757
rect 2036 1689 2070 1691
rect 2036 1657 2070 1689
rect 2036 1587 2070 1619
rect 2036 1585 2070 1587
rect 2036 1519 2070 1547
rect 2036 1513 2070 1519
rect 2036 1451 2070 1475
rect 2036 1441 2070 1451
rect 2036 1383 2070 1403
rect 2036 1369 2070 1383
rect 2036 1315 2070 1331
rect 2036 1297 2070 1315
rect 2036 1247 2070 1259
rect 2036 1225 2070 1247
rect 2036 1179 2070 1187
rect 2036 1153 2070 1179
rect 2036 1111 2070 1115
rect 2036 1081 2070 1111
rect 2036 1009 2070 1043
rect 2036 941 2070 971
rect 2036 937 2070 941
rect 2036 873 2070 899
rect 2036 865 2070 873
rect 2036 805 2070 827
rect 2036 793 2070 805
rect 2036 737 2070 755
rect 2036 721 2070 737
rect 2036 669 2070 683
rect 2036 649 2070 669
rect 2036 601 2070 611
rect 2036 577 2070 601
rect 2036 533 2070 539
rect 2036 505 2070 533
rect 2036 465 2070 467
rect 2036 433 2070 465
rect 2036 363 2070 395
rect 2036 361 2070 363
rect 2036 295 2070 323
rect 2036 289 2070 295
rect 2036 227 2070 251
rect 2036 217 2070 227
rect 2036 159 2070 179
rect 2036 145 2070 159
rect 2036 91 2070 107
rect 2036 73 2070 91
rect 2124 1961 2158 1979
rect 2124 1945 2158 1961
rect 2124 1893 2158 1907
rect 2124 1873 2158 1893
rect 2124 1825 2158 1835
rect 2124 1801 2158 1825
rect 2124 1757 2158 1763
rect 2124 1729 2158 1757
rect 2124 1689 2158 1691
rect 2124 1657 2158 1689
rect 2124 1587 2158 1619
rect 2124 1585 2158 1587
rect 2124 1519 2158 1547
rect 2124 1513 2158 1519
rect 2124 1451 2158 1475
rect 2124 1441 2158 1451
rect 2124 1383 2158 1403
rect 2124 1369 2158 1383
rect 2124 1315 2158 1331
rect 2124 1297 2158 1315
rect 2124 1247 2158 1259
rect 2124 1225 2158 1247
rect 2124 1179 2158 1187
rect 2124 1153 2158 1179
rect 2124 1111 2158 1115
rect 2124 1081 2158 1111
rect 2124 1009 2158 1043
rect 2124 941 2158 971
rect 2124 937 2158 941
rect 2124 873 2158 899
rect 2124 865 2158 873
rect 2124 805 2158 827
rect 2124 793 2158 805
rect 2124 737 2158 755
rect 2124 721 2158 737
rect 2124 669 2158 683
rect 2124 649 2158 669
rect 2124 601 2158 611
rect 2124 577 2158 601
rect 2124 533 2158 539
rect 2124 505 2158 533
rect 2124 465 2158 467
rect 2124 433 2158 465
rect 2124 363 2158 395
rect 2124 361 2158 363
rect 2124 295 2158 323
rect 2124 289 2158 295
rect 2124 227 2158 251
rect 2124 217 2158 227
rect 2124 159 2158 179
rect 2124 145 2158 159
rect 2124 91 2158 107
rect 2124 73 2158 91
rect 2300 2135 2334 2169
rect 2212 1961 2246 1979
rect 2212 1945 2246 1961
rect 2212 1893 2246 1907
rect 2212 1873 2246 1893
rect 2212 1825 2246 1835
rect 2212 1801 2246 1825
rect 2212 1757 2246 1763
rect 2212 1729 2246 1757
rect 2212 1689 2246 1691
rect 2212 1657 2246 1689
rect 2212 1587 2246 1619
rect 2212 1585 2246 1587
rect 2212 1519 2246 1547
rect 2212 1513 2246 1519
rect 2212 1451 2246 1475
rect 2212 1441 2246 1451
rect 2212 1383 2246 1403
rect 2212 1369 2246 1383
rect 2212 1315 2246 1331
rect 2212 1297 2246 1315
rect 2212 1247 2246 1259
rect 2212 1225 2246 1247
rect 2212 1179 2246 1187
rect 2212 1153 2246 1179
rect 2212 1111 2246 1115
rect 2212 1081 2246 1111
rect 2212 1009 2246 1043
rect 2212 941 2246 971
rect 2212 937 2246 941
rect 2212 873 2246 899
rect 2212 865 2246 873
rect 2212 805 2246 827
rect 2212 793 2246 805
rect 2212 737 2246 755
rect 2212 721 2246 737
rect 2212 669 2246 683
rect 2212 649 2246 669
rect 2212 601 2246 611
rect 2212 577 2246 601
rect 2212 533 2246 539
rect 2212 505 2246 533
rect 2212 465 2246 467
rect 2212 433 2246 465
rect 2212 363 2246 395
rect 2212 361 2246 363
rect 2212 295 2246 323
rect 2212 289 2246 295
rect 2212 227 2246 251
rect 2212 217 2246 227
rect 2212 159 2246 179
rect 2212 145 2246 159
rect 2212 91 2246 107
rect 2212 73 2246 91
rect 2300 1961 2334 1979
rect 2300 1945 2334 1961
rect 2300 1893 2334 1907
rect 2300 1873 2334 1893
rect 2300 1825 2334 1835
rect 2300 1801 2334 1825
rect 2300 1757 2334 1763
rect 2300 1729 2334 1757
rect 2300 1689 2334 1691
rect 2300 1657 2334 1689
rect 2300 1587 2334 1619
rect 2300 1585 2334 1587
rect 2300 1519 2334 1547
rect 2300 1513 2334 1519
rect 2300 1451 2334 1475
rect 2300 1441 2334 1451
rect 2300 1383 2334 1403
rect 2300 1369 2334 1383
rect 2300 1315 2334 1331
rect 2300 1297 2334 1315
rect 2300 1247 2334 1259
rect 2300 1225 2334 1247
rect 2300 1179 2334 1187
rect 2300 1153 2334 1179
rect 2300 1111 2334 1115
rect 2300 1081 2334 1111
rect 2300 1009 2334 1043
rect 2300 941 2334 971
rect 2300 937 2334 941
rect 2300 873 2334 899
rect 2300 865 2334 873
rect 2300 805 2334 827
rect 2300 793 2334 805
rect 2300 737 2334 755
rect 2300 721 2334 737
rect 2300 669 2334 683
rect 2300 649 2334 669
rect 2300 601 2334 611
rect 2300 577 2334 601
rect 2300 533 2334 539
rect 2300 505 2334 533
rect 2300 465 2334 467
rect 2300 433 2334 465
rect 2300 363 2334 395
rect 2300 361 2334 363
rect 2300 295 2334 323
rect 2300 289 2334 295
rect 2300 227 2334 251
rect 2300 217 2334 227
rect 2300 159 2334 179
rect 2300 145 2334 159
rect 2300 91 2334 107
rect 2300 73 2334 91
rect 2476 2135 2510 2169
rect 2388 1961 2422 1979
rect 2388 1945 2422 1961
rect 2388 1893 2422 1907
rect 2388 1873 2422 1893
rect 2388 1825 2422 1835
rect 2388 1801 2422 1825
rect 2388 1757 2422 1763
rect 2388 1729 2422 1757
rect 2388 1689 2422 1691
rect 2388 1657 2422 1689
rect 2388 1587 2422 1619
rect 2388 1585 2422 1587
rect 2388 1519 2422 1547
rect 2388 1513 2422 1519
rect 2388 1451 2422 1475
rect 2388 1441 2422 1451
rect 2388 1383 2422 1403
rect 2388 1369 2422 1383
rect 2388 1315 2422 1331
rect 2388 1297 2422 1315
rect 2388 1247 2422 1259
rect 2388 1225 2422 1247
rect 2388 1179 2422 1187
rect 2388 1153 2422 1179
rect 2388 1111 2422 1115
rect 2388 1081 2422 1111
rect 2388 1009 2422 1043
rect 2388 941 2422 971
rect 2388 937 2422 941
rect 2388 873 2422 899
rect 2388 865 2422 873
rect 2388 805 2422 827
rect 2388 793 2422 805
rect 2388 737 2422 755
rect 2388 721 2422 737
rect 2388 669 2422 683
rect 2388 649 2422 669
rect 2388 601 2422 611
rect 2388 577 2422 601
rect 2388 533 2422 539
rect 2388 505 2422 533
rect 2388 465 2422 467
rect 2388 433 2422 465
rect 2388 363 2422 395
rect 2388 361 2422 363
rect 2388 295 2422 323
rect 2388 289 2422 295
rect 2388 227 2422 251
rect 2388 217 2422 227
rect 2388 159 2422 179
rect 2388 145 2422 159
rect 2388 91 2422 107
rect 2388 73 2422 91
rect 2476 1961 2510 1979
rect 2476 1945 2510 1961
rect 2476 1893 2510 1907
rect 2476 1873 2510 1893
rect 2476 1825 2510 1835
rect 2476 1801 2510 1825
rect 2476 1757 2510 1763
rect 2476 1729 2510 1757
rect 2476 1689 2510 1691
rect 2476 1657 2510 1689
rect 2476 1587 2510 1619
rect 2476 1585 2510 1587
rect 2476 1519 2510 1547
rect 2476 1513 2510 1519
rect 2476 1451 2510 1475
rect 2476 1441 2510 1451
rect 2476 1383 2510 1403
rect 2476 1369 2510 1383
rect 2476 1315 2510 1331
rect 2476 1297 2510 1315
rect 2476 1247 2510 1259
rect 2476 1225 2510 1247
rect 2476 1179 2510 1187
rect 2476 1153 2510 1179
rect 2476 1111 2510 1115
rect 2476 1081 2510 1111
rect 2476 1009 2510 1043
rect 2476 941 2510 971
rect 2476 937 2510 941
rect 2476 873 2510 899
rect 2476 865 2510 873
rect 2476 805 2510 827
rect 2476 793 2510 805
rect 2476 737 2510 755
rect 2476 721 2510 737
rect 2476 669 2510 683
rect 2476 649 2510 669
rect 2476 601 2510 611
rect 2476 577 2510 601
rect 2476 533 2510 539
rect 2476 505 2510 533
rect 2476 465 2510 467
rect 2476 433 2510 465
rect 2476 363 2510 395
rect 2476 361 2510 363
rect 2476 295 2510 323
rect 2476 289 2510 295
rect 2476 227 2510 251
rect 2476 217 2510 227
rect 2476 159 2510 179
rect 2476 145 2510 159
rect 2476 91 2510 107
rect 2476 73 2510 91
rect 2652 2135 2686 2169
rect 2564 1961 2598 1979
rect 2564 1945 2598 1961
rect 2564 1893 2598 1907
rect 2564 1873 2598 1893
rect 2564 1825 2598 1835
rect 2564 1801 2598 1825
rect 2564 1757 2598 1763
rect 2564 1729 2598 1757
rect 2564 1689 2598 1691
rect 2564 1657 2598 1689
rect 2564 1587 2598 1619
rect 2564 1585 2598 1587
rect 2564 1519 2598 1547
rect 2564 1513 2598 1519
rect 2564 1451 2598 1475
rect 2564 1441 2598 1451
rect 2564 1383 2598 1403
rect 2564 1369 2598 1383
rect 2564 1315 2598 1331
rect 2564 1297 2598 1315
rect 2564 1247 2598 1259
rect 2564 1225 2598 1247
rect 2564 1179 2598 1187
rect 2564 1153 2598 1179
rect 2564 1111 2598 1115
rect 2564 1081 2598 1111
rect 2564 1009 2598 1043
rect 2564 941 2598 971
rect 2564 937 2598 941
rect 2564 873 2598 899
rect 2564 865 2598 873
rect 2564 805 2598 827
rect 2564 793 2598 805
rect 2564 737 2598 755
rect 2564 721 2598 737
rect 2564 669 2598 683
rect 2564 649 2598 669
rect 2564 601 2598 611
rect 2564 577 2598 601
rect 2564 533 2598 539
rect 2564 505 2598 533
rect 2564 465 2598 467
rect 2564 433 2598 465
rect 2564 363 2598 395
rect 2564 361 2598 363
rect 2564 295 2598 323
rect 2564 289 2598 295
rect 2564 227 2598 251
rect 2564 217 2598 227
rect 2564 159 2598 179
rect 2564 145 2598 159
rect 2564 91 2598 107
rect 2564 73 2598 91
rect 2652 1961 2686 1979
rect 2652 1945 2686 1961
rect 2652 1893 2686 1907
rect 2652 1873 2686 1893
rect 2652 1825 2686 1835
rect 2652 1801 2686 1825
rect 2652 1757 2686 1763
rect 2652 1729 2686 1757
rect 2652 1689 2686 1691
rect 2652 1657 2686 1689
rect 2652 1587 2686 1619
rect 2652 1585 2686 1587
rect 2652 1519 2686 1547
rect 2652 1513 2686 1519
rect 2652 1451 2686 1475
rect 2652 1441 2686 1451
rect 2652 1383 2686 1403
rect 2652 1369 2686 1383
rect 2652 1315 2686 1331
rect 2652 1297 2686 1315
rect 2652 1247 2686 1259
rect 2652 1225 2686 1247
rect 2652 1179 2686 1187
rect 2652 1153 2686 1179
rect 2652 1111 2686 1115
rect 2652 1081 2686 1111
rect 2652 1009 2686 1043
rect 2652 941 2686 971
rect 2652 937 2686 941
rect 2652 873 2686 899
rect 2652 865 2686 873
rect 2652 805 2686 827
rect 2652 793 2686 805
rect 2652 737 2686 755
rect 2652 721 2686 737
rect 2652 669 2686 683
rect 2652 649 2686 669
rect 2652 601 2686 611
rect 2652 577 2686 601
rect 2652 533 2686 539
rect 2652 505 2686 533
rect 2652 465 2686 467
rect 2652 433 2686 465
rect 2652 363 2686 395
rect 2652 361 2686 363
rect 2652 295 2686 323
rect 2652 289 2686 295
rect 2652 227 2686 251
rect 2652 217 2686 227
rect 2652 159 2686 179
rect 2652 145 2686 159
rect 2652 91 2686 107
rect 2652 73 2686 91
rect 628 -63 662 -58
rect 628 -92 662 -63
rect 980 -63 1014 -58
rect 980 -92 1014 -63
rect 1332 -63 1366 -58
rect 1332 -92 1366 -63
rect 1684 -63 1718 -58
rect 1684 -92 1718 -63
rect 2036 -63 2070 -58
rect 2036 -92 2070 -63
rect 2388 -63 2422 -58
rect 2388 -92 2422 -63
rect 2564 -63 2598 -58
rect 2564 -92 2598 -63
rect 96 -245 130 -211
rect 168 -245 202 -211
rect 240 -245 274 -211
rect 312 -245 346 -211
rect 384 -245 418 -211
rect 456 -245 490 -211
rect 804 -227 838 -222
rect 804 -256 838 -227
rect 1156 -227 1190 -222
rect 1156 -256 1190 -227
rect 1508 -227 1542 -222
rect 1508 -256 1542 -227
rect 1860 -227 1894 -222
rect 1860 -256 1894 -227
rect 2212 -227 2246 -222
rect 2212 -256 2246 -227
<< metal1 >>
rect 609 2378 2089 2396
rect 609 2344 628 2378
rect 662 2344 980 2378
rect 1014 2344 1332 2378
rect 1366 2344 1684 2378
rect 1718 2344 2036 2378
rect 2070 2344 2089 2378
rect 609 2326 2089 2344
rect 81 2273 2617 2291
rect 81 2239 100 2273
rect 134 2239 276 2273
rect 310 2239 452 2273
rect 486 2239 804 2273
rect 838 2239 1156 2273
rect 1190 2239 1508 2273
rect 1542 2239 1860 2273
rect 1894 2239 2212 2273
rect 2246 2239 2388 2273
rect 2422 2239 2564 2273
rect 2598 2239 2617 2273
rect 81 2221 2617 2239
rect -7 2169 2705 2187
rect -7 2135 12 2169
rect 46 2135 188 2169
rect 222 2135 364 2169
rect 398 2135 540 2169
rect 574 2135 716 2169
rect 750 2135 892 2169
rect 926 2135 1068 2169
rect 1102 2135 1244 2169
rect 1278 2135 1420 2169
rect 1454 2135 1596 2169
rect 1630 2135 1772 2169
rect 1806 2135 1948 2169
rect 1982 2135 2124 2169
rect 2158 2135 2300 2169
rect 2334 2135 2476 2169
rect 2510 2135 2652 2169
rect 2686 2135 2705 2169
rect -7 2117 2705 2135
rect 6 1979 52 2026
rect 6 1945 12 1979
rect 46 1945 52 1979
rect 6 1907 52 1945
rect 6 1873 12 1907
rect 46 1873 52 1907
rect 6 1835 52 1873
rect 6 1801 12 1835
rect 46 1801 52 1835
rect 6 1763 52 1801
rect 6 1729 12 1763
rect 46 1729 52 1763
rect 6 1691 52 1729
rect 6 1657 12 1691
rect 46 1657 52 1691
rect 6 1619 52 1657
rect 6 1585 12 1619
rect 46 1585 52 1619
rect 6 1547 52 1585
rect 6 1513 12 1547
rect 46 1513 52 1547
rect 6 1475 52 1513
rect 6 1441 12 1475
rect 46 1441 52 1475
rect 6 1403 52 1441
rect 6 1369 12 1403
rect 46 1369 52 1403
rect 6 1331 52 1369
rect 6 1297 12 1331
rect 46 1297 52 1331
rect 6 1259 52 1297
rect 6 1225 12 1259
rect 46 1225 52 1259
rect 6 1187 52 1225
rect 6 1153 12 1187
rect 46 1153 52 1187
rect 6 1115 52 1153
rect 6 1081 12 1115
rect 46 1081 52 1115
rect 6 1043 52 1081
rect 6 1009 12 1043
rect 46 1009 52 1043
rect 6 971 52 1009
rect 6 937 12 971
rect 46 937 52 971
rect 6 899 52 937
rect 6 865 12 899
rect 46 865 52 899
rect 6 827 52 865
rect 6 793 12 827
rect 46 793 52 827
rect 6 755 52 793
rect 6 721 12 755
rect 46 721 52 755
rect 6 683 52 721
rect 6 649 12 683
rect 46 649 52 683
rect 6 611 52 649
rect 6 577 12 611
rect 46 577 52 611
rect 6 539 52 577
rect 6 505 12 539
rect 46 505 52 539
rect 6 467 52 505
rect 6 433 12 467
rect 46 433 52 467
rect 6 395 52 433
rect 6 361 12 395
rect 46 361 52 395
rect 6 323 52 361
rect 6 289 12 323
rect 46 289 52 323
rect 6 251 52 289
rect 6 217 12 251
rect 46 217 52 251
rect 6 179 52 217
rect 6 145 12 179
rect 46 145 52 179
rect 6 107 52 145
rect 6 73 12 107
rect 46 73 52 107
rect 6 26 52 73
rect 94 1979 140 2026
rect 94 1945 100 1979
rect 134 1945 140 1979
rect 94 1907 140 1945
rect 94 1873 100 1907
rect 134 1873 140 1907
rect 94 1835 140 1873
rect 94 1801 100 1835
rect 134 1801 140 1835
rect 94 1763 140 1801
rect 94 1729 100 1763
rect 134 1729 140 1763
rect 94 1691 140 1729
rect 94 1657 100 1691
rect 134 1657 140 1691
rect 94 1619 140 1657
rect 94 1585 100 1619
rect 134 1585 140 1619
rect 94 1547 140 1585
rect 94 1513 100 1547
rect 134 1513 140 1547
rect 94 1475 140 1513
rect 94 1441 100 1475
rect 134 1441 140 1475
rect 94 1403 140 1441
rect 94 1369 100 1403
rect 134 1369 140 1403
rect 94 1331 140 1369
rect 94 1297 100 1331
rect 134 1297 140 1331
rect 94 1259 140 1297
rect 94 1225 100 1259
rect 134 1225 140 1259
rect 94 1187 140 1225
rect 94 1153 100 1187
rect 134 1153 140 1187
rect 94 1115 140 1153
rect 94 1081 100 1115
rect 134 1081 140 1115
rect 94 1043 140 1081
rect 94 1009 100 1043
rect 134 1009 140 1043
rect 94 971 140 1009
rect 94 937 100 971
rect 134 937 140 971
rect 94 899 140 937
rect 94 865 100 899
rect 134 865 140 899
rect 94 827 140 865
rect 94 793 100 827
rect 134 793 140 827
rect 94 755 140 793
rect 94 721 100 755
rect 134 721 140 755
rect 94 683 140 721
rect 94 649 100 683
rect 134 649 140 683
rect 94 611 140 649
rect 94 577 100 611
rect 134 577 140 611
rect 94 539 140 577
rect 94 505 100 539
rect 134 505 140 539
rect 94 467 140 505
rect 94 433 100 467
rect 134 433 140 467
rect 94 395 140 433
rect 94 361 100 395
rect 134 361 140 395
rect 94 323 140 361
rect 94 289 100 323
rect 134 289 140 323
rect 94 251 140 289
rect 94 217 100 251
rect 134 217 140 251
rect 94 179 140 217
rect 94 145 100 179
rect 134 145 140 179
rect 94 107 140 145
rect 94 73 100 107
rect 134 73 140 107
rect 94 26 140 73
rect 182 1979 228 2026
rect 182 1945 188 1979
rect 222 1945 228 1979
rect 182 1907 228 1945
rect 182 1873 188 1907
rect 222 1873 228 1907
rect 182 1835 228 1873
rect 182 1801 188 1835
rect 222 1801 228 1835
rect 182 1763 228 1801
rect 182 1729 188 1763
rect 222 1729 228 1763
rect 182 1691 228 1729
rect 182 1657 188 1691
rect 222 1657 228 1691
rect 182 1619 228 1657
rect 182 1585 188 1619
rect 222 1585 228 1619
rect 182 1547 228 1585
rect 182 1513 188 1547
rect 222 1513 228 1547
rect 182 1475 228 1513
rect 182 1441 188 1475
rect 222 1441 228 1475
rect 182 1403 228 1441
rect 182 1369 188 1403
rect 222 1369 228 1403
rect 182 1331 228 1369
rect 182 1297 188 1331
rect 222 1297 228 1331
rect 182 1259 228 1297
rect 182 1225 188 1259
rect 222 1225 228 1259
rect 182 1187 228 1225
rect 182 1153 188 1187
rect 222 1153 228 1187
rect 182 1115 228 1153
rect 182 1081 188 1115
rect 222 1081 228 1115
rect 182 1043 228 1081
rect 182 1009 188 1043
rect 222 1009 228 1043
rect 182 971 228 1009
rect 182 937 188 971
rect 222 937 228 971
rect 182 899 228 937
rect 182 865 188 899
rect 222 865 228 899
rect 182 827 228 865
rect 182 793 188 827
rect 222 793 228 827
rect 182 755 228 793
rect 182 721 188 755
rect 222 721 228 755
rect 182 683 228 721
rect 182 649 188 683
rect 222 649 228 683
rect 182 611 228 649
rect 182 577 188 611
rect 222 577 228 611
rect 182 539 228 577
rect 182 505 188 539
rect 222 505 228 539
rect 182 467 228 505
rect 182 433 188 467
rect 222 433 228 467
rect 182 395 228 433
rect 182 361 188 395
rect 222 361 228 395
rect 182 323 228 361
rect 182 289 188 323
rect 222 289 228 323
rect 182 251 228 289
rect 182 217 188 251
rect 222 217 228 251
rect 182 179 228 217
rect 182 145 188 179
rect 222 145 228 179
rect 182 107 228 145
rect 182 73 188 107
rect 222 73 228 107
rect 182 26 228 73
rect 270 1979 316 2026
rect 270 1945 276 1979
rect 310 1945 316 1979
rect 270 1907 316 1945
rect 270 1873 276 1907
rect 310 1873 316 1907
rect 270 1835 316 1873
rect 270 1801 276 1835
rect 310 1801 316 1835
rect 270 1763 316 1801
rect 270 1729 276 1763
rect 310 1729 316 1763
rect 270 1691 316 1729
rect 270 1657 276 1691
rect 310 1657 316 1691
rect 270 1619 316 1657
rect 270 1585 276 1619
rect 310 1585 316 1619
rect 270 1547 316 1585
rect 270 1513 276 1547
rect 310 1513 316 1547
rect 270 1475 316 1513
rect 270 1441 276 1475
rect 310 1441 316 1475
rect 270 1403 316 1441
rect 270 1369 276 1403
rect 310 1369 316 1403
rect 270 1331 316 1369
rect 270 1297 276 1331
rect 310 1297 316 1331
rect 270 1259 316 1297
rect 270 1225 276 1259
rect 310 1225 316 1259
rect 270 1187 316 1225
rect 270 1153 276 1187
rect 310 1153 316 1187
rect 270 1115 316 1153
rect 270 1081 276 1115
rect 310 1081 316 1115
rect 270 1043 316 1081
rect 270 1009 276 1043
rect 310 1009 316 1043
rect 270 971 316 1009
rect 270 937 276 971
rect 310 937 316 971
rect 270 899 316 937
rect 270 865 276 899
rect 310 865 316 899
rect 270 827 316 865
rect 270 793 276 827
rect 310 793 316 827
rect 270 755 316 793
rect 270 721 276 755
rect 310 721 316 755
rect 270 683 316 721
rect 270 649 276 683
rect 310 649 316 683
rect 270 611 316 649
rect 270 577 276 611
rect 310 577 316 611
rect 270 539 316 577
rect 270 505 276 539
rect 310 505 316 539
rect 270 467 316 505
rect 270 433 276 467
rect 310 433 316 467
rect 270 395 316 433
rect 270 361 276 395
rect 310 361 316 395
rect 270 323 316 361
rect 270 289 276 323
rect 310 289 316 323
rect 270 251 316 289
rect 270 217 276 251
rect 310 217 316 251
rect 270 179 316 217
rect 270 145 276 179
rect 310 145 316 179
rect 270 107 316 145
rect 270 73 276 107
rect 310 73 316 107
rect 270 26 316 73
rect 358 1979 404 2026
rect 358 1945 364 1979
rect 398 1945 404 1979
rect 358 1907 404 1945
rect 358 1873 364 1907
rect 398 1873 404 1907
rect 358 1835 404 1873
rect 358 1801 364 1835
rect 398 1801 404 1835
rect 358 1763 404 1801
rect 358 1729 364 1763
rect 398 1729 404 1763
rect 358 1691 404 1729
rect 358 1657 364 1691
rect 398 1657 404 1691
rect 358 1619 404 1657
rect 358 1585 364 1619
rect 398 1585 404 1619
rect 358 1547 404 1585
rect 358 1513 364 1547
rect 398 1513 404 1547
rect 358 1475 404 1513
rect 358 1441 364 1475
rect 398 1441 404 1475
rect 358 1403 404 1441
rect 358 1369 364 1403
rect 398 1369 404 1403
rect 358 1331 404 1369
rect 358 1297 364 1331
rect 398 1297 404 1331
rect 358 1259 404 1297
rect 358 1225 364 1259
rect 398 1225 404 1259
rect 358 1187 404 1225
rect 358 1153 364 1187
rect 398 1153 404 1187
rect 358 1115 404 1153
rect 358 1081 364 1115
rect 398 1081 404 1115
rect 358 1043 404 1081
rect 358 1009 364 1043
rect 398 1009 404 1043
rect 358 971 404 1009
rect 358 937 364 971
rect 398 937 404 971
rect 358 899 404 937
rect 358 865 364 899
rect 398 865 404 899
rect 358 827 404 865
rect 358 793 364 827
rect 398 793 404 827
rect 358 755 404 793
rect 358 721 364 755
rect 398 721 404 755
rect 358 683 404 721
rect 358 649 364 683
rect 398 649 404 683
rect 358 611 404 649
rect 358 577 364 611
rect 398 577 404 611
rect 358 539 404 577
rect 358 505 364 539
rect 398 505 404 539
rect 358 467 404 505
rect 358 433 364 467
rect 398 433 404 467
rect 358 395 404 433
rect 358 361 364 395
rect 398 361 404 395
rect 358 323 404 361
rect 358 289 364 323
rect 398 289 404 323
rect 358 251 404 289
rect 358 217 364 251
rect 398 217 404 251
rect 358 179 404 217
rect 358 145 364 179
rect 398 145 404 179
rect 358 107 404 145
rect 358 73 364 107
rect 398 73 404 107
rect 358 26 404 73
rect 446 1979 492 2026
rect 446 1945 452 1979
rect 486 1945 492 1979
rect 446 1907 492 1945
rect 446 1873 452 1907
rect 486 1873 492 1907
rect 446 1835 492 1873
rect 446 1801 452 1835
rect 486 1801 492 1835
rect 446 1763 492 1801
rect 446 1729 452 1763
rect 486 1729 492 1763
rect 446 1691 492 1729
rect 446 1657 452 1691
rect 486 1657 492 1691
rect 446 1619 492 1657
rect 446 1585 452 1619
rect 486 1585 492 1619
rect 446 1547 492 1585
rect 446 1513 452 1547
rect 486 1513 492 1547
rect 446 1475 492 1513
rect 446 1441 452 1475
rect 486 1441 492 1475
rect 446 1403 492 1441
rect 446 1369 452 1403
rect 486 1369 492 1403
rect 446 1331 492 1369
rect 446 1297 452 1331
rect 486 1297 492 1331
rect 446 1259 492 1297
rect 446 1225 452 1259
rect 486 1225 492 1259
rect 446 1187 492 1225
rect 446 1153 452 1187
rect 486 1153 492 1187
rect 446 1115 492 1153
rect 446 1081 452 1115
rect 486 1081 492 1115
rect 446 1043 492 1081
rect 446 1009 452 1043
rect 486 1009 492 1043
rect 446 971 492 1009
rect 446 937 452 971
rect 486 937 492 971
rect 446 899 492 937
rect 446 865 452 899
rect 486 865 492 899
rect 446 827 492 865
rect 446 793 452 827
rect 486 793 492 827
rect 446 755 492 793
rect 446 721 452 755
rect 486 721 492 755
rect 446 683 492 721
rect 446 649 452 683
rect 486 649 492 683
rect 446 611 492 649
rect 446 577 452 611
rect 486 577 492 611
rect 446 539 492 577
rect 446 505 452 539
rect 486 505 492 539
rect 446 467 492 505
rect 446 433 452 467
rect 486 433 492 467
rect 446 395 492 433
rect 446 361 452 395
rect 486 361 492 395
rect 446 323 492 361
rect 446 289 452 323
rect 486 289 492 323
rect 446 251 492 289
rect 446 217 452 251
rect 486 217 492 251
rect 446 179 492 217
rect 446 145 452 179
rect 486 145 492 179
rect 446 107 492 145
rect 446 73 452 107
rect 486 73 492 107
rect 446 26 492 73
rect 534 1979 580 2026
rect 534 1945 540 1979
rect 574 1945 580 1979
rect 534 1907 580 1945
rect 534 1873 540 1907
rect 574 1873 580 1907
rect 534 1835 580 1873
rect 534 1801 540 1835
rect 574 1801 580 1835
rect 534 1763 580 1801
rect 534 1729 540 1763
rect 574 1729 580 1763
rect 534 1691 580 1729
rect 534 1657 540 1691
rect 574 1657 580 1691
rect 534 1619 580 1657
rect 534 1585 540 1619
rect 574 1585 580 1619
rect 534 1547 580 1585
rect 534 1513 540 1547
rect 574 1513 580 1547
rect 534 1475 580 1513
rect 534 1441 540 1475
rect 574 1441 580 1475
rect 534 1403 580 1441
rect 534 1369 540 1403
rect 574 1369 580 1403
rect 534 1331 580 1369
rect 534 1297 540 1331
rect 574 1297 580 1331
rect 534 1259 580 1297
rect 534 1225 540 1259
rect 574 1225 580 1259
rect 534 1187 580 1225
rect 534 1153 540 1187
rect 574 1153 580 1187
rect 534 1115 580 1153
rect 534 1081 540 1115
rect 574 1081 580 1115
rect 534 1043 580 1081
rect 534 1009 540 1043
rect 574 1009 580 1043
rect 534 971 580 1009
rect 534 937 540 971
rect 574 937 580 971
rect 534 899 580 937
rect 534 865 540 899
rect 574 865 580 899
rect 534 827 580 865
rect 534 793 540 827
rect 574 793 580 827
rect 534 755 580 793
rect 534 721 540 755
rect 574 721 580 755
rect 534 683 580 721
rect 534 649 540 683
rect 574 649 580 683
rect 534 611 580 649
rect 534 577 540 611
rect 574 577 580 611
rect 534 539 580 577
rect 534 505 540 539
rect 574 505 580 539
rect 534 467 580 505
rect 534 433 540 467
rect 574 433 580 467
rect 534 395 580 433
rect 534 361 540 395
rect 574 361 580 395
rect 534 323 580 361
rect 534 289 540 323
rect 574 289 580 323
rect 534 251 580 289
rect 534 217 540 251
rect 574 217 580 251
rect 534 179 580 217
rect 534 145 540 179
rect 574 145 580 179
rect 534 107 580 145
rect 534 73 540 107
rect 574 73 580 107
rect 534 26 580 73
rect 622 1979 668 2026
rect 622 1945 628 1979
rect 662 1945 668 1979
rect 622 1907 668 1945
rect 622 1873 628 1907
rect 662 1873 668 1907
rect 622 1835 668 1873
rect 622 1801 628 1835
rect 662 1801 668 1835
rect 622 1763 668 1801
rect 622 1729 628 1763
rect 662 1729 668 1763
rect 622 1691 668 1729
rect 622 1657 628 1691
rect 662 1657 668 1691
rect 622 1619 668 1657
rect 622 1585 628 1619
rect 662 1585 668 1619
rect 622 1547 668 1585
rect 622 1513 628 1547
rect 662 1513 668 1547
rect 622 1475 668 1513
rect 622 1441 628 1475
rect 662 1441 668 1475
rect 622 1403 668 1441
rect 622 1369 628 1403
rect 662 1369 668 1403
rect 622 1331 668 1369
rect 622 1297 628 1331
rect 662 1297 668 1331
rect 622 1259 668 1297
rect 622 1225 628 1259
rect 662 1225 668 1259
rect 622 1187 668 1225
rect 622 1153 628 1187
rect 662 1153 668 1187
rect 622 1115 668 1153
rect 622 1081 628 1115
rect 662 1081 668 1115
rect 622 1043 668 1081
rect 622 1009 628 1043
rect 662 1009 668 1043
rect 622 971 668 1009
rect 622 937 628 971
rect 662 937 668 971
rect 622 899 668 937
rect 622 865 628 899
rect 662 865 668 899
rect 622 827 668 865
rect 622 793 628 827
rect 662 793 668 827
rect 622 755 668 793
rect 622 721 628 755
rect 662 721 668 755
rect 622 683 668 721
rect 622 649 628 683
rect 662 649 668 683
rect 622 611 668 649
rect 622 577 628 611
rect 662 577 668 611
rect 622 539 668 577
rect 622 505 628 539
rect 662 505 668 539
rect 622 467 668 505
rect 622 433 628 467
rect 662 433 668 467
rect 622 395 668 433
rect 622 361 628 395
rect 662 361 668 395
rect 622 323 668 361
rect 622 289 628 323
rect 662 289 668 323
rect 622 251 668 289
rect 622 217 628 251
rect 662 217 668 251
rect 622 179 668 217
rect 622 145 628 179
rect 662 145 668 179
rect 622 107 668 145
rect 622 73 628 107
rect 662 73 668 107
rect 622 26 668 73
rect 710 1979 756 2026
rect 710 1945 716 1979
rect 750 1945 756 1979
rect 710 1907 756 1945
rect 710 1873 716 1907
rect 750 1873 756 1907
rect 710 1835 756 1873
rect 710 1801 716 1835
rect 750 1801 756 1835
rect 710 1763 756 1801
rect 710 1729 716 1763
rect 750 1729 756 1763
rect 710 1691 756 1729
rect 710 1657 716 1691
rect 750 1657 756 1691
rect 710 1619 756 1657
rect 710 1585 716 1619
rect 750 1585 756 1619
rect 710 1547 756 1585
rect 710 1513 716 1547
rect 750 1513 756 1547
rect 710 1475 756 1513
rect 710 1441 716 1475
rect 750 1441 756 1475
rect 710 1403 756 1441
rect 710 1369 716 1403
rect 750 1369 756 1403
rect 710 1331 756 1369
rect 710 1297 716 1331
rect 750 1297 756 1331
rect 710 1259 756 1297
rect 710 1225 716 1259
rect 750 1225 756 1259
rect 710 1187 756 1225
rect 710 1153 716 1187
rect 750 1153 756 1187
rect 710 1115 756 1153
rect 710 1081 716 1115
rect 750 1081 756 1115
rect 710 1043 756 1081
rect 710 1009 716 1043
rect 750 1009 756 1043
rect 710 971 756 1009
rect 710 937 716 971
rect 750 937 756 971
rect 710 899 756 937
rect 710 865 716 899
rect 750 865 756 899
rect 710 827 756 865
rect 710 793 716 827
rect 750 793 756 827
rect 710 755 756 793
rect 710 721 716 755
rect 750 721 756 755
rect 710 683 756 721
rect 710 649 716 683
rect 750 649 756 683
rect 710 611 756 649
rect 710 577 716 611
rect 750 577 756 611
rect 710 539 756 577
rect 710 505 716 539
rect 750 505 756 539
rect 710 467 756 505
rect 710 433 716 467
rect 750 433 756 467
rect 710 395 756 433
rect 710 361 716 395
rect 750 361 756 395
rect 710 323 756 361
rect 710 289 716 323
rect 750 289 756 323
rect 710 251 756 289
rect 710 217 716 251
rect 750 217 756 251
rect 710 179 756 217
rect 710 145 716 179
rect 750 145 756 179
rect 710 107 756 145
rect 710 73 716 107
rect 750 73 756 107
rect 710 26 756 73
rect 798 1979 844 2026
rect 798 1945 804 1979
rect 838 1945 844 1979
rect 798 1907 844 1945
rect 798 1873 804 1907
rect 838 1873 844 1907
rect 798 1835 844 1873
rect 798 1801 804 1835
rect 838 1801 844 1835
rect 798 1763 844 1801
rect 798 1729 804 1763
rect 838 1729 844 1763
rect 798 1691 844 1729
rect 798 1657 804 1691
rect 838 1657 844 1691
rect 798 1619 844 1657
rect 798 1585 804 1619
rect 838 1585 844 1619
rect 798 1547 844 1585
rect 798 1513 804 1547
rect 838 1513 844 1547
rect 798 1475 844 1513
rect 798 1441 804 1475
rect 838 1441 844 1475
rect 798 1403 844 1441
rect 798 1369 804 1403
rect 838 1369 844 1403
rect 798 1331 844 1369
rect 798 1297 804 1331
rect 838 1297 844 1331
rect 798 1259 844 1297
rect 798 1225 804 1259
rect 838 1225 844 1259
rect 798 1187 844 1225
rect 798 1153 804 1187
rect 838 1153 844 1187
rect 798 1115 844 1153
rect 798 1081 804 1115
rect 838 1081 844 1115
rect 798 1043 844 1081
rect 798 1009 804 1043
rect 838 1009 844 1043
rect 798 971 844 1009
rect 798 937 804 971
rect 838 937 844 971
rect 798 899 844 937
rect 798 865 804 899
rect 838 865 844 899
rect 798 827 844 865
rect 798 793 804 827
rect 838 793 844 827
rect 798 755 844 793
rect 798 721 804 755
rect 838 721 844 755
rect 798 683 844 721
rect 798 649 804 683
rect 838 649 844 683
rect 798 611 844 649
rect 798 577 804 611
rect 838 577 844 611
rect 798 539 844 577
rect 798 505 804 539
rect 838 505 844 539
rect 798 467 844 505
rect 798 433 804 467
rect 838 433 844 467
rect 798 395 844 433
rect 798 361 804 395
rect 838 361 844 395
rect 798 323 844 361
rect 798 289 804 323
rect 838 289 844 323
rect 798 251 844 289
rect 798 217 804 251
rect 838 217 844 251
rect 798 179 844 217
rect 798 145 804 179
rect 838 145 844 179
rect 798 107 844 145
rect 798 73 804 107
rect 838 73 844 107
rect 798 26 844 73
rect 886 1979 932 2026
rect 886 1945 892 1979
rect 926 1945 932 1979
rect 886 1907 932 1945
rect 886 1873 892 1907
rect 926 1873 932 1907
rect 886 1835 932 1873
rect 886 1801 892 1835
rect 926 1801 932 1835
rect 886 1763 932 1801
rect 886 1729 892 1763
rect 926 1729 932 1763
rect 886 1691 932 1729
rect 886 1657 892 1691
rect 926 1657 932 1691
rect 886 1619 932 1657
rect 886 1585 892 1619
rect 926 1585 932 1619
rect 886 1547 932 1585
rect 886 1513 892 1547
rect 926 1513 932 1547
rect 886 1475 932 1513
rect 886 1441 892 1475
rect 926 1441 932 1475
rect 886 1403 932 1441
rect 886 1369 892 1403
rect 926 1369 932 1403
rect 886 1331 932 1369
rect 886 1297 892 1331
rect 926 1297 932 1331
rect 886 1259 932 1297
rect 886 1225 892 1259
rect 926 1225 932 1259
rect 886 1187 932 1225
rect 886 1153 892 1187
rect 926 1153 932 1187
rect 886 1115 932 1153
rect 886 1081 892 1115
rect 926 1081 932 1115
rect 886 1043 932 1081
rect 886 1009 892 1043
rect 926 1009 932 1043
rect 886 971 932 1009
rect 886 937 892 971
rect 926 937 932 971
rect 886 899 932 937
rect 886 865 892 899
rect 926 865 932 899
rect 886 827 932 865
rect 886 793 892 827
rect 926 793 932 827
rect 886 755 932 793
rect 886 721 892 755
rect 926 721 932 755
rect 886 683 932 721
rect 886 649 892 683
rect 926 649 932 683
rect 886 611 932 649
rect 886 577 892 611
rect 926 577 932 611
rect 886 539 932 577
rect 886 505 892 539
rect 926 505 932 539
rect 886 467 932 505
rect 886 433 892 467
rect 926 433 932 467
rect 886 395 932 433
rect 886 361 892 395
rect 926 361 932 395
rect 886 323 932 361
rect 886 289 892 323
rect 926 289 932 323
rect 886 251 932 289
rect 886 217 892 251
rect 926 217 932 251
rect 886 179 932 217
rect 886 145 892 179
rect 926 145 932 179
rect 886 107 932 145
rect 886 73 892 107
rect 926 73 932 107
rect 886 26 932 73
rect 974 1979 1020 2026
rect 974 1945 980 1979
rect 1014 1945 1020 1979
rect 974 1907 1020 1945
rect 974 1873 980 1907
rect 1014 1873 1020 1907
rect 974 1835 1020 1873
rect 974 1801 980 1835
rect 1014 1801 1020 1835
rect 974 1763 1020 1801
rect 974 1729 980 1763
rect 1014 1729 1020 1763
rect 974 1691 1020 1729
rect 974 1657 980 1691
rect 1014 1657 1020 1691
rect 974 1619 1020 1657
rect 974 1585 980 1619
rect 1014 1585 1020 1619
rect 974 1547 1020 1585
rect 974 1513 980 1547
rect 1014 1513 1020 1547
rect 974 1475 1020 1513
rect 974 1441 980 1475
rect 1014 1441 1020 1475
rect 974 1403 1020 1441
rect 974 1369 980 1403
rect 1014 1369 1020 1403
rect 974 1331 1020 1369
rect 974 1297 980 1331
rect 1014 1297 1020 1331
rect 974 1259 1020 1297
rect 974 1225 980 1259
rect 1014 1225 1020 1259
rect 974 1187 1020 1225
rect 974 1153 980 1187
rect 1014 1153 1020 1187
rect 974 1115 1020 1153
rect 974 1081 980 1115
rect 1014 1081 1020 1115
rect 974 1043 1020 1081
rect 974 1009 980 1043
rect 1014 1009 1020 1043
rect 974 971 1020 1009
rect 974 937 980 971
rect 1014 937 1020 971
rect 974 899 1020 937
rect 974 865 980 899
rect 1014 865 1020 899
rect 974 827 1020 865
rect 974 793 980 827
rect 1014 793 1020 827
rect 974 755 1020 793
rect 974 721 980 755
rect 1014 721 1020 755
rect 974 683 1020 721
rect 974 649 980 683
rect 1014 649 1020 683
rect 974 611 1020 649
rect 974 577 980 611
rect 1014 577 1020 611
rect 974 539 1020 577
rect 974 505 980 539
rect 1014 505 1020 539
rect 974 467 1020 505
rect 974 433 980 467
rect 1014 433 1020 467
rect 974 395 1020 433
rect 974 361 980 395
rect 1014 361 1020 395
rect 974 323 1020 361
rect 974 289 980 323
rect 1014 289 1020 323
rect 974 251 1020 289
rect 974 217 980 251
rect 1014 217 1020 251
rect 974 179 1020 217
rect 974 145 980 179
rect 1014 145 1020 179
rect 974 107 1020 145
rect 974 73 980 107
rect 1014 73 1020 107
rect 974 26 1020 73
rect 1062 1979 1108 2026
rect 1062 1945 1068 1979
rect 1102 1945 1108 1979
rect 1062 1907 1108 1945
rect 1062 1873 1068 1907
rect 1102 1873 1108 1907
rect 1062 1835 1108 1873
rect 1062 1801 1068 1835
rect 1102 1801 1108 1835
rect 1062 1763 1108 1801
rect 1062 1729 1068 1763
rect 1102 1729 1108 1763
rect 1062 1691 1108 1729
rect 1062 1657 1068 1691
rect 1102 1657 1108 1691
rect 1062 1619 1108 1657
rect 1062 1585 1068 1619
rect 1102 1585 1108 1619
rect 1062 1547 1108 1585
rect 1062 1513 1068 1547
rect 1102 1513 1108 1547
rect 1062 1475 1108 1513
rect 1062 1441 1068 1475
rect 1102 1441 1108 1475
rect 1062 1403 1108 1441
rect 1062 1369 1068 1403
rect 1102 1369 1108 1403
rect 1062 1331 1108 1369
rect 1062 1297 1068 1331
rect 1102 1297 1108 1331
rect 1062 1259 1108 1297
rect 1062 1225 1068 1259
rect 1102 1225 1108 1259
rect 1062 1187 1108 1225
rect 1062 1153 1068 1187
rect 1102 1153 1108 1187
rect 1062 1115 1108 1153
rect 1062 1081 1068 1115
rect 1102 1081 1108 1115
rect 1062 1043 1108 1081
rect 1062 1009 1068 1043
rect 1102 1009 1108 1043
rect 1062 971 1108 1009
rect 1062 937 1068 971
rect 1102 937 1108 971
rect 1062 899 1108 937
rect 1062 865 1068 899
rect 1102 865 1108 899
rect 1062 827 1108 865
rect 1062 793 1068 827
rect 1102 793 1108 827
rect 1062 755 1108 793
rect 1062 721 1068 755
rect 1102 721 1108 755
rect 1062 683 1108 721
rect 1062 649 1068 683
rect 1102 649 1108 683
rect 1062 611 1108 649
rect 1062 577 1068 611
rect 1102 577 1108 611
rect 1062 539 1108 577
rect 1062 505 1068 539
rect 1102 505 1108 539
rect 1062 467 1108 505
rect 1062 433 1068 467
rect 1102 433 1108 467
rect 1062 395 1108 433
rect 1062 361 1068 395
rect 1102 361 1108 395
rect 1062 323 1108 361
rect 1062 289 1068 323
rect 1102 289 1108 323
rect 1062 251 1108 289
rect 1062 217 1068 251
rect 1102 217 1108 251
rect 1062 179 1108 217
rect 1062 145 1068 179
rect 1102 145 1108 179
rect 1062 107 1108 145
rect 1062 73 1068 107
rect 1102 73 1108 107
rect 1062 26 1108 73
rect 1150 1979 1196 2026
rect 1150 1945 1156 1979
rect 1190 1945 1196 1979
rect 1150 1907 1196 1945
rect 1150 1873 1156 1907
rect 1190 1873 1196 1907
rect 1150 1835 1196 1873
rect 1150 1801 1156 1835
rect 1190 1801 1196 1835
rect 1150 1763 1196 1801
rect 1150 1729 1156 1763
rect 1190 1729 1196 1763
rect 1150 1691 1196 1729
rect 1150 1657 1156 1691
rect 1190 1657 1196 1691
rect 1150 1619 1196 1657
rect 1150 1585 1156 1619
rect 1190 1585 1196 1619
rect 1150 1547 1196 1585
rect 1150 1513 1156 1547
rect 1190 1513 1196 1547
rect 1150 1475 1196 1513
rect 1150 1441 1156 1475
rect 1190 1441 1196 1475
rect 1150 1403 1196 1441
rect 1150 1369 1156 1403
rect 1190 1369 1196 1403
rect 1150 1331 1196 1369
rect 1150 1297 1156 1331
rect 1190 1297 1196 1331
rect 1150 1259 1196 1297
rect 1150 1225 1156 1259
rect 1190 1225 1196 1259
rect 1150 1187 1196 1225
rect 1150 1153 1156 1187
rect 1190 1153 1196 1187
rect 1150 1115 1196 1153
rect 1150 1081 1156 1115
rect 1190 1081 1196 1115
rect 1150 1043 1196 1081
rect 1150 1009 1156 1043
rect 1190 1009 1196 1043
rect 1150 971 1196 1009
rect 1150 937 1156 971
rect 1190 937 1196 971
rect 1150 899 1196 937
rect 1150 865 1156 899
rect 1190 865 1196 899
rect 1150 827 1196 865
rect 1150 793 1156 827
rect 1190 793 1196 827
rect 1150 755 1196 793
rect 1150 721 1156 755
rect 1190 721 1196 755
rect 1150 683 1196 721
rect 1150 649 1156 683
rect 1190 649 1196 683
rect 1150 611 1196 649
rect 1150 577 1156 611
rect 1190 577 1196 611
rect 1150 539 1196 577
rect 1150 505 1156 539
rect 1190 505 1196 539
rect 1150 467 1196 505
rect 1150 433 1156 467
rect 1190 433 1196 467
rect 1150 395 1196 433
rect 1150 361 1156 395
rect 1190 361 1196 395
rect 1150 323 1196 361
rect 1150 289 1156 323
rect 1190 289 1196 323
rect 1150 251 1196 289
rect 1150 217 1156 251
rect 1190 217 1196 251
rect 1150 179 1196 217
rect 1150 145 1156 179
rect 1190 145 1196 179
rect 1150 107 1196 145
rect 1150 73 1156 107
rect 1190 73 1196 107
rect 1150 26 1196 73
rect 1238 1979 1284 2026
rect 1238 1945 1244 1979
rect 1278 1945 1284 1979
rect 1238 1907 1284 1945
rect 1238 1873 1244 1907
rect 1278 1873 1284 1907
rect 1238 1835 1284 1873
rect 1238 1801 1244 1835
rect 1278 1801 1284 1835
rect 1238 1763 1284 1801
rect 1238 1729 1244 1763
rect 1278 1729 1284 1763
rect 1238 1691 1284 1729
rect 1238 1657 1244 1691
rect 1278 1657 1284 1691
rect 1238 1619 1284 1657
rect 1238 1585 1244 1619
rect 1278 1585 1284 1619
rect 1238 1547 1284 1585
rect 1238 1513 1244 1547
rect 1278 1513 1284 1547
rect 1238 1475 1284 1513
rect 1238 1441 1244 1475
rect 1278 1441 1284 1475
rect 1238 1403 1284 1441
rect 1238 1369 1244 1403
rect 1278 1369 1284 1403
rect 1238 1331 1284 1369
rect 1238 1297 1244 1331
rect 1278 1297 1284 1331
rect 1238 1259 1284 1297
rect 1238 1225 1244 1259
rect 1278 1225 1284 1259
rect 1238 1187 1284 1225
rect 1238 1153 1244 1187
rect 1278 1153 1284 1187
rect 1238 1115 1284 1153
rect 1238 1081 1244 1115
rect 1278 1081 1284 1115
rect 1238 1043 1284 1081
rect 1238 1009 1244 1043
rect 1278 1009 1284 1043
rect 1238 971 1284 1009
rect 1238 937 1244 971
rect 1278 937 1284 971
rect 1238 899 1284 937
rect 1238 865 1244 899
rect 1278 865 1284 899
rect 1238 827 1284 865
rect 1238 793 1244 827
rect 1278 793 1284 827
rect 1238 755 1284 793
rect 1238 721 1244 755
rect 1278 721 1284 755
rect 1238 683 1284 721
rect 1238 649 1244 683
rect 1278 649 1284 683
rect 1238 611 1284 649
rect 1238 577 1244 611
rect 1278 577 1284 611
rect 1238 539 1284 577
rect 1238 505 1244 539
rect 1278 505 1284 539
rect 1238 467 1284 505
rect 1238 433 1244 467
rect 1278 433 1284 467
rect 1238 395 1284 433
rect 1238 361 1244 395
rect 1278 361 1284 395
rect 1238 323 1284 361
rect 1238 289 1244 323
rect 1278 289 1284 323
rect 1238 251 1284 289
rect 1238 217 1244 251
rect 1278 217 1284 251
rect 1238 179 1284 217
rect 1238 145 1244 179
rect 1278 145 1284 179
rect 1238 107 1284 145
rect 1238 73 1244 107
rect 1278 73 1284 107
rect 1238 26 1284 73
rect 1326 1979 1372 2026
rect 1326 1945 1332 1979
rect 1366 1945 1372 1979
rect 1326 1907 1372 1945
rect 1326 1873 1332 1907
rect 1366 1873 1372 1907
rect 1326 1835 1372 1873
rect 1326 1801 1332 1835
rect 1366 1801 1372 1835
rect 1326 1763 1372 1801
rect 1326 1729 1332 1763
rect 1366 1729 1372 1763
rect 1326 1691 1372 1729
rect 1326 1657 1332 1691
rect 1366 1657 1372 1691
rect 1326 1619 1372 1657
rect 1326 1585 1332 1619
rect 1366 1585 1372 1619
rect 1326 1547 1372 1585
rect 1326 1513 1332 1547
rect 1366 1513 1372 1547
rect 1326 1475 1372 1513
rect 1326 1441 1332 1475
rect 1366 1441 1372 1475
rect 1326 1403 1372 1441
rect 1326 1369 1332 1403
rect 1366 1369 1372 1403
rect 1326 1331 1372 1369
rect 1326 1297 1332 1331
rect 1366 1297 1372 1331
rect 1326 1259 1372 1297
rect 1326 1225 1332 1259
rect 1366 1225 1372 1259
rect 1326 1187 1372 1225
rect 1326 1153 1332 1187
rect 1366 1153 1372 1187
rect 1326 1115 1372 1153
rect 1326 1081 1332 1115
rect 1366 1081 1372 1115
rect 1326 1043 1372 1081
rect 1326 1009 1332 1043
rect 1366 1009 1372 1043
rect 1326 971 1372 1009
rect 1326 937 1332 971
rect 1366 937 1372 971
rect 1326 899 1372 937
rect 1326 865 1332 899
rect 1366 865 1372 899
rect 1326 827 1372 865
rect 1326 793 1332 827
rect 1366 793 1372 827
rect 1326 755 1372 793
rect 1326 721 1332 755
rect 1366 721 1372 755
rect 1326 683 1372 721
rect 1326 649 1332 683
rect 1366 649 1372 683
rect 1326 611 1372 649
rect 1326 577 1332 611
rect 1366 577 1372 611
rect 1326 539 1372 577
rect 1326 505 1332 539
rect 1366 505 1372 539
rect 1326 467 1372 505
rect 1326 433 1332 467
rect 1366 433 1372 467
rect 1326 395 1372 433
rect 1326 361 1332 395
rect 1366 361 1372 395
rect 1326 323 1372 361
rect 1326 289 1332 323
rect 1366 289 1372 323
rect 1326 251 1372 289
rect 1326 217 1332 251
rect 1366 217 1372 251
rect 1326 179 1372 217
rect 1326 145 1332 179
rect 1366 145 1372 179
rect 1326 107 1372 145
rect 1326 73 1332 107
rect 1366 73 1372 107
rect 1326 26 1372 73
rect 1414 1979 1460 2026
rect 1414 1945 1420 1979
rect 1454 1945 1460 1979
rect 1414 1907 1460 1945
rect 1414 1873 1420 1907
rect 1454 1873 1460 1907
rect 1414 1835 1460 1873
rect 1414 1801 1420 1835
rect 1454 1801 1460 1835
rect 1414 1763 1460 1801
rect 1414 1729 1420 1763
rect 1454 1729 1460 1763
rect 1414 1691 1460 1729
rect 1414 1657 1420 1691
rect 1454 1657 1460 1691
rect 1414 1619 1460 1657
rect 1414 1585 1420 1619
rect 1454 1585 1460 1619
rect 1414 1547 1460 1585
rect 1414 1513 1420 1547
rect 1454 1513 1460 1547
rect 1414 1475 1460 1513
rect 1414 1441 1420 1475
rect 1454 1441 1460 1475
rect 1414 1403 1460 1441
rect 1414 1369 1420 1403
rect 1454 1369 1460 1403
rect 1414 1331 1460 1369
rect 1414 1297 1420 1331
rect 1454 1297 1460 1331
rect 1414 1259 1460 1297
rect 1414 1225 1420 1259
rect 1454 1225 1460 1259
rect 1414 1187 1460 1225
rect 1414 1153 1420 1187
rect 1454 1153 1460 1187
rect 1414 1115 1460 1153
rect 1414 1081 1420 1115
rect 1454 1081 1460 1115
rect 1414 1043 1460 1081
rect 1414 1009 1420 1043
rect 1454 1009 1460 1043
rect 1414 971 1460 1009
rect 1414 937 1420 971
rect 1454 937 1460 971
rect 1414 899 1460 937
rect 1414 865 1420 899
rect 1454 865 1460 899
rect 1414 827 1460 865
rect 1414 793 1420 827
rect 1454 793 1460 827
rect 1414 755 1460 793
rect 1414 721 1420 755
rect 1454 721 1460 755
rect 1414 683 1460 721
rect 1414 649 1420 683
rect 1454 649 1460 683
rect 1414 611 1460 649
rect 1414 577 1420 611
rect 1454 577 1460 611
rect 1414 539 1460 577
rect 1414 505 1420 539
rect 1454 505 1460 539
rect 1414 467 1460 505
rect 1414 433 1420 467
rect 1454 433 1460 467
rect 1414 395 1460 433
rect 1414 361 1420 395
rect 1454 361 1460 395
rect 1414 323 1460 361
rect 1414 289 1420 323
rect 1454 289 1460 323
rect 1414 251 1460 289
rect 1414 217 1420 251
rect 1454 217 1460 251
rect 1414 179 1460 217
rect 1414 145 1420 179
rect 1454 145 1460 179
rect 1414 107 1460 145
rect 1414 73 1420 107
rect 1454 73 1460 107
rect 1414 26 1460 73
rect 1502 1979 1548 2026
rect 1502 1945 1508 1979
rect 1542 1945 1548 1979
rect 1502 1907 1548 1945
rect 1502 1873 1508 1907
rect 1542 1873 1548 1907
rect 1502 1835 1548 1873
rect 1502 1801 1508 1835
rect 1542 1801 1548 1835
rect 1502 1763 1548 1801
rect 1502 1729 1508 1763
rect 1542 1729 1548 1763
rect 1502 1691 1548 1729
rect 1502 1657 1508 1691
rect 1542 1657 1548 1691
rect 1502 1619 1548 1657
rect 1502 1585 1508 1619
rect 1542 1585 1548 1619
rect 1502 1547 1548 1585
rect 1502 1513 1508 1547
rect 1542 1513 1548 1547
rect 1502 1475 1548 1513
rect 1502 1441 1508 1475
rect 1542 1441 1548 1475
rect 1502 1403 1548 1441
rect 1502 1369 1508 1403
rect 1542 1369 1548 1403
rect 1502 1331 1548 1369
rect 1502 1297 1508 1331
rect 1542 1297 1548 1331
rect 1502 1259 1548 1297
rect 1502 1225 1508 1259
rect 1542 1225 1548 1259
rect 1502 1187 1548 1225
rect 1502 1153 1508 1187
rect 1542 1153 1548 1187
rect 1502 1115 1548 1153
rect 1502 1081 1508 1115
rect 1542 1081 1548 1115
rect 1502 1043 1548 1081
rect 1502 1009 1508 1043
rect 1542 1009 1548 1043
rect 1502 971 1548 1009
rect 1502 937 1508 971
rect 1542 937 1548 971
rect 1502 899 1548 937
rect 1502 865 1508 899
rect 1542 865 1548 899
rect 1502 827 1548 865
rect 1502 793 1508 827
rect 1542 793 1548 827
rect 1502 755 1548 793
rect 1502 721 1508 755
rect 1542 721 1548 755
rect 1502 683 1548 721
rect 1502 649 1508 683
rect 1542 649 1548 683
rect 1502 611 1548 649
rect 1502 577 1508 611
rect 1542 577 1548 611
rect 1502 539 1548 577
rect 1502 505 1508 539
rect 1542 505 1548 539
rect 1502 467 1548 505
rect 1502 433 1508 467
rect 1542 433 1548 467
rect 1502 395 1548 433
rect 1502 361 1508 395
rect 1542 361 1548 395
rect 1502 323 1548 361
rect 1502 289 1508 323
rect 1542 289 1548 323
rect 1502 251 1548 289
rect 1502 217 1508 251
rect 1542 217 1548 251
rect 1502 179 1548 217
rect 1502 145 1508 179
rect 1542 145 1548 179
rect 1502 107 1548 145
rect 1502 73 1508 107
rect 1542 73 1548 107
rect 1502 26 1548 73
rect 1590 1979 1636 2026
rect 1590 1945 1596 1979
rect 1630 1945 1636 1979
rect 1590 1907 1636 1945
rect 1590 1873 1596 1907
rect 1630 1873 1636 1907
rect 1590 1835 1636 1873
rect 1590 1801 1596 1835
rect 1630 1801 1636 1835
rect 1590 1763 1636 1801
rect 1590 1729 1596 1763
rect 1630 1729 1636 1763
rect 1590 1691 1636 1729
rect 1590 1657 1596 1691
rect 1630 1657 1636 1691
rect 1590 1619 1636 1657
rect 1590 1585 1596 1619
rect 1630 1585 1636 1619
rect 1590 1547 1636 1585
rect 1590 1513 1596 1547
rect 1630 1513 1636 1547
rect 1590 1475 1636 1513
rect 1590 1441 1596 1475
rect 1630 1441 1636 1475
rect 1590 1403 1636 1441
rect 1590 1369 1596 1403
rect 1630 1369 1636 1403
rect 1590 1331 1636 1369
rect 1590 1297 1596 1331
rect 1630 1297 1636 1331
rect 1590 1259 1636 1297
rect 1590 1225 1596 1259
rect 1630 1225 1636 1259
rect 1590 1187 1636 1225
rect 1590 1153 1596 1187
rect 1630 1153 1636 1187
rect 1590 1115 1636 1153
rect 1590 1081 1596 1115
rect 1630 1081 1636 1115
rect 1590 1043 1636 1081
rect 1590 1009 1596 1043
rect 1630 1009 1636 1043
rect 1590 971 1636 1009
rect 1590 937 1596 971
rect 1630 937 1636 971
rect 1590 899 1636 937
rect 1590 865 1596 899
rect 1630 865 1636 899
rect 1590 827 1636 865
rect 1590 793 1596 827
rect 1630 793 1636 827
rect 1590 755 1636 793
rect 1590 721 1596 755
rect 1630 721 1636 755
rect 1590 683 1636 721
rect 1590 649 1596 683
rect 1630 649 1636 683
rect 1590 611 1636 649
rect 1590 577 1596 611
rect 1630 577 1636 611
rect 1590 539 1636 577
rect 1590 505 1596 539
rect 1630 505 1636 539
rect 1590 467 1636 505
rect 1590 433 1596 467
rect 1630 433 1636 467
rect 1590 395 1636 433
rect 1590 361 1596 395
rect 1630 361 1636 395
rect 1590 323 1636 361
rect 1590 289 1596 323
rect 1630 289 1636 323
rect 1590 251 1636 289
rect 1590 217 1596 251
rect 1630 217 1636 251
rect 1590 179 1636 217
rect 1590 145 1596 179
rect 1630 145 1636 179
rect 1590 107 1636 145
rect 1590 73 1596 107
rect 1630 73 1636 107
rect 1590 26 1636 73
rect 1678 1979 1724 2026
rect 1678 1945 1684 1979
rect 1718 1945 1724 1979
rect 1678 1907 1724 1945
rect 1678 1873 1684 1907
rect 1718 1873 1724 1907
rect 1678 1835 1724 1873
rect 1678 1801 1684 1835
rect 1718 1801 1724 1835
rect 1678 1763 1724 1801
rect 1678 1729 1684 1763
rect 1718 1729 1724 1763
rect 1678 1691 1724 1729
rect 1678 1657 1684 1691
rect 1718 1657 1724 1691
rect 1678 1619 1724 1657
rect 1678 1585 1684 1619
rect 1718 1585 1724 1619
rect 1678 1547 1724 1585
rect 1678 1513 1684 1547
rect 1718 1513 1724 1547
rect 1678 1475 1724 1513
rect 1678 1441 1684 1475
rect 1718 1441 1724 1475
rect 1678 1403 1724 1441
rect 1678 1369 1684 1403
rect 1718 1369 1724 1403
rect 1678 1331 1724 1369
rect 1678 1297 1684 1331
rect 1718 1297 1724 1331
rect 1678 1259 1724 1297
rect 1678 1225 1684 1259
rect 1718 1225 1724 1259
rect 1678 1187 1724 1225
rect 1678 1153 1684 1187
rect 1718 1153 1724 1187
rect 1678 1115 1724 1153
rect 1678 1081 1684 1115
rect 1718 1081 1724 1115
rect 1678 1043 1724 1081
rect 1678 1009 1684 1043
rect 1718 1009 1724 1043
rect 1678 971 1724 1009
rect 1678 937 1684 971
rect 1718 937 1724 971
rect 1678 899 1724 937
rect 1678 865 1684 899
rect 1718 865 1724 899
rect 1678 827 1724 865
rect 1678 793 1684 827
rect 1718 793 1724 827
rect 1678 755 1724 793
rect 1678 721 1684 755
rect 1718 721 1724 755
rect 1678 683 1724 721
rect 1678 649 1684 683
rect 1718 649 1724 683
rect 1678 611 1724 649
rect 1678 577 1684 611
rect 1718 577 1724 611
rect 1678 539 1724 577
rect 1678 505 1684 539
rect 1718 505 1724 539
rect 1678 467 1724 505
rect 1678 433 1684 467
rect 1718 433 1724 467
rect 1678 395 1724 433
rect 1678 361 1684 395
rect 1718 361 1724 395
rect 1678 323 1724 361
rect 1678 289 1684 323
rect 1718 289 1724 323
rect 1678 251 1724 289
rect 1678 217 1684 251
rect 1718 217 1724 251
rect 1678 179 1724 217
rect 1678 145 1684 179
rect 1718 145 1724 179
rect 1678 107 1724 145
rect 1678 73 1684 107
rect 1718 73 1724 107
rect 1678 26 1724 73
rect 1766 1979 1812 2026
rect 1766 1945 1772 1979
rect 1806 1945 1812 1979
rect 1766 1907 1812 1945
rect 1766 1873 1772 1907
rect 1806 1873 1812 1907
rect 1766 1835 1812 1873
rect 1766 1801 1772 1835
rect 1806 1801 1812 1835
rect 1766 1763 1812 1801
rect 1766 1729 1772 1763
rect 1806 1729 1812 1763
rect 1766 1691 1812 1729
rect 1766 1657 1772 1691
rect 1806 1657 1812 1691
rect 1766 1619 1812 1657
rect 1766 1585 1772 1619
rect 1806 1585 1812 1619
rect 1766 1547 1812 1585
rect 1766 1513 1772 1547
rect 1806 1513 1812 1547
rect 1766 1475 1812 1513
rect 1766 1441 1772 1475
rect 1806 1441 1812 1475
rect 1766 1403 1812 1441
rect 1766 1369 1772 1403
rect 1806 1369 1812 1403
rect 1766 1331 1812 1369
rect 1766 1297 1772 1331
rect 1806 1297 1812 1331
rect 1766 1259 1812 1297
rect 1766 1225 1772 1259
rect 1806 1225 1812 1259
rect 1766 1187 1812 1225
rect 1766 1153 1772 1187
rect 1806 1153 1812 1187
rect 1766 1115 1812 1153
rect 1766 1081 1772 1115
rect 1806 1081 1812 1115
rect 1766 1043 1812 1081
rect 1766 1009 1772 1043
rect 1806 1009 1812 1043
rect 1766 971 1812 1009
rect 1766 937 1772 971
rect 1806 937 1812 971
rect 1766 899 1812 937
rect 1766 865 1772 899
rect 1806 865 1812 899
rect 1766 827 1812 865
rect 1766 793 1772 827
rect 1806 793 1812 827
rect 1766 755 1812 793
rect 1766 721 1772 755
rect 1806 721 1812 755
rect 1766 683 1812 721
rect 1766 649 1772 683
rect 1806 649 1812 683
rect 1766 611 1812 649
rect 1766 577 1772 611
rect 1806 577 1812 611
rect 1766 539 1812 577
rect 1766 505 1772 539
rect 1806 505 1812 539
rect 1766 467 1812 505
rect 1766 433 1772 467
rect 1806 433 1812 467
rect 1766 395 1812 433
rect 1766 361 1772 395
rect 1806 361 1812 395
rect 1766 323 1812 361
rect 1766 289 1772 323
rect 1806 289 1812 323
rect 1766 251 1812 289
rect 1766 217 1772 251
rect 1806 217 1812 251
rect 1766 179 1812 217
rect 1766 145 1772 179
rect 1806 145 1812 179
rect 1766 107 1812 145
rect 1766 73 1772 107
rect 1806 73 1812 107
rect 1766 26 1812 73
rect 1854 1979 1900 2026
rect 1854 1945 1860 1979
rect 1894 1945 1900 1979
rect 1854 1907 1900 1945
rect 1854 1873 1860 1907
rect 1894 1873 1900 1907
rect 1854 1835 1900 1873
rect 1854 1801 1860 1835
rect 1894 1801 1900 1835
rect 1854 1763 1900 1801
rect 1854 1729 1860 1763
rect 1894 1729 1900 1763
rect 1854 1691 1900 1729
rect 1854 1657 1860 1691
rect 1894 1657 1900 1691
rect 1854 1619 1900 1657
rect 1854 1585 1860 1619
rect 1894 1585 1900 1619
rect 1854 1547 1900 1585
rect 1854 1513 1860 1547
rect 1894 1513 1900 1547
rect 1854 1475 1900 1513
rect 1854 1441 1860 1475
rect 1894 1441 1900 1475
rect 1854 1403 1900 1441
rect 1854 1369 1860 1403
rect 1894 1369 1900 1403
rect 1854 1331 1900 1369
rect 1854 1297 1860 1331
rect 1894 1297 1900 1331
rect 1854 1259 1900 1297
rect 1854 1225 1860 1259
rect 1894 1225 1900 1259
rect 1854 1187 1900 1225
rect 1854 1153 1860 1187
rect 1894 1153 1900 1187
rect 1854 1115 1900 1153
rect 1854 1081 1860 1115
rect 1894 1081 1900 1115
rect 1854 1043 1900 1081
rect 1854 1009 1860 1043
rect 1894 1009 1900 1043
rect 1854 971 1900 1009
rect 1854 937 1860 971
rect 1894 937 1900 971
rect 1854 899 1900 937
rect 1854 865 1860 899
rect 1894 865 1900 899
rect 1854 827 1900 865
rect 1854 793 1860 827
rect 1894 793 1900 827
rect 1854 755 1900 793
rect 1854 721 1860 755
rect 1894 721 1900 755
rect 1854 683 1900 721
rect 1854 649 1860 683
rect 1894 649 1900 683
rect 1854 611 1900 649
rect 1854 577 1860 611
rect 1894 577 1900 611
rect 1854 539 1900 577
rect 1854 505 1860 539
rect 1894 505 1900 539
rect 1854 467 1900 505
rect 1854 433 1860 467
rect 1894 433 1900 467
rect 1854 395 1900 433
rect 1854 361 1860 395
rect 1894 361 1900 395
rect 1854 323 1900 361
rect 1854 289 1860 323
rect 1894 289 1900 323
rect 1854 251 1900 289
rect 1854 217 1860 251
rect 1894 217 1900 251
rect 1854 179 1900 217
rect 1854 145 1860 179
rect 1894 145 1900 179
rect 1854 107 1900 145
rect 1854 73 1860 107
rect 1894 73 1900 107
rect 1854 26 1900 73
rect 1942 1979 1988 2026
rect 1942 1945 1948 1979
rect 1982 1945 1988 1979
rect 1942 1907 1988 1945
rect 1942 1873 1948 1907
rect 1982 1873 1988 1907
rect 1942 1835 1988 1873
rect 1942 1801 1948 1835
rect 1982 1801 1988 1835
rect 1942 1763 1988 1801
rect 1942 1729 1948 1763
rect 1982 1729 1988 1763
rect 1942 1691 1988 1729
rect 1942 1657 1948 1691
rect 1982 1657 1988 1691
rect 1942 1619 1988 1657
rect 1942 1585 1948 1619
rect 1982 1585 1988 1619
rect 1942 1547 1988 1585
rect 1942 1513 1948 1547
rect 1982 1513 1988 1547
rect 1942 1475 1988 1513
rect 1942 1441 1948 1475
rect 1982 1441 1988 1475
rect 1942 1403 1988 1441
rect 1942 1369 1948 1403
rect 1982 1369 1988 1403
rect 1942 1331 1988 1369
rect 1942 1297 1948 1331
rect 1982 1297 1988 1331
rect 1942 1259 1988 1297
rect 1942 1225 1948 1259
rect 1982 1225 1988 1259
rect 1942 1187 1988 1225
rect 1942 1153 1948 1187
rect 1982 1153 1988 1187
rect 1942 1115 1988 1153
rect 1942 1081 1948 1115
rect 1982 1081 1988 1115
rect 1942 1043 1988 1081
rect 1942 1009 1948 1043
rect 1982 1009 1988 1043
rect 1942 971 1988 1009
rect 1942 937 1948 971
rect 1982 937 1988 971
rect 1942 899 1988 937
rect 1942 865 1948 899
rect 1982 865 1988 899
rect 1942 827 1988 865
rect 1942 793 1948 827
rect 1982 793 1988 827
rect 1942 755 1988 793
rect 1942 721 1948 755
rect 1982 721 1988 755
rect 1942 683 1988 721
rect 1942 649 1948 683
rect 1982 649 1988 683
rect 1942 611 1988 649
rect 1942 577 1948 611
rect 1982 577 1988 611
rect 1942 539 1988 577
rect 1942 505 1948 539
rect 1982 505 1988 539
rect 1942 467 1988 505
rect 1942 433 1948 467
rect 1982 433 1988 467
rect 1942 395 1988 433
rect 1942 361 1948 395
rect 1982 361 1988 395
rect 1942 323 1988 361
rect 1942 289 1948 323
rect 1982 289 1988 323
rect 1942 251 1988 289
rect 1942 217 1948 251
rect 1982 217 1988 251
rect 1942 179 1988 217
rect 1942 145 1948 179
rect 1982 145 1988 179
rect 1942 107 1988 145
rect 1942 73 1948 107
rect 1982 73 1988 107
rect 1942 26 1988 73
rect 2030 1979 2076 2026
rect 2030 1945 2036 1979
rect 2070 1945 2076 1979
rect 2030 1907 2076 1945
rect 2030 1873 2036 1907
rect 2070 1873 2076 1907
rect 2030 1835 2076 1873
rect 2030 1801 2036 1835
rect 2070 1801 2076 1835
rect 2030 1763 2076 1801
rect 2030 1729 2036 1763
rect 2070 1729 2076 1763
rect 2030 1691 2076 1729
rect 2030 1657 2036 1691
rect 2070 1657 2076 1691
rect 2030 1619 2076 1657
rect 2030 1585 2036 1619
rect 2070 1585 2076 1619
rect 2030 1547 2076 1585
rect 2030 1513 2036 1547
rect 2070 1513 2076 1547
rect 2030 1475 2076 1513
rect 2030 1441 2036 1475
rect 2070 1441 2076 1475
rect 2030 1403 2076 1441
rect 2030 1369 2036 1403
rect 2070 1369 2076 1403
rect 2030 1331 2076 1369
rect 2030 1297 2036 1331
rect 2070 1297 2076 1331
rect 2030 1259 2076 1297
rect 2030 1225 2036 1259
rect 2070 1225 2076 1259
rect 2030 1187 2076 1225
rect 2030 1153 2036 1187
rect 2070 1153 2076 1187
rect 2030 1115 2076 1153
rect 2030 1081 2036 1115
rect 2070 1081 2076 1115
rect 2030 1043 2076 1081
rect 2030 1009 2036 1043
rect 2070 1009 2076 1043
rect 2030 971 2076 1009
rect 2030 937 2036 971
rect 2070 937 2076 971
rect 2030 899 2076 937
rect 2030 865 2036 899
rect 2070 865 2076 899
rect 2030 827 2076 865
rect 2030 793 2036 827
rect 2070 793 2076 827
rect 2030 755 2076 793
rect 2030 721 2036 755
rect 2070 721 2076 755
rect 2030 683 2076 721
rect 2030 649 2036 683
rect 2070 649 2076 683
rect 2030 611 2076 649
rect 2030 577 2036 611
rect 2070 577 2076 611
rect 2030 539 2076 577
rect 2030 505 2036 539
rect 2070 505 2076 539
rect 2030 467 2076 505
rect 2030 433 2036 467
rect 2070 433 2076 467
rect 2030 395 2076 433
rect 2030 361 2036 395
rect 2070 361 2076 395
rect 2030 323 2076 361
rect 2030 289 2036 323
rect 2070 289 2076 323
rect 2030 251 2076 289
rect 2030 217 2036 251
rect 2070 217 2076 251
rect 2030 179 2076 217
rect 2030 145 2036 179
rect 2070 145 2076 179
rect 2030 107 2076 145
rect 2030 73 2036 107
rect 2070 73 2076 107
rect 2030 26 2076 73
rect 2118 1979 2164 2026
rect 2118 1945 2124 1979
rect 2158 1945 2164 1979
rect 2118 1907 2164 1945
rect 2118 1873 2124 1907
rect 2158 1873 2164 1907
rect 2118 1835 2164 1873
rect 2118 1801 2124 1835
rect 2158 1801 2164 1835
rect 2118 1763 2164 1801
rect 2118 1729 2124 1763
rect 2158 1729 2164 1763
rect 2118 1691 2164 1729
rect 2118 1657 2124 1691
rect 2158 1657 2164 1691
rect 2118 1619 2164 1657
rect 2118 1585 2124 1619
rect 2158 1585 2164 1619
rect 2118 1547 2164 1585
rect 2118 1513 2124 1547
rect 2158 1513 2164 1547
rect 2118 1475 2164 1513
rect 2118 1441 2124 1475
rect 2158 1441 2164 1475
rect 2118 1403 2164 1441
rect 2118 1369 2124 1403
rect 2158 1369 2164 1403
rect 2118 1331 2164 1369
rect 2118 1297 2124 1331
rect 2158 1297 2164 1331
rect 2118 1259 2164 1297
rect 2118 1225 2124 1259
rect 2158 1225 2164 1259
rect 2118 1187 2164 1225
rect 2118 1153 2124 1187
rect 2158 1153 2164 1187
rect 2118 1115 2164 1153
rect 2118 1081 2124 1115
rect 2158 1081 2164 1115
rect 2118 1043 2164 1081
rect 2118 1009 2124 1043
rect 2158 1009 2164 1043
rect 2118 971 2164 1009
rect 2118 937 2124 971
rect 2158 937 2164 971
rect 2118 899 2164 937
rect 2118 865 2124 899
rect 2158 865 2164 899
rect 2118 827 2164 865
rect 2118 793 2124 827
rect 2158 793 2164 827
rect 2118 755 2164 793
rect 2118 721 2124 755
rect 2158 721 2164 755
rect 2118 683 2164 721
rect 2118 649 2124 683
rect 2158 649 2164 683
rect 2118 611 2164 649
rect 2118 577 2124 611
rect 2158 577 2164 611
rect 2118 539 2164 577
rect 2118 505 2124 539
rect 2158 505 2164 539
rect 2118 467 2164 505
rect 2118 433 2124 467
rect 2158 433 2164 467
rect 2118 395 2164 433
rect 2118 361 2124 395
rect 2158 361 2164 395
rect 2118 323 2164 361
rect 2118 289 2124 323
rect 2158 289 2164 323
rect 2118 251 2164 289
rect 2118 217 2124 251
rect 2158 217 2164 251
rect 2118 179 2164 217
rect 2118 145 2124 179
rect 2158 145 2164 179
rect 2118 107 2164 145
rect 2118 73 2124 107
rect 2158 73 2164 107
rect 2118 26 2164 73
rect 2206 1979 2252 2026
rect 2206 1945 2212 1979
rect 2246 1945 2252 1979
rect 2206 1907 2252 1945
rect 2206 1873 2212 1907
rect 2246 1873 2252 1907
rect 2206 1835 2252 1873
rect 2206 1801 2212 1835
rect 2246 1801 2252 1835
rect 2206 1763 2252 1801
rect 2206 1729 2212 1763
rect 2246 1729 2252 1763
rect 2206 1691 2252 1729
rect 2206 1657 2212 1691
rect 2246 1657 2252 1691
rect 2206 1619 2252 1657
rect 2206 1585 2212 1619
rect 2246 1585 2252 1619
rect 2206 1547 2252 1585
rect 2206 1513 2212 1547
rect 2246 1513 2252 1547
rect 2206 1475 2252 1513
rect 2206 1441 2212 1475
rect 2246 1441 2252 1475
rect 2206 1403 2252 1441
rect 2206 1369 2212 1403
rect 2246 1369 2252 1403
rect 2206 1331 2252 1369
rect 2206 1297 2212 1331
rect 2246 1297 2252 1331
rect 2206 1259 2252 1297
rect 2206 1225 2212 1259
rect 2246 1225 2252 1259
rect 2206 1187 2252 1225
rect 2206 1153 2212 1187
rect 2246 1153 2252 1187
rect 2206 1115 2252 1153
rect 2206 1081 2212 1115
rect 2246 1081 2252 1115
rect 2206 1043 2252 1081
rect 2206 1009 2212 1043
rect 2246 1009 2252 1043
rect 2206 971 2252 1009
rect 2206 937 2212 971
rect 2246 937 2252 971
rect 2206 899 2252 937
rect 2206 865 2212 899
rect 2246 865 2252 899
rect 2206 827 2252 865
rect 2206 793 2212 827
rect 2246 793 2252 827
rect 2206 755 2252 793
rect 2206 721 2212 755
rect 2246 721 2252 755
rect 2206 683 2252 721
rect 2206 649 2212 683
rect 2246 649 2252 683
rect 2206 611 2252 649
rect 2206 577 2212 611
rect 2246 577 2252 611
rect 2206 539 2252 577
rect 2206 505 2212 539
rect 2246 505 2252 539
rect 2206 467 2252 505
rect 2206 433 2212 467
rect 2246 433 2252 467
rect 2206 395 2252 433
rect 2206 361 2212 395
rect 2246 361 2252 395
rect 2206 323 2252 361
rect 2206 289 2212 323
rect 2246 289 2252 323
rect 2206 251 2252 289
rect 2206 217 2212 251
rect 2246 217 2252 251
rect 2206 179 2252 217
rect 2206 145 2212 179
rect 2246 145 2252 179
rect 2206 107 2252 145
rect 2206 73 2212 107
rect 2246 73 2252 107
rect 2206 26 2252 73
rect 2294 1979 2340 2026
rect 2294 1945 2300 1979
rect 2334 1945 2340 1979
rect 2294 1907 2340 1945
rect 2294 1873 2300 1907
rect 2334 1873 2340 1907
rect 2294 1835 2340 1873
rect 2294 1801 2300 1835
rect 2334 1801 2340 1835
rect 2294 1763 2340 1801
rect 2294 1729 2300 1763
rect 2334 1729 2340 1763
rect 2294 1691 2340 1729
rect 2294 1657 2300 1691
rect 2334 1657 2340 1691
rect 2294 1619 2340 1657
rect 2294 1585 2300 1619
rect 2334 1585 2340 1619
rect 2294 1547 2340 1585
rect 2294 1513 2300 1547
rect 2334 1513 2340 1547
rect 2294 1475 2340 1513
rect 2294 1441 2300 1475
rect 2334 1441 2340 1475
rect 2294 1403 2340 1441
rect 2294 1369 2300 1403
rect 2334 1369 2340 1403
rect 2294 1331 2340 1369
rect 2294 1297 2300 1331
rect 2334 1297 2340 1331
rect 2294 1259 2340 1297
rect 2294 1225 2300 1259
rect 2334 1225 2340 1259
rect 2294 1187 2340 1225
rect 2294 1153 2300 1187
rect 2334 1153 2340 1187
rect 2294 1115 2340 1153
rect 2294 1081 2300 1115
rect 2334 1081 2340 1115
rect 2294 1043 2340 1081
rect 2294 1009 2300 1043
rect 2334 1009 2340 1043
rect 2294 971 2340 1009
rect 2294 937 2300 971
rect 2334 937 2340 971
rect 2294 899 2340 937
rect 2294 865 2300 899
rect 2334 865 2340 899
rect 2294 827 2340 865
rect 2294 793 2300 827
rect 2334 793 2340 827
rect 2294 755 2340 793
rect 2294 721 2300 755
rect 2334 721 2340 755
rect 2294 683 2340 721
rect 2294 649 2300 683
rect 2334 649 2340 683
rect 2294 611 2340 649
rect 2294 577 2300 611
rect 2334 577 2340 611
rect 2294 539 2340 577
rect 2294 505 2300 539
rect 2334 505 2340 539
rect 2294 467 2340 505
rect 2294 433 2300 467
rect 2334 433 2340 467
rect 2294 395 2340 433
rect 2294 361 2300 395
rect 2334 361 2340 395
rect 2294 323 2340 361
rect 2294 289 2300 323
rect 2334 289 2340 323
rect 2294 251 2340 289
rect 2294 217 2300 251
rect 2334 217 2340 251
rect 2294 179 2340 217
rect 2294 145 2300 179
rect 2334 145 2340 179
rect 2294 107 2340 145
rect 2294 73 2300 107
rect 2334 73 2340 107
rect 2294 26 2340 73
rect 2382 1979 2428 2026
rect 2382 1945 2388 1979
rect 2422 1945 2428 1979
rect 2382 1907 2428 1945
rect 2382 1873 2388 1907
rect 2422 1873 2428 1907
rect 2382 1835 2428 1873
rect 2382 1801 2388 1835
rect 2422 1801 2428 1835
rect 2382 1763 2428 1801
rect 2382 1729 2388 1763
rect 2422 1729 2428 1763
rect 2382 1691 2428 1729
rect 2382 1657 2388 1691
rect 2422 1657 2428 1691
rect 2382 1619 2428 1657
rect 2382 1585 2388 1619
rect 2422 1585 2428 1619
rect 2382 1547 2428 1585
rect 2382 1513 2388 1547
rect 2422 1513 2428 1547
rect 2382 1475 2428 1513
rect 2382 1441 2388 1475
rect 2422 1441 2428 1475
rect 2382 1403 2428 1441
rect 2382 1369 2388 1403
rect 2422 1369 2428 1403
rect 2382 1331 2428 1369
rect 2382 1297 2388 1331
rect 2422 1297 2428 1331
rect 2382 1259 2428 1297
rect 2382 1225 2388 1259
rect 2422 1225 2428 1259
rect 2382 1187 2428 1225
rect 2382 1153 2388 1187
rect 2422 1153 2428 1187
rect 2382 1115 2428 1153
rect 2382 1081 2388 1115
rect 2422 1081 2428 1115
rect 2382 1043 2428 1081
rect 2382 1009 2388 1043
rect 2422 1009 2428 1043
rect 2382 971 2428 1009
rect 2382 937 2388 971
rect 2422 937 2428 971
rect 2382 899 2428 937
rect 2382 865 2388 899
rect 2422 865 2428 899
rect 2382 827 2428 865
rect 2382 793 2388 827
rect 2422 793 2428 827
rect 2382 755 2428 793
rect 2382 721 2388 755
rect 2422 721 2428 755
rect 2382 683 2428 721
rect 2382 649 2388 683
rect 2422 649 2428 683
rect 2382 611 2428 649
rect 2382 577 2388 611
rect 2422 577 2428 611
rect 2382 539 2428 577
rect 2382 505 2388 539
rect 2422 505 2428 539
rect 2382 467 2428 505
rect 2382 433 2388 467
rect 2422 433 2428 467
rect 2382 395 2428 433
rect 2382 361 2388 395
rect 2422 361 2428 395
rect 2382 323 2428 361
rect 2382 289 2388 323
rect 2422 289 2428 323
rect 2382 251 2428 289
rect 2382 217 2388 251
rect 2422 217 2428 251
rect 2382 179 2428 217
rect 2382 145 2388 179
rect 2422 145 2428 179
rect 2382 107 2428 145
rect 2382 73 2388 107
rect 2422 73 2428 107
rect 2382 26 2428 73
rect 2470 1979 2516 2026
rect 2470 1945 2476 1979
rect 2510 1945 2516 1979
rect 2470 1907 2516 1945
rect 2470 1873 2476 1907
rect 2510 1873 2516 1907
rect 2470 1835 2516 1873
rect 2470 1801 2476 1835
rect 2510 1801 2516 1835
rect 2470 1763 2516 1801
rect 2470 1729 2476 1763
rect 2510 1729 2516 1763
rect 2470 1691 2516 1729
rect 2470 1657 2476 1691
rect 2510 1657 2516 1691
rect 2470 1619 2516 1657
rect 2470 1585 2476 1619
rect 2510 1585 2516 1619
rect 2470 1547 2516 1585
rect 2470 1513 2476 1547
rect 2510 1513 2516 1547
rect 2470 1475 2516 1513
rect 2470 1441 2476 1475
rect 2510 1441 2516 1475
rect 2470 1403 2516 1441
rect 2470 1369 2476 1403
rect 2510 1369 2516 1403
rect 2470 1331 2516 1369
rect 2470 1297 2476 1331
rect 2510 1297 2516 1331
rect 2470 1259 2516 1297
rect 2470 1225 2476 1259
rect 2510 1225 2516 1259
rect 2470 1187 2516 1225
rect 2470 1153 2476 1187
rect 2510 1153 2516 1187
rect 2470 1115 2516 1153
rect 2470 1081 2476 1115
rect 2510 1081 2516 1115
rect 2470 1043 2516 1081
rect 2470 1009 2476 1043
rect 2510 1009 2516 1043
rect 2470 971 2516 1009
rect 2470 937 2476 971
rect 2510 937 2516 971
rect 2470 899 2516 937
rect 2470 865 2476 899
rect 2510 865 2516 899
rect 2470 827 2516 865
rect 2470 793 2476 827
rect 2510 793 2516 827
rect 2470 755 2516 793
rect 2470 721 2476 755
rect 2510 721 2516 755
rect 2470 683 2516 721
rect 2470 649 2476 683
rect 2510 649 2516 683
rect 2470 611 2516 649
rect 2470 577 2476 611
rect 2510 577 2516 611
rect 2470 539 2516 577
rect 2470 505 2476 539
rect 2510 505 2516 539
rect 2470 467 2516 505
rect 2470 433 2476 467
rect 2510 433 2516 467
rect 2470 395 2516 433
rect 2470 361 2476 395
rect 2510 361 2516 395
rect 2470 323 2516 361
rect 2470 289 2476 323
rect 2510 289 2516 323
rect 2470 251 2516 289
rect 2470 217 2476 251
rect 2510 217 2516 251
rect 2470 179 2516 217
rect 2470 145 2476 179
rect 2510 145 2516 179
rect 2470 107 2516 145
rect 2470 73 2476 107
rect 2510 73 2516 107
rect 2470 26 2516 73
rect 2558 1979 2604 2026
rect 2558 1945 2564 1979
rect 2598 1945 2604 1979
rect 2558 1907 2604 1945
rect 2558 1873 2564 1907
rect 2598 1873 2604 1907
rect 2558 1835 2604 1873
rect 2558 1801 2564 1835
rect 2598 1801 2604 1835
rect 2558 1763 2604 1801
rect 2558 1729 2564 1763
rect 2598 1729 2604 1763
rect 2558 1691 2604 1729
rect 2558 1657 2564 1691
rect 2598 1657 2604 1691
rect 2558 1619 2604 1657
rect 2558 1585 2564 1619
rect 2598 1585 2604 1619
rect 2558 1547 2604 1585
rect 2558 1513 2564 1547
rect 2598 1513 2604 1547
rect 2558 1475 2604 1513
rect 2558 1441 2564 1475
rect 2598 1441 2604 1475
rect 2558 1403 2604 1441
rect 2558 1369 2564 1403
rect 2598 1369 2604 1403
rect 2558 1331 2604 1369
rect 2558 1297 2564 1331
rect 2598 1297 2604 1331
rect 2558 1259 2604 1297
rect 2558 1225 2564 1259
rect 2598 1225 2604 1259
rect 2558 1187 2604 1225
rect 2558 1153 2564 1187
rect 2598 1153 2604 1187
rect 2558 1115 2604 1153
rect 2558 1081 2564 1115
rect 2598 1081 2604 1115
rect 2558 1043 2604 1081
rect 2558 1009 2564 1043
rect 2598 1009 2604 1043
rect 2558 971 2604 1009
rect 2558 937 2564 971
rect 2598 937 2604 971
rect 2558 899 2604 937
rect 2558 865 2564 899
rect 2598 865 2604 899
rect 2558 827 2604 865
rect 2558 793 2564 827
rect 2598 793 2604 827
rect 2558 755 2604 793
rect 2558 721 2564 755
rect 2598 721 2604 755
rect 2558 683 2604 721
rect 2558 649 2564 683
rect 2598 649 2604 683
rect 2558 611 2604 649
rect 2558 577 2564 611
rect 2598 577 2604 611
rect 2558 539 2604 577
rect 2558 505 2564 539
rect 2598 505 2604 539
rect 2558 467 2604 505
rect 2558 433 2564 467
rect 2598 433 2604 467
rect 2558 395 2604 433
rect 2558 361 2564 395
rect 2598 361 2604 395
rect 2558 323 2604 361
rect 2558 289 2564 323
rect 2598 289 2604 323
rect 2558 251 2604 289
rect 2558 217 2564 251
rect 2598 217 2604 251
rect 2558 179 2604 217
rect 2558 145 2564 179
rect 2598 145 2604 179
rect 2558 107 2604 145
rect 2558 73 2564 107
rect 2598 73 2604 107
rect 2558 26 2604 73
rect 2646 1979 2692 2026
rect 2646 1945 2652 1979
rect 2686 1945 2692 1979
rect 2646 1907 2692 1945
rect 2646 1873 2652 1907
rect 2686 1873 2692 1907
rect 2646 1835 2692 1873
rect 2646 1801 2652 1835
rect 2686 1801 2692 1835
rect 2646 1763 2692 1801
rect 2646 1729 2652 1763
rect 2686 1729 2692 1763
rect 2646 1691 2692 1729
rect 2646 1657 2652 1691
rect 2686 1657 2692 1691
rect 2646 1619 2692 1657
rect 2646 1585 2652 1619
rect 2686 1585 2692 1619
rect 2646 1547 2692 1585
rect 2646 1513 2652 1547
rect 2686 1513 2692 1547
rect 2646 1475 2692 1513
rect 2646 1441 2652 1475
rect 2686 1441 2692 1475
rect 2646 1403 2692 1441
rect 2646 1369 2652 1403
rect 2686 1369 2692 1403
rect 2646 1331 2692 1369
rect 2646 1297 2652 1331
rect 2686 1297 2692 1331
rect 2646 1259 2692 1297
rect 2646 1225 2652 1259
rect 2686 1225 2692 1259
rect 2646 1187 2692 1225
rect 2646 1153 2652 1187
rect 2686 1153 2692 1187
rect 2646 1115 2692 1153
rect 2646 1081 2652 1115
rect 2686 1081 2692 1115
rect 2646 1043 2692 1081
rect 2646 1009 2652 1043
rect 2686 1009 2692 1043
rect 2646 971 2692 1009
rect 2646 937 2652 971
rect 2686 937 2692 971
rect 2646 899 2692 937
rect 2646 865 2652 899
rect 2686 865 2692 899
rect 2646 827 2692 865
rect 2646 793 2652 827
rect 2686 793 2692 827
rect 2646 755 2692 793
rect 2646 721 2652 755
rect 2686 721 2692 755
rect 2646 683 2692 721
rect 2646 649 2652 683
rect 2686 649 2692 683
rect 2646 611 2692 649
rect 2646 577 2652 611
rect 2686 577 2692 611
rect 2646 539 2692 577
rect 2646 505 2652 539
rect 2686 505 2692 539
rect 2646 467 2692 505
rect 2646 433 2652 467
rect 2686 433 2692 467
rect 2646 395 2692 433
rect 2646 361 2652 395
rect 2686 361 2692 395
rect 2646 323 2692 361
rect 2646 289 2652 323
rect 2686 289 2692 323
rect 2646 251 2692 289
rect 2646 217 2652 251
rect 2686 217 2692 251
rect 2646 179 2692 217
rect 2646 145 2652 179
rect 2686 145 2692 179
rect 2646 107 2692 145
rect 2646 73 2652 107
rect 2686 73 2692 107
rect 2646 26 2692 73
rect -773 -58 2112 -14
rect -773 -92 628 -58
rect 662 -92 980 -58
rect 1014 -92 1332 -58
rect 1366 -92 1684 -58
rect 1718 -92 2036 -58
rect 2070 -92 2112 -58
rect -773 -136 2112 -92
rect 2346 -58 2640 -14
rect 2346 -92 2388 -58
rect 2422 -92 2564 -58
rect 2598 -92 2640 -58
rect 2346 -136 2640 -92
rect 2346 -164 2464 -136
rect 48 -211 2464 -164
rect 48 -245 96 -211
rect 130 -245 168 -211
rect 202 -245 240 -211
rect 274 -245 312 -211
rect 346 -245 384 -211
rect 418 -245 456 -211
rect 490 -222 2464 -211
rect 490 -245 804 -222
rect 48 -256 804 -245
rect 838 -256 1156 -222
rect 1190 -256 1508 -222
rect 1542 -256 1860 -222
rect 1894 -256 2212 -222
rect 2246 -256 2464 -222
rect 48 -299 2464 -256
rect 48 -301 2346 -299
rect 48 -302 608 -301
use sky130_fd_pr__nfet_01v8_lvt_9WNFGV  sky130_fd_pr__nfet_01v8_lvt_9WNFGV_0
timestamp 1637060811
transform 1 0 73 0 1 1026
box -99 -1026 99 1026
<< labels >>
rlabel metal1 s 1492 2396 1492 2396 4 D2
port 1 nsew
rlabel metal1 s 1485 2291 1485 2291 4 S1
port 2 nsew
rlabel metal1 s 1349 -301 1349 -301 4 G2
port 3 nsew
rlabel metal1 s 1435 -136 1435 -136 4 G1
port 4 nsew
<< end >>
