magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< locali >>
rect 18272 22242 18538 22348
rect 18272 22136 18340 22242
rect 18446 22136 18538 22242
rect 18272 22048 18538 22136
rect 18490 20974 18668 21012
rect 18490 20940 18546 20974
rect 18580 20940 18668 20974
rect 18490 20902 18668 20940
rect 18490 20868 18546 20902
rect 18580 20868 18668 20902
rect 18490 20846 18668 20868
<< viali >>
rect 18340 22136 18446 22242
rect 18546 20940 18580 20974
rect 18546 20868 18580 20902
<< metal1 >>
rect 18272 22242 18538 22348
rect 18272 22136 18340 22242
rect 18446 22136 18538 22242
rect 18272 22048 18538 22136
rect 20464 21232 20838 22156
rect 25816 21116 26320 22228
rect 30742 21182 31106 22222
rect 18490 20974 18668 21012
rect 18490 20947 18546 20974
rect 18580 20947 18668 20974
rect 18490 20895 18537 20947
rect 18589 20895 18668 20947
rect 18490 20868 18546 20895
rect 18580 20868 18668 20895
rect 18490 20846 18668 20868
<< via1 >>
rect 18537 20940 18546 20947
rect 18546 20940 18580 20947
rect 18580 20940 18589 20947
rect 18537 20902 18589 20940
rect 18537 20895 18546 20902
rect 18546 20895 18580 20902
rect 18580 20895 18589 20902
<< metal2 >>
rect 17276 38148 18560 38378
rect 36786 22436 38266 22442
rect 36662 22379 38266 22436
rect 36662 22243 37833 22379
rect 38209 22243 38266 22379
rect 36662 22178 38266 22243
rect 18490 20947 18668 21012
rect 18490 20895 18537 20947
rect 18589 20895 18668 20947
rect 18490 20846 18668 20895
rect 36662 20830 37170 22178
rect 17242 4246 40488 4350
rect 17242 4030 39594 4246
rect 40290 4030 40488 4246
rect 17242 3944 40488 4030
<< via2 >>
rect 37833 22243 38209 22379
rect 39594 4030 40290 4246
<< metal3 >>
rect 37780 22383 38272 22442
rect 37780 22239 37829 22383
rect 38213 22239 38272 22383
rect 37780 22172 38272 22239
rect 39562 4246 40322 4262
rect 39562 4030 39594 4246
rect 40290 4030 40322 4246
rect 39562 4014 40322 4030
<< via3 >>
rect 37829 22379 38213 22383
rect 37829 22243 37833 22379
rect 37833 22243 38209 22379
rect 38209 22243 38213 22379
rect 37829 22239 38213 22243
<< metal4 >>
rect 39350 22486 42378 22966
rect 37780 22383 42378 22486
rect 37780 22239 37829 22383
rect 38213 22239 42378 22383
rect 37780 22156 42378 22239
rect 39290 21656 42378 22156
use pmos40  pmos40_0
timestamp 1636132012
transform 1 0 18406 0 -1 21364
box 0 0 18908 16664
use pmos40  pmos40_1
timestamp 1636132012
transform 1 0 18280 0 -1 38724
box 0 0 18908 16664
use cap225_layout  cap225_layout_0
timestamp 1636132012
transform 1 0 129394 0 1 89866
box -90032 -89592 7438 8920
use recitifer_layout  recitifer_layout_0
timestamp 1636132012
transform 1 0 930 0 1 29318
box -910 -29318 17472 9474
<< labels >>
rlabel metal1 s 26132 21614 26132 21614 4 VOUT_C
port 1 nsew
rlabel metal2 s 38716 4124 38716 4124 4 VSS
port 2 nsew
rlabel metal2 s 18060 38258 18060 38258 4 VIN1
port 3 nsew
rlabel metal4 s 38484 22386 38484 22386 4 VIN2
port 4 nsew
<< end >>
