magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< locali >>
rect 32542 2293 39918 2352
rect 32542 2115 39500 2293
rect 39822 2115 39918 2293
rect 32542 2056 39918 2115
<< viali >>
rect 39500 2115 39822 2293
<< metal1 >>
rect 18072 2496 22216 2592
rect 18072 2188 18168 2496
rect 18348 2188 22216 2496
rect 18072 2102 22216 2188
rect 33624 1654 33908 4786
rect 39350 2294 39912 2344
rect 39350 2293 39507 2294
rect 39815 2293 39912 2294
rect 39350 2115 39500 2293
rect 39822 2115 39912 2293
rect 39350 2114 39507 2115
rect 39815 2114 39912 2115
rect 39350 2058 39912 2114
rect 33274 1650 34032 1654
rect 33274 1470 33407 1650
rect 33971 1470 34032 1650
rect 33274 1418 34032 1470
rect 33274 1378 33954 1418
<< via1 >>
rect 18168 2188 18348 2496
rect 39507 2293 39815 2294
rect 39507 2115 39815 2293
rect 39507 2114 39815 2115
rect 33407 1470 33971 1650
<< metal2 >>
rect 18160 38322 18366 38332
rect 18160 38186 18195 38322
rect 18331 38186 18366 38322
rect 18160 38176 18366 38186
rect 18052 2496 18418 2588
rect 18052 2188 18168 2496
rect 18348 2188 18418 2496
rect 18052 2096 18418 2188
rect 39350 2294 39912 2344
rect 39350 2114 39507 2294
rect 39815 2114 39912 2294
rect 39350 2058 39912 2114
rect 30098 1650 34060 1704
rect 30098 1470 33407 1650
rect 33971 1470 34060 1650
rect 30098 1384 34060 1470
rect 27588 707 33540 794
rect 27588 411 33241 707
rect 33457 411 33540 707
rect 27588 354 33540 411
<< via2 >>
rect 18195 38186 18331 38322
rect 18190 2194 18326 2490
rect 39513 2136 39809 2272
rect 33241 411 33457 707
<< metal3 >>
rect 18076 38322 18422 38364
rect 18076 38186 18195 38322
rect 18331 38186 18422 38322
rect 18076 2490 18422 38186
rect 18076 2194 18190 2490
rect 18326 2194 18422 2490
rect 18076 2102 18422 2194
rect 39476 2272 39846 2300
rect 39476 2136 39513 2272
rect 39809 2136 39846 2272
rect 39476 2108 39846 2136
rect 33154 711 33608 848
rect 33154 407 33237 711
rect 33461 407 33608 711
rect 33154 252 33608 407
<< via3 >>
rect 33237 707 33461 711
rect 33237 411 33241 707
rect 33241 411 33457 707
rect 33457 411 33461 707
rect 33237 407 33461 411
<< metal4 >>
rect 42048 854 43364 3186
rect 33190 711 43364 854
rect 33190 407 33237 711
rect 33461 407 43364 711
rect 33190 272 43364 407
use RX_layout  RX_layout_0
timestamp 1636132012
transform 1 0 -22 0 1 -2
box 20 0 136832 98786
use Comparator_jafar  Comparator_jafar_0
timestamp 1636132012
transform 1 0 18424 0 1 634
box 3752 -276 14192 2976
<< end >>
