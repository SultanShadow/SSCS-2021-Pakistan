magic
tech sky130A
magscale 1 2
timestamp 1635855079
<< error_p >>
rect -317 572 -259 578
rect -125 572 -67 578
rect 67 572 125 578
rect 259 572 317 578
rect -317 538 -305 572
rect -125 538 -113 572
rect 67 538 79 572
rect 259 538 271 572
rect -317 532 -259 538
rect -125 532 -67 538
rect 67 532 125 538
rect 259 532 317 538
rect -413 -538 -355 -532
rect -221 -538 -163 -532
rect -29 -538 29 -532
rect 163 -538 221 -532
rect 355 -538 413 -532
rect -413 -572 -401 -538
rect -221 -572 -209 -538
rect -29 -572 -17 -538
rect 163 -572 175 -538
rect 355 -572 367 -538
rect -413 -578 -355 -572
rect -221 -578 -163 -572
rect -29 -578 29 -572
rect 163 -578 221 -572
rect 355 -578 413 -572
<< pwell >>
rect -589 -700 589 700
<< nmoslvt >>
rect -399 -500 -369 500
rect -303 -500 -273 500
rect -207 -500 -177 500
rect -111 -500 -81 500
rect -15 -500 15 500
rect 81 -500 111 500
rect 177 -500 207 500
rect 273 -500 303 500
rect 369 -500 399 500
<< ndiff >>
rect -461 459 -399 500
rect -461 425 -449 459
rect -415 425 -399 459
rect -461 391 -399 425
rect -461 357 -449 391
rect -415 357 -399 391
rect -461 323 -399 357
rect -461 289 -449 323
rect -415 289 -399 323
rect -461 255 -399 289
rect -461 221 -449 255
rect -415 221 -399 255
rect -461 187 -399 221
rect -461 153 -449 187
rect -415 153 -399 187
rect -461 119 -399 153
rect -461 85 -449 119
rect -415 85 -399 119
rect -461 51 -399 85
rect -461 17 -449 51
rect -415 17 -399 51
rect -461 -17 -399 17
rect -461 -51 -449 -17
rect -415 -51 -399 -17
rect -461 -85 -399 -51
rect -461 -119 -449 -85
rect -415 -119 -399 -85
rect -461 -153 -399 -119
rect -461 -187 -449 -153
rect -415 -187 -399 -153
rect -461 -221 -399 -187
rect -461 -255 -449 -221
rect -415 -255 -399 -221
rect -461 -289 -399 -255
rect -461 -323 -449 -289
rect -415 -323 -399 -289
rect -461 -357 -399 -323
rect -461 -391 -449 -357
rect -415 -391 -399 -357
rect -461 -425 -399 -391
rect -461 -459 -449 -425
rect -415 -459 -399 -425
rect -461 -500 -399 -459
rect -369 459 -303 500
rect -369 425 -353 459
rect -319 425 -303 459
rect -369 391 -303 425
rect -369 357 -353 391
rect -319 357 -303 391
rect -369 323 -303 357
rect -369 289 -353 323
rect -319 289 -303 323
rect -369 255 -303 289
rect -369 221 -353 255
rect -319 221 -303 255
rect -369 187 -303 221
rect -369 153 -353 187
rect -319 153 -303 187
rect -369 119 -303 153
rect -369 85 -353 119
rect -319 85 -303 119
rect -369 51 -303 85
rect -369 17 -353 51
rect -319 17 -303 51
rect -369 -17 -303 17
rect -369 -51 -353 -17
rect -319 -51 -303 -17
rect -369 -85 -303 -51
rect -369 -119 -353 -85
rect -319 -119 -303 -85
rect -369 -153 -303 -119
rect -369 -187 -353 -153
rect -319 -187 -303 -153
rect -369 -221 -303 -187
rect -369 -255 -353 -221
rect -319 -255 -303 -221
rect -369 -289 -303 -255
rect -369 -323 -353 -289
rect -319 -323 -303 -289
rect -369 -357 -303 -323
rect -369 -391 -353 -357
rect -319 -391 -303 -357
rect -369 -425 -303 -391
rect -369 -459 -353 -425
rect -319 -459 -303 -425
rect -369 -500 -303 -459
rect -273 459 -207 500
rect -273 425 -257 459
rect -223 425 -207 459
rect -273 391 -207 425
rect -273 357 -257 391
rect -223 357 -207 391
rect -273 323 -207 357
rect -273 289 -257 323
rect -223 289 -207 323
rect -273 255 -207 289
rect -273 221 -257 255
rect -223 221 -207 255
rect -273 187 -207 221
rect -273 153 -257 187
rect -223 153 -207 187
rect -273 119 -207 153
rect -273 85 -257 119
rect -223 85 -207 119
rect -273 51 -207 85
rect -273 17 -257 51
rect -223 17 -207 51
rect -273 -17 -207 17
rect -273 -51 -257 -17
rect -223 -51 -207 -17
rect -273 -85 -207 -51
rect -273 -119 -257 -85
rect -223 -119 -207 -85
rect -273 -153 -207 -119
rect -273 -187 -257 -153
rect -223 -187 -207 -153
rect -273 -221 -207 -187
rect -273 -255 -257 -221
rect -223 -255 -207 -221
rect -273 -289 -207 -255
rect -273 -323 -257 -289
rect -223 -323 -207 -289
rect -273 -357 -207 -323
rect -273 -391 -257 -357
rect -223 -391 -207 -357
rect -273 -425 -207 -391
rect -273 -459 -257 -425
rect -223 -459 -207 -425
rect -273 -500 -207 -459
rect -177 459 -111 500
rect -177 425 -161 459
rect -127 425 -111 459
rect -177 391 -111 425
rect -177 357 -161 391
rect -127 357 -111 391
rect -177 323 -111 357
rect -177 289 -161 323
rect -127 289 -111 323
rect -177 255 -111 289
rect -177 221 -161 255
rect -127 221 -111 255
rect -177 187 -111 221
rect -177 153 -161 187
rect -127 153 -111 187
rect -177 119 -111 153
rect -177 85 -161 119
rect -127 85 -111 119
rect -177 51 -111 85
rect -177 17 -161 51
rect -127 17 -111 51
rect -177 -17 -111 17
rect -177 -51 -161 -17
rect -127 -51 -111 -17
rect -177 -85 -111 -51
rect -177 -119 -161 -85
rect -127 -119 -111 -85
rect -177 -153 -111 -119
rect -177 -187 -161 -153
rect -127 -187 -111 -153
rect -177 -221 -111 -187
rect -177 -255 -161 -221
rect -127 -255 -111 -221
rect -177 -289 -111 -255
rect -177 -323 -161 -289
rect -127 -323 -111 -289
rect -177 -357 -111 -323
rect -177 -391 -161 -357
rect -127 -391 -111 -357
rect -177 -425 -111 -391
rect -177 -459 -161 -425
rect -127 -459 -111 -425
rect -177 -500 -111 -459
rect -81 459 -15 500
rect -81 425 -65 459
rect -31 425 -15 459
rect -81 391 -15 425
rect -81 357 -65 391
rect -31 357 -15 391
rect -81 323 -15 357
rect -81 289 -65 323
rect -31 289 -15 323
rect -81 255 -15 289
rect -81 221 -65 255
rect -31 221 -15 255
rect -81 187 -15 221
rect -81 153 -65 187
rect -31 153 -15 187
rect -81 119 -15 153
rect -81 85 -65 119
rect -31 85 -15 119
rect -81 51 -15 85
rect -81 17 -65 51
rect -31 17 -15 51
rect -81 -17 -15 17
rect -81 -51 -65 -17
rect -31 -51 -15 -17
rect -81 -85 -15 -51
rect -81 -119 -65 -85
rect -31 -119 -15 -85
rect -81 -153 -15 -119
rect -81 -187 -65 -153
rect -31 -187 -15 -153
rect -81 -221 -15 -187
rect -81 -255 -65 -221
rect -31 -255 -15 -221
rect -81 -289 -15 -255
rect -81 -323 -65 -289
rect -31 -323 -15 -289
rect -81 -357 -15 -323
rect -81 -391 -65 -357
rect -31 -391 -15 -357
rect -81 -425 -15 -391
rect -81 -459 -65 -425
rect -31 -459 -15 -425
rect -81 -500 -15 -459
rect 15 459 81 500
rect 15 425 31 459
rect 65 425 81 459
rect 15 391 81 425
rect 15 357 31 391
rect 65 357 81 391
rect 15 323 81 357
rect 15 289 31 323
rect 65 289 81 323
rect 15 255 81 289
rect 15 221 31 255
rect 65 221 81 255
rect 15 187 81 221
rect 15 153 31 187
rect 65 153 81 187
rect 15 119 81 153
rect 15 85 31 119
rect 65 85 81 119
rect 15 51 81 85
rect 15 17 31 51
rect 65 17 81 51
rect 15 -17 81 17
rect 15 -51 31 -17
rect 65 -51 81 -17
rect 15 -85 81 -51
rect 15 -119 31 -85
rect 65 -119 81 -85
rect 15 -153 81 -119
rect 15 -187 31 -153
rect 65 -187 81 -153
rect 15 -221 81 -187
rect 15 -255 31 -221
rect 65 -255 81 -221
rect 15 -289 81 -255
rect 15 -323 31 -289
rect 65 -323 81 -289
rect 15 -357 81 -323
rect 15 -391 31 -357
rect 65 -391 81 -357
rect 15 -425 81 -391
rect 15 -459 31 -425
rect 65 -459 81 -425
rect 15 -500 81 -459
rect 111 459 177 500
rect 111 425 127 459
rect 161 425 177 459
rect 111 391 177 425
rect 111 357 127 391
rect 161 357 177 391
rect 111 323 177 357
rect 111 289 127 323
rect 161 289 177 323
rect 111 255 177 289
rect 111 221 127 255
rect 161 221 177 255
rect 111 187 177 221
rect 111 153 127 187
rect 161 153 177 187
rect 111 119 177 153
rect 111 85 127 119
rect 161 85 177 119
rect 111 51 177 85
rect 111 17 127 51
rect 161 17 177 51
rect 111 -17 177 17
rect 111 -51 127 -17
rect 161 -51 177 -17
rect 111 -85 177 -51
rect 111 -119 127 -85
rect 161 -119 177 -85
rect 111 -153 177 -119
rect 111 -187 127 -153
rect 161 -187 177 -153
rect 111 -221 177 -187
rect 111 -255 127 -221
rect 161 -255 177 -221
rect 111 -289 177 -255
rect 111 -323 127 -289
rect 161 -323 177 -289
rect 111 -357 177 -323
rect 111 -391 127 -357
rect 161 -391 177 -357
rect 111 -425 177 -391
rect 111 -459 127 -425
rect 161 -459 177 -425
rect 111 -500 177 -459
rect 207 459 273 500
rect 207 425 223 459
rect 257 425 273 459
rect 207 391 273 425
rect 207 357 223 391
rect 257 357 273 391
rect 207 323 273 357
rect 207 289 223 323
rect 257 289 273 323
rect 207 255 273 289
rect 207 221 223 255
rect 257 221 273 255
rect 207 187 273 221
rect 207 153 223 187
rect 257 153 273 187
rect 207 119 273 153
rect 207 85 223 119
rect 257 85 273 119
rect 207 51 273 85
rect 207 17 223 51
rect 257 17 273 51
rect 207 -17 273 17
rect 207 -51 223 -17
rect 257 -51 273 -17
rect 207 -85 273 -51
rect 207 -119 223 -85
rect 257 -119 273 -85
rect 207 -153 273 -119
rect 207 -187 223 -153
rect 257 -187 273 -153
rect 207 -221 273 -187
rect 207 -255 223 -221
rect 257 -255 273 -221
rect 207 -289 273 -255
rect 207 -323 223 -289
rect 257 -323 273 -289
rect 207 -357 273 -323
rect 207 -391 223 -357
rect 257 -391 273 -357
rect 207 -425 273 -391
rect 207 -459 223 -425
rect 257 -459 273 -425
rect 207 -500 273 -459
rect 303 459 369 500
rect 303 425 319 459
rect 353 425 369 459
rect 303 391 369 425
rect 303 357 319 391
rect 353 357 369 391
rect 303 323 369 357
rect 303 289 319 323
rect 353 289 369 323
rect 303 255 369 289
rect 303 221 319 255
rect 353 221 369 255
rect 303 187 369 221
rect 303 153 319 187
rect 353 153 369 187
rect 303 119 369 153
rect 303 85 319 119
rect 353 85 369 119
rect 303 51 369 85
rect 303 17 319 51
rect 353 17 369 51
rect 303 -17 369 17
rect 303 -51 319 -17
rect 353 -51 369 -17
rect 303 -85 369 -51
rect 303 -119 319 -85
rect 353 -119 369 -85
rect 303 -153 369 -119
rect 303 -187 319 -153
rect 353 -187 369 -153
rect 303 -221 369 -187
rect 303 -255 319 -221
rect 353 -255 369 -221
rect 303 -289 369 -255
rect 303 -323 319 -289
rect 353 -323 369 -289
rect 303 -357 369 -323
rect 303 -391 319 -357
rect 353 -391 369 -357
rect 303 -425 369 -391
rect 303 -459 319 -425
rect 353 -459 369 -425
rect 303 -500 369 -459
rect 399 459 461 500
rect 399 425 415 459
rect 449 425 461 459
rect 399 391 461 425
rect 399 357 415 391
rect 449 357 461 391
rect 399 323 461 357
rect 399 289 415 323
rect 449 289 461 323
rect 399 255 461 289
rect 399 221 415 255
rect 449 221 461 255
rect 399 187 461 221
rect 399 153 415 187
rect 449 153 461 187
rect 399 119 461 153
rect 399 85 415 119
rect 449 85 461 119
rect 399 51 461 85
rect 399 17 415 51
rect 449 17 461 51
rect 399 -17 461 17
rect 399 -51 415 -17
rect 449 -51 461 -17
rect 399 -85 461 -51
rect 399 -119 415 -85
rect 449 -119 461 -85
rect 399 -153 461 -119
rect 399 -187 415 -153
rect 449 -187 461 -153
rect 399 -221 461 -187
rect 399 -255 415 -221
rect 449 -255 461 -221
rect 399 -289 461 -255
rect 399 -323 415 -289
rect 449 -323 461 -289
rect 399 -357 461 -323
rect 399 -391 415 -357
rect 449 -391 461 -357
rect 399 -425 461 -391
rect 399 -459 415 -425
rect 449 -459 461 -425
rect 399 -500 461 -459
<< ndiffc >>
rect -449 425 -415 459
rect -449 357 -415 391
rect -449 289 -415 323
rect -449 221 -415 255
rect -449 153 -415 187
rect -449 85 -415 119
rect -449 17 -415 51
rect -449 -51 -415 -17
rect -449 -119 -415 -85
rect -449 -187 -415 -153
rect -449 -255 -415 -221
rect -449 -323 -415 -289
rect -449 -391 -415 -357
rect -449 -459 -415 -425
rect -353 425 -319 459
rect -353 357 -319 391
rect -353 289 -319 323
rect -353 221 -319 255
rect -353 153 -319 187
rect -353 85 -319 119
rect -353 17 -319 51
rect -353 -51 -319 -17
rect -353 -119 -319 -85
rect -353 -187 -319 -153
rect -353 -255 -319 -221
rect -353 -323 -319 -289
rect -353 -391 -319 -357
rect -353 -459 -319 -425
rect -257 425 -223 459
rect -257 357 -223 391
rect -257 289 -223 323
rect -257 221 -223 255
rect -257 153 -223 187
rect -257 85 -223 119
rect -257 17 -223 51
rect -257 -51 -223 -17
rect -257 -119 -223 -85
rect -257 -187 -223 -153
rect -257 -255 -223 -221
rect -257 -323 -223 -289
rect -257 -391 -223 -357
rect -257 -459 -223 -425
rect -161 425 -127 459
rect -161 357 -127 391
rect -161 289 -127 323
rect -161 221 -127 255
rect -161 153 -127 187
rect -161 85 -127 119
rect -161 17 -127 51
rect -161 -51 -127 -17
rect -161 -119 -127 -85
rect -161 -187 -127 -153
rect -161 -255 -127 -221
rect -161 -323 -127 -289
rect -161 -391 -127 -357
rect -161 -459 -127 -425
rect -65 425 -31 459
rect -65 357 -31 391
rect -65 289 -31 323
rect -65 221 -31 255
rect -65 153 -31 187
rect -65 85 -31 119
rect -65 17 -31 51
rect -65 -51 -31 -17
rect -65 -119 -31 -85
rect -65 -187 -31 -153
rect -65 -255 -31 -221
rect -65 -323 -31 -289
rect -65 -391 -31 -357
rect -65 -459 -31 -425
rect 31 425 65 459
rect 31 357 65 391
rect 31 289 65 323
rect 31 221 65 255
rect 31 153 65 187
rect 31 85 65 119
rect 31 17 65 51
rect 31 -51 65 -17
rect 31 -119 65 -85
rect 31 -187 65 -153
rect 31 -255 65 -221
rect 31 -323 65 -289
rect 31 -391 65 -357
rect 31 -459 65 -425
rect 127 425 161 459
rect 127 357 161 391
rect 127 289 161 323
rect 127 221 161 255
rect 127 153 161 187
rect 127 85 161 119
rect 127 17 161 51
rect 127 -51 161 -17
rect 127 -119 161 -85
rect 127 -187 161 -153
rect 127 -255 161 -221
rect 127 -323 161 -289
rect 127 -391 161 -357
rect 127 -459 161 -425
rect 223 425 257 459
rect 223 357 257 391
rect 223 289 257 323
rect 223 221 257 255
rect 223 153 257 187
rect 223 85 257 119
rect 223 17 257 51
rect 223 -51 257 -17
rect 223 -119 257 -85
rect 223 -187 257 -153
rect 223 -255 257 -221
rect 223 -323 257 -289
rect 223 -391 257 -357
rect 223 -459 257 -425
rect 319 425 353 459
rect 319 357 353 391
rect 319 289 353 323
rect 319 221 353 255
rect 319 153 353 187
rect 319 85 353 119
rect 319 17 353 51
rect 319 -51 353 -17
rect 319 -119 353 -85
rect 319 -187 353 -153
rect 319 -255 353 -221
rect 319 -323 353 -289
rect 319 -391 353 -357
rect 319 -459 353 -425
rect 415 425 449 459
rect 415 357 449 391
rect 415 289 449 323
rect 415 221 449 255
rect 415 153 449 187
rect 415 85 449 119
rect 415 17 449 51
rect 415 -51 449 -17
rect 415 -119 449 -85
rect 415 -187 449 -153
rect 415 -255 449 -221
rect 415 -323 449 -289
rect 415 -391 449 -357
rect 415 -459 449 -425
<< psubdiff >>
rect -563 640 -459 674
rect -425 640 -391 674
rect -357 640 -323 674
rect -289 640 -255 674
rect -221 640 -187 674
rect -153 640 -119 674
rect -85 640 -51 674
rect -17 640 17 674
rect 51 640 85 674
rect 119 640 153 674
rect 187 640 221 674
rect 255 640 289 674
rect 323 640 357 674
rect 391 640 425 674
rect 459 640 563 674
rect -563 561 -529 640
rect -563 493 -529 527
rect 529 561 563 640
rect -563 425 -529 459
rect -563 357 -529 391
rect -563 289 -529 323
rect -563 221 -529 255
rect -563 153 -529 187
rect -563 85 -529 119
rect -563 17 -529 51
rect -563 -51 -529 -17
rect -563 -119 -529 -85
rect -563 -187 -529 -153
rect -563 -255 -529 -221
rect -563 -323 -529 -289
rect -563 -391 -529 -357
rect -563 -459 -529 -425
rect -563 -527 -529 -493
rect 529 493 563 527
rect 529 425 563 459
rect 529 357 563 391
rect 529 289 563 323
rect 529 221 563 255
rect 529 153 563 187
rect 529 85 563 119
rect 529 17 563 51
rect 529 -51 563 -17
rect 529 -119 563 -85
rect 529 -187 563 -153
rect 529 -255 563 -221
rect 529 -323 563 -289
rect 529 -391 563 -357
rect 529 -459 563 -425
rect -563 -640 -529 -561
rect 529 -527 563 -493
rect 529 -640 563 -561
rect -563 -674 -459 -640
rect -425 -674 -391 -640
rect -357 -674 -323 -640
rect -289 -674 -255 -640
rect -221 -674 -187 -640
rect -153 -674 -119 -640
rect -85 -674 -51 -640
rect -17 -674 17 -640
rect 51 -674 85 -640
rect 119 -674 153 -640
rect 187 -674 221 -640
rect 255 -674 289 -640
rect 323 -674 357 -640
rect 391 -674 425 -640
rect 459 -674 563 -640
<< psubdiffcont >>
rect -459 640 -425 674
rect -391 640 -357 674
rect -323 640 -289 674
rect -255 640 -221 674
rect -187 640 -153 674
rect -119 640 -85 674
rect -51 640 -17 674
rect 17 640 51 674
rect 85 640 119 674
rect 153 640 187 674
rect 221 640 255 674
rect 289 640 323 674
rect 357 640 391 674
rect 425 640 459 674
rect -563 527 -529 561
rect 529 527 563 561
rect -563 459 -529 493
rect -563 391 -529 425
rect -563 323 -529 357
rect -563 255 -529 289
rect -563 187 -529 221
rect -563 119 -529 153
rect -563 51 -529 85
rect -563 -17 -529 17
rect -563 -85 -529 -51
rect -563 -153 -529 -119
rect -563 -221 -529 -187
rect -563 -289 -529 -255
rect -563 -357 -529 -323
rect -563 -425 -529 -391
rect -563 -493 -529 -459
rect 529 459 563 493
rect 529 391 563 425
rect 529 323 563 357
rect 529 255 563 289
rect 529 187 563 221
rect 529 119 563 153
rect 529 51 563 85
rect 529 -17 563 17
rect 529 -85 563 -51
rect 529 -153 563 -119
rect 529 -221 563 -187
rect 529 -289 563 -255
rect 529 -357 563 -323
rect 529 -425 563 -391
rect 529 -493 563 -459
rect -563 -561 -529 -527
rect 529 -561 563 -527
rect -459 -674 -425 -640
rect -391 -674 -357 -640
rect -323 -674 -289 -640
rect -255 -674 -221 -640
rect -187 -674 -153 -640
rect -119 -674 -85 -640
rect -51 -674 -17 -640
rect 17 -674 51 -640
rect 85 -674 119 -640
rect 153 -674 187 -640
rect 221 -674 255 -640
rect 289 -674 323 -640
rect 357 -674 391 -640
rect 425 -674 459 -640
<< poly >>
rect -321 572 -255 588
rect -321 538 -305 572
rect -271 538 -255 572
rect -399 500 -369 526
rect -321 522 -255 538
rect -129 572 -63 588
rect -129 538 -113 572
rect -79 538 -63 572
rect -303 500 -273 522
rect -207 500 -177 526
rect -129 522 -63 538
rect 63 572 129 588
rect 63 538 79 572
rect 113 538 129 572
rect -111 500 -81 522
rect -15 500 15 526
rect 63 522 129 538
rect 255 572 321 588
rect 255 538 271 572
rect 305 538 321 572
rect 81 500 111 522
rect 177 500 207 526
rect 255 522 321 538
rect 273 500 303 522
rect 369 500 399 526
rect -399 -522 -369 -500
rect -417 -538 -351 -522
rect -303 -526 -273 -500
rect -207 -522 -177 -500
rect -417 -572 -401 -538
rect -367 -572 -351 -538
rect -417 -588 -351 -572
rect -225 -538 -159 -522
rect -111 -526 -81 -500
rect -15 -522 15 -500
rect -225 -572 -209 -538
rect -175 -572 -159 -538
rect -225 -588 -159 -572
rect -33 -538 33 -522
rect 81 -526 111 -500
rect 177 -522 207 -500
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect -33 -588 33 -572
rect 159 -538 225 -522
rect 273 -526 303 -500
rect 369 -522 399 -500
rect 159 -572 175 -538
rect 209 -572 225 -538
rect 159 -588 225 -572
rect 351 -538 417 -522
rect 351 -572 367 -538
rect 401 -572 417 -538
rect 351 -588 417 -572
<< polycont >>
rect -305 538 -271 572
rect -113 538 -79 572
rect 79 538 113 572
rect 271 538 305 572
rect -401 -572 -367 -538
rect -209 -572 -175 -538
rect -17 -572 17 -538
rect 175 -572 209 -538
rect 367 -572 401 -538
<< locali >>
rect -563 640 -459 674
rect -425 640 -391 674
rect -357 640 -323 674
rect -289 640 -255 674
rect -221 640 -187 674
rect -153 640 -119 674
rect -85 640 -51 674
rect -17 640 17 674
rect 51 640 85 674
rect 119 640 153 674
rect 187 640 221 674
rect 255 640 289 674
rect 323 640 357 674
rect 391 640 425 674
rect 459 640 563 674
rect -563 561 -529 640
rect -321 538 -305 572
rect -271 538 -255 572
rect -129 538 -113 572
rect -79 538 -63 572
rect 63 538 79 572
rect 113 538 129 572
rect 255 538 271 572
rect 305 538 321 572
rect 529 561 563 640
rect -563 493 -529 527
rect -563 425 -529 459
rect -563 357 -529 391
rect -563 289 -529 323
rect -563 221 -529 255
rect -563 153 -529 187
rect -563 85 -529 119
rect -563 17 -529 51
rect -563 -51 -529 -17
rect -563 -119 -529 -85
rect -563 -187 -529 -153
rect -563 -255 -529 -221
rect -563 -323 -529 -289
rect -563 -391 -529 -357
rect -563 -459 -529 -425
rect -563 -527 -529 -493
rect -449 485 -415 504
rect -449 413 -415 425
rect -449 341 -415 357
rect -449 269 -415 289
rect -449 197 -415 221
rect -449 125 -415 153
rect -449 53 -415 85
rect -449 -17 -415 17
rect -449 -85 -415 -53
rect -449 -153 -415 -125
rect -449 -221 -415 -197
rect -449 -289 -415 -269
rect -449 -357 -415 -341
rect -449 -425 -415 -413
rect -449 -504 -415 -485
rect -353 485 -319 504
rect -353 413 -319 425
rect -353 341 -319 357
rect -353 269 -319 289
rect -353 197 -319 221
rect -353 125 -319 153
rect -353 53 -319 85
rect -353 -17 -319 17
rect -353 -85 -319 -53
rect -353 -153 -319 -125
rect -353 -221 -319 -197
rect -353 -289 -319 -269
rect -353 -357 -319 -341
rect -353 -425 -319 -413
rect -353 -504 -319 -485
rect -257 485 -223 504
rect -257 413 -223 425
rect -257 341 -223 357
rect -257 269 -223 289
rect -257 197 -223 221
rect -257 125 -223 153
rect -257 53 -223 85
rect -257 -17 -223 17
rect -257 -85 -223 -53
rect -257 -153 -223 -125
rect -257 -221 -223 -197
rect -257 -289 -223 -269
rect -257 -357 -223 -341
rect -257 -425 -223 -413
rect -257 -504 -223 -485
rect -161 485 -127 504
rect -161 413 -127 425
rect -161 341 -127 357
rect -161 269 -127 289
rect -161 197 -127 221
rect -161 125 -127 153
rect -161 53 -127 85
rect -161 -17 -127 17
rect -161 -85 -127 -53
rect -161 -153 -127 -125
rect -161 -221 -127 -197
rect -161 -289 -127 -269
rect -161 -357 -127 -341
rect -161 -425 -127 -413
rect -161 -504 -127 -485
rect -65 485 -31 504
rect -65 413 -31 425
rect -65 341 -31 357
rect -65 269 -31 289
rect -65 197 -31 221
rect -65 125 -31 153
rect -65 53 -31 85
rect -65 -17 -31 17
rect -65 -85 -31 -53
rect -65 -153 -31 -125
rect -65 -221 -31 -197
rect -65 -289 -31 -269
rect -65 -357 -31 -341
rect -65 -425 -31 -413
rect -65 -504 -31 -485
rect 31 485 65 504
rect 31 413 65 425
rect 31 341 65 357
rect 31 269 65 289
rect 31 197 65 221
rect 31 125 65 153
rect 31 53 65 85
rect 31 -17 65 17
rect 31 -85 65 -53
rect 31 -153 65 -125
rect 31 -221 65 -197
rect 31 -289 65 -269
rect 31 -357 65 -341
rect 31 -425 65 -413
rect 31 -504 65 -485
rect 127 485 161 504
rect 127 413 161 425
rect 127 341 161 357
rect 127 269 161 289
rect 127 197 161 221
rect 127 125 161 153
rect 127 53 161 85
rect 127 -17 161 17
rect 127 -85 161 -53
rect 127 -153 161 -125
rect 127 -221 161 -197
rect 127 -289 161 -269
rect 127 -357 161 -341
rect 127 -425 161 -413
rect 127 -504 161 -485
rect 223 485 257 504
rect 223 413 257 425
rect 223 341 257 357
rect 223 269 257 289
rect 223 197 257 221
rect 223 125 257 153
rect 223 53 257 85
rect 223 -17 257 17
rect 223 -85 257 -53
rect 223 -153 257 -125
rect 223 -221 257 -197
rect 223 -289 257 -269
rect 223 -357 257 -341
rect 223 -425 257 -413
rect 223 -504 257 -485
rect 319 485 353 504
rect 319 413 353 425
rect 319 341 353 357
rect 319 269 353 289
rect 319 197 353 221
rect 319 125 353 153
rect 319 53 353 85
rect 319 -17 353 17
rect 319 -85 353 -53
rect 319 -153 353 -125
rect 319 -221 353 -197
rect 319 -289 353 -269
rect 319 -357 353 -341
rect 319 -425 353 -413
rect 319 -504 353 -485
rect 415 485 449 504
rect 415 413 449 425
rect 415 341 449 357
rect 415 269 449 289
rect 415 197 449 221
rect 415 125 449 153
rect 415 53 449 85
rect 415 -17 449 17
rect 415 -85 449 -53
rect 415 -153 449 -125
rect 415 -221 449 -197
rect 415 -289 449 -269
rect 415 -357 449 -341
rect 415 -425 449 -413
rect 415 -504 449 -485
rect 529 493 563 527
rect 529 425 563 459
rect 529 357 563 391
rect 529 289 563 323
rect 529 221 563 255
rect 529 153 563 187
rect 529 85 563 119
rect 529 17 563 51
rect 529 -51 563 -17
rect 529 -119 563 -85
rect 529 -187 563 -153
rect 529 -255 563 -221
rect 529 -323 563 -289
rect 529 -391 563 -357
rect 529 -459 563 -425
rect 529 -527 563 -493
rect -563 -640 -529 -561
rect -417 -572 -401 -538
rect -367 -572 -351 -538
rect -225 -572 -209 -538
rect -175 -572 -159 -538
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect 159 -572 175 -538
rect 209 -572 225 -538
rect 351 -572 367 -538
rect 401 -572 417 -538
rect 529 -640 563 -561
rect -563 -674 -459 -640
rect -425 -674 -391 -640
rect -357 -674 -323 -640
rect -289 -674 -255 -640
rect -221 -674 -187 -640
rect -153 -674 -119 -640
rect -85 -674 -51 -640
rect -17 -674 17 -640
rect 51 -674 85 -640
rect 119 -674 153 -640
rect 187 -674 221 -640
rect 255 -674 289 -640
rect 323 -674 357 -640
rect 391 -674 425 -640
rect 459 -674 563 -640
<< viali >>
rect -305 538 -271 572
rect -113 538 -79 572
rect 79 538 113 572
rect 271 538 305 572
rect -449 459 -415 485
rect -449 451 -415 459
rect -449 391 -415 413
rect -449 379 -415 391
rect -449 323 -415 341
rect -449 307 -415 323
rect -449 255 -415 269
rect -449 235 -415 255
rect -449 187 -415 197
rect -449 163 -415 187
rect -449 119 -415 125
rect -449 91 -415 119
rect -449 51 -415 53
rect -449 19 -415 51
rect -449 -51 -415 -19
rect -449 -53 -415 -51
rect -449 -119 -415 -91
rect -449 -125 -415 -119
rect -449 -187 -415 -163
rect -449 -197 -415 -187
rect -449 -255 -415 -235
rect -449 -269 -415 -255
rect -449 -323 -415 -307
rect -449 -341 -415 -323
rect -449 -391 -415 -379
rect -449 -413 -415 -391
rect -449 -459 -415 -451
rect -449 -485 -415 -459
rect -353 459 -319 485
rect -353 451 -319 459
rect -353 391 -319 413
rect -353 379 -319 391
rect -353 323 -319 341
rect -353 307 -319 323
rect -353 255 -319 269
rect -353 235 -319 255
rect -353 187 -319 197
rect -353 163 -319 187
rect -353 119 -319 125
rect -353 91 -319 119
rect -353 51 -319 53
rect -353 19 -319 51
rect -353 -51 -319 -19
rect -353 -53 -319 -51
rect -353 -119 -319 -91
rect -353 -125 -319 -119
rect -353 -187 -319 -163
rect -353 -197 -319 -187
rect -353 -255 -319 -235
rect -353 -269 -319 -255
rect -353 -323 -319 -307
rect -353 -341 -319 -323
rect -353 -391 -319 -379
rect -353 -413 -319 -391
rect -353 -459 -319 -451
rect -353 -485 -319 -459
rect -257 459 -223 485
rect -257 451 -223 459
rect -257 391 -223 413
rect -257 379 -223 391
rect -257 323 -223 341
rect -257 307 -223 323
rect -257 255 -223 269
rect -257 235 -223 255
rect -257 187 -223 197
rect -257 163 -223 187
rect -257 119 -223 125
rect -257 91 -223 119
rect -257 51 -223 53
rect -257 19 -223 51
rect -257 -51 -223 -19
rect -257 -53 -223 -51
rect -257 -119 -223 -91
rect -257 -125 -223 -119
rect -257 -187 -223 -163
rect -257 -197 -223 -187
rect -257 -255 -223 -235
rect -257 -269 -223 -255
rect -257 -323 -223 -307
rect -257 -341 -223 -323
rect -257 -391 -223 -379
rect -257 -413 -223 -391
rect -257 -459 -223 -451
rect -257 -485 -223 -459
rect -161 459 -127 485
rect -161 451 -127 459
rect -161 391 -127 413
rect -161 379 -127 391
rect -161 323 -127 341
rect -161 307 -127 323
rect -161 255 -127 269
rect -161 235 -127 255
rect -161 187 -127 197
rect -161 163 -127 187
rect -161 119 -127 125
rect -161 91 -127 119
rect -161 51 -127 53
rect -161 19 -127 51
rect -161 -51 -127 -19
rect -161 -53 -127 -51
rect -161 -119 -127 -91
rect -161 -125 -127 -119
rect -161 -187 -127 -163
rect -161 -197 -127 -187
rect -161 -255 -127 -235
rect -161 -269 -127 -255
rect -161 -323 -127 -307
rect -161 -341 -127 -323
rect -161 -391 -127 -379
rect -161 -413 -127 -391
rect -161 -459 -127 -451
rect -161 -485 -127 -459
rect -65 459 -31 485
rect -65 451 -31 459
rect -65 391 -31 413
rect -65 379 -31 391
rect -65 323 -31 341
rect -65 307 -31 323
rect -65 255 -31 269
rect -65 235 -31 255
rect -65 187 -31 197
rect -65 163 -31 187
rect -65 119 -31 125
rect -65 91 -31 119
rect -65 51 -31 53
rect -65 19 -31 51
rect -65 -51 -31 -19
rect -65 -53 -31 -51
rect -65 -119 -31 -91
rect -65 -125 -31 -119
rect -65 -187 -31 -163
rect -65 -197 -31 -187
rect -65 -255 -31 -235
rect -65 -269 -31 -255
rect -65 -323 -31 -307
rect -65 -341 -31 -323
rect -65 -391 -31 -379
rect -65 -413 -31 -391
rect -65 -459 -31 -451
rect -65 -485 -31 -459
rect 31 459 65 485
rect 31 451 65 459
rect 31 391 65 413
rect 31 379 65 391
rect 31 323 65 341
rect 31 307 65 323
rect 31 255 65 269
rect 31 235 65 255
rect 31 187 65 197
rect 31 163 65 187
rect 31 119 65 125
rect 31 91 65 119
rect 31 51 65 53
rect 31 19 65 51
rect 31 -51 65 -19
rect 31 -53 65 -51
rect 31 -119 65 -91
rect 31 -125 65 -119
rect 31 -187 65 -163
rect 31 -197 65 -187
rect 31 -255 65 -235
rect 31 -269 65 -255
rect 31 -323 65 -307
rect 31 -341 65 -323
rect 31 -391 65 -379
rect 31 -413 65 -391
rect 31 -459 65 -451
rect 31 -485 65 -459
rect 127 459 161 485
rect 127 451 161 459
rect 127 391 161 413
rect 127 379 161 391
rect 127 323 161 341
rect 127 307 161 323
rect 127 255 161 269
rect 127 235 161 255
rect 127 187 161 197
rect 127 163 161 187
rect 127 119 161 125
rect 127 91 161 119
rect 127 51 161 53
rect 127 19 161 51
rect 127 -51 161 -19
rect 127 -53 161 -51
rect 127 -119 161 -91
rect 127 -125 161 -119
rect 127 -187 161 -163
rect 127 -197 161 -187
rect 127 -255 161 -235
rect 127 -269 161 -255
rect 127 -323 161 -307
rect 127 -341 161 -323
rect 127 -391 161 -379
rect 127 -413 161 -391
rect 127 -459 161 -451
rect 127 -485 161 -459
rect 223 459 257 485
rect 223 451 257 459
rect 223 391 257 413
rect 223 379 257 391
rect 223 323 257 341
rect 223 307 257 323
rect 223 255 257 269
rect 223 235 257 255
rect 223 187 257 197
rect 223 163 257 187
rect 223 119 257 125
rect 223 91 257 119
rect 223 51 257 53
rect 223 19 257 51
rect 223 -51 257 -19
rect 223 -53 257 -51
rect 223 -119 257 -91
rect 223 -125 257 -119
rect 223 -187 257 -163
rect 223 -197 257 -187
rect 223 -255 257 -235
rect 223 -269 257 -255
rect 223 -323 257 -307
rect 223 -341 257 -323
rect 223 -391 257 -379
rect 223 -413 257 -391
rect 223 -459 257 -451
rect 223 -485 257 -459
rect 319 459 353 485
rect 319 451 353 459
rect 319 391 353 413
rect 319 379 353 391
rect 319 323 353 341
rect 319 307 353 323
rect 319 255 353 269
rect 319 235 353 255
rect 319 187 353 197
rect 319 163 353 187
rect 319 119 353 125
rect 319 91 353 119
rect 319 51 353 53
rect 319 19 353 51
rect 319 -51 353 -19
rect 319 -53 353 -51
rect 319 -119 353 -91
rect 319 -125 353 -119
rect 319 -187 353 -163
rect 319 -197 353 -187
rect 319 -255 353 -235
rect 319 -269 353 -255
rect 319 -323 353 -307
rect 319 -341 353 -323
rect 319 -391 353 -379
rect 319 -413 353 -391
rect 319 -459 353 -451
rect 319 -485 353 -459
rect 415 459 449 485
rect 415 451 449 459
rect 415 391 449 413
rect 415 379 449 391
rect 415 323 449 341
rect 415 307 449 323
rect 415 255 449 269
rect 415 235 449 255
rect 415 187 449 197
rect 415 163 449 187
rect 415 119 449 125
rect 415 91 449 119
rect 415 51 449 53
rect 415 19 449 51
rect 415 -51 449 -19
rect 415 -53 449 -51
rect 415 -119 449 -91
rect 415 -125 449 -119
rect 415 -187 449 -163
rect 415 -197 449 -187
rect 415 -255 449 -235
rect 415 -269 449 -255
rect 415 -323 449 -307
rect 415 -341 449 -323
rect 415 -391 449 -379
rect 415 -413 449 -391
rect 415 -459 449 -451
rect 415 -485 449 -459
rect -401 -572 -367 -538
rect -209 -572 -175 -538
rect -17 -572 17 -538
rect 175 -572 209 -538
rect 367 -572 401 -538
<< metal1 >>
rect -317 572 -259 578
rect -317 538 -305 572
rect -271 538 -259 572
rect -317 532 -259 538
rect -125 572 -67 578
rect -125 538 -113 572
rect -79 538 -67 572
rect -125 532 -67 538
rect 67 572 125 578
rect 67 538 79 572
rect 113 538 125 572
rect 67 532 125 538
rect 259 572 317 578
rect 259 538 271 572
rect 305 538 317 572
rect 259 532 317 538
rect -455 485 -409 500
rect -455 451 -449 485
rect -415 451 -409 485
rect -455 413 -409 451
rect -455 379 -449 413
rect -415 379 -409 413
rect -455 341 -409 379
rect -455 307 -449 341
rect -415 307 -409 341
rect -455 269 -409 307
rect -455 235 -449 269
rect -415 235 -409 269
rect -455 197 -409 235
rect -455 163 -449 197
rect -415 163 -409 197
rect -455 125 -409 163
rect -455 91 -449 125
rect -415 91 -409 125
rect -455 53 -409 91
rect -455 19 -449 53
rect -415 19 -409 53
rect -455 -19 -409 19
rect -455 -53 -449 -19
rect -415 -53 -409 -19
rect -455 -91 -409 -53
rect -455 -125 -449 -91
rect -415 -125 -409 -91
rect -455 -163 -409 -125
rect -455 -197 -449 -163
rect -415 -197 -409 -163
rect -455 -235 -409 -197
rect -455 -269 -449 -235
rect -415 -269 -409 -235
rect -455 -307 -409 -269
rect -455 -341 -449 -307
rect -415 -341 -409 -307
rect -455 -379 -409 -341
rect -455 -413 -449 -379
rect -415 -413 -409 -379
rect -455 -451 -409 -413
rect -455 -485 -449 -451
rect -415 -485 -409 -451
rect -455 -500 -409 -485
rect -359 485 -313 500
rect -359 451 -353 485
rect -319 451 -313 485
rect -359 413 -313 451
rect -359 379 -353 413
rect -319 379 -313 413
rect -359 341 -313 379
rect -359 307 -353 341
rect -319 307 -313 341
rect -359 269 -313 307
rect -359 235 -353 269
rect -319 235 -313 269
rect -359 197 -313 235
rect -359 163 -353 197
rect -319 163 -313 197
rect -359 125 -313 163
rect -359 91 -353 125
rect -319 91 -313 125
rect -359 53 -313 91
rect -359 19 -353 53
rect -319 19 -313 53
rect -359 -19 -313 19
rect -359 -53 -353 -19
rect -319 -53 -313 -19
rect -359 -91 -313 -53
rect -359 -125 -353 -91
rect -319 -125 -313 -91
rect -359 -163 -313 -125
rect -359 -197 -353 -163
rect -319 -197 -313 -163
rect -359 -235 -313 -197
rect -359 -269 -353 -235
rect -319 -269 -313 -235
rect -359 -307 -313 -269
rect -359 -341 -353 -307
rect -319 -341 -313 -307
rect -359 -379 -313 -341
rect -359 -413 -353 -379
rect -319 -413 -313 -379
rect -359 -451 -313 -413
rect -359 -485 -353 -451
rect -319 -485 -313 -451
rect -359 -500 -313 -485
rect -263 485 -217 500
rect -263 451 -257 485
rect -223 451 -217 485
rect -263 413 -217 451
rect -263 379 -257 413
rect -223 379 -217 413
rect -263 341 -217 379
rect -263 307 -257 341
rect -223 307 -217 341
rect -263 269 -217 307
rect -263 235 -257 269
rect -223 235 -217 269
rect -263 197 -217 235
rect -263 163 -257 197
rect -223 163 -217 197
rect -263 125 -217 163
rect -263 91 -257 125
rect -223 91 -217 125
rect -263 53 -217 91
rect -263 19 -257 53
rect -223 19 -217 53
rect -263 -19 -217 19
rect -263 -53 -257 -19
rect -223 -53 -217 -19
rect -263 -91 -217 -53
rect -263 -125 -257 -91
rect -223 -125 -217 -91
rect -263 -163 -217 -125
rect -263 -197 -257 -163
rect -223 -197 -217 -163
rect -263 -235 -217 -197
rect -263 -269 -257 -235
rect -223 -269 -217 -235
rect -263 -307 -217 -269
rect -263 -341 -257 -307
rect -223 -341 -217 -307
rect -263 -379 -217 -341
rect -263 -413 -257 -379
rect -223 -413 -217 -379
rect -263 -451 -217 -413
rect -263 -485 -257 -451
rect -223 -485 -217 -451
rect -263 -500 -217 -485
rect -167 485 -121 500
rect -167 451 -161 485
rect -127 451 -121 485
rect -167 413 -121 451
rect -167 379 -161 413
rect -127 379 -121 413
rect -167 341 -121 379
rect -167 307 -161 341
rect -127 307 -121 341
rect -167 269 -121 307
rect -167 235 -161 269
rect -127 235 -121 269
rect -167 197 -121 235
rect -167 163 -161 197
rect -127 163 -121 197
rect -167 125 -121 163
rect -167 91 -161 125
rect -127 91 -121 125
rect -167 53 -121 91
rect -167 19 -161 53
rect -127 19 -121 53
rect -167 -19 -121 19
rect -167 -53 -161 -19
rect -127 -53 -121 -19
rect -167 -91 -121 -53
rect -167 -125 -161 -91
rect -127 -125 -121 -91
rect -167 -163 -121 -125
rect -167 -197 -161 -163
rect -127 -197 -121 -163
rect -167 -235 -121 -197
rect -167 -269 -161 -235
rect -127 -269 -121 -235
rect -167 -307 -121 -269
rect -167 -341 -161 -307
rect -127 -341 -121 -307
rect -167 -379 -121 -341
rect -167 -413 -161 -379
rect -127 -413 -121 -379
rect -167 -451 -121 -413
rect -167 -485 -161 -451
rect -127 -485 -121 -451
rect -167 -500 -121 -485
rect -71 485 -25 500
rect -71 451 -65 485
rect -31 451 -25 485
rect -71 413 -25 451
rect -71 379 -65 413
rect -31 379 -25 413
rect -71 341 -25 379
rect -71 307 -65 341
rect -31 307 -25 341
rect -71 269 -25 307
rect -71 235 -65 269
rect -31 235 -25 269
rect -71 197 -25 235
rect -71 163 -65 197
rect -31 163 -25 197
rect -71 125 -25 163
rect -71 91 -65 125
rect -31 91 -25 125
rect -71 53 -25 91
rect -71 19 -65 53
rect -31 19 -25 53
rect -71 -19 -25 19
rect -71 -53 -65 -19
rect -31 -53 -25 -19
rect -71 -91 -25 -53
rect -71 -125 -65 -91
rect -31 -125 -25 -91
rect -71 -163 -25 -125
rect -71 -197 -65 -163
rect -31 -197 -25 -163
rect -71 -235 -25 -197
rect -71 -269 -65 -235
rect -31 -269 -25 -235
rect -71 -307 -25 -269
rect -71 -341 -65 -307
rect -31 -341 -25 -307
rect -71 -379 -25 -341
rect -71 -413 -65 -379
rect -31 -413 -25 -379
rect -71 -451 -25 -413
rect -71 -485 -65 -451
rect -31 -485 -25 -451
rect -71 -500 -25 -485
rect 25 485 71 500
rect 25 451 31 485
rect 65 451 71 485
rect 25 413 71 451
rect 25 379 31 413
rect 65 379 71 413
rect 25 341 71 379
rect 25 307 31 341
rect 65 307 71 341
rect 25 269 71 307
rect 25 235 31 269
rect 65 235 71 269
rect 25 197 71 235
rect 25 163 31 197
rect 65 163 71 197
rect 25 125 71 163
rect 25 91 31 125
rect 65 91 71 125
rect 25 53 71 91
rect 25 19 31 53
rect 65 19 71 53
rect 25 -19 71 19
rect 25 -53 31 -19
rect 65 -53 71 -19
rect 25 -91 71 -53
rect 25 -125 31 -91
rect 65 -125 71 -91
rect 25 -163 71 -125
rect 25 -197 31 -163
rect 65 -197 71 -163
rect 25 -235 71 -197
rect 25 -269 31 -235
rect 65 -269 71 -235
rect 25 -307 71 -269
rect 25 -341 31 -307
rect 65 -341 71 -307
rect 25 -379 71 -341
rect 25 -413 31 -379
rect 65 -413 71 -379
rect 25 -451 71 -413
rect 25 -485 31 -451
rect 65 -485 71 -451
rect 25 -500 71 -485
rect 121 485 167 500
rect 121 451 127 485
rect 161 451 167 485
rect 121 413 167 451
rect 121 379 127 413
rect 161 379 167 413
rect 121 341 167 379
rect 121 307 127 341
rect 161 307 167 341
rect 121 269 167 307
rect 121 235 127 269
rect 161 235 167 269
rect 121 197 167 235
rect 121 163 127 197
rect 161 163 167 197
rect 121 125 167 163
rect 121 91 127 125
rect 161 91 167 125
rect 121 53 167 91
rect 121 19 127 53
rect 161 19 167 53
rect 121 -19 167 19
rect 121 -53 127 -19
rect 161 -53 167 -19
rect 121 -91 167 -53
rect 121 -125 127 -91
rect 161 -125 167 -91
rect 121 -163 167 -125
rect 121 -197 127 -163
rect 161 -197 167 -163
rect 121 -235 167 -197
rect 121 -269 127 -235
rect 161 -269 167 -235
rect 121 -307 167 -269
rect 121 -341 127 -307
rect 161 -341 167 -307
rect 121 -379 167 -341
rect 121 -413 127 -379
rect 161 -413 167 -379
rect 121 -451 167 -413
rect 121 -485 127 -451
rect 161 -485 167 -451
rect 121 -500 167 -485
rect 217 485 263 500
rect 217 451 223 485
rect 257 451 263 485
rect 217 413 263 451
rect 217 379 223 413
rect 257 379 263 413
rect 217 341 263 379
rect 217 307 223 341
rect 257 307 263 341
rect 217 269 263 307
rect 217 235 223 269
rect 257 235 263 269
rect 217 197 263 235
rect 217 163 223 197
rect 257 163 263 197
rect 217 125 263 163
rect 217 91 223 125
rect 257 91 263 125
rect 217 53 263 91
rect 217 19 223 53
rect 257 19 263 53
rect 217 -19 263 19
rect 217 -53 223 -19
rect 257 -53 263 -19
rect 217 -91 263 -53
rect 217 -125 223 -91
rect 257 -125 263 -91
rect 217 -163 263 -125
rect 217 -197 223 -163
rect 257 -197 263 -163
rect 217 -235 263 -197
rect 217 -269 223 -235
rect 257 -269 263 -235
rect 217 -307 263 -269
rect 217 -341 223 -307
rect 257 -341 263 -307
rect 217 -379 263 -341
rect 217 -413 223 -379
rect 257 -413 263 -379
rect 217 -451 263 -413
rect 217 -485 223 -451
rect 257 -485 263 -451
rect 217 -500 263 -485
rect 313 485 359 500
rect 313 451 319 485
rect 353 451 359 485
rect 313 413 359 451
rect 313 379 319 413
rect 353 379 359 413
rect 313 341 359 379
rect 313 307 319 341
rect 353 307 359 341
rect 313 269 359 307
rect 313 235 319 269
rect 353 235 359 269
rect 313 197 359 235
rect 313 163 319 197
rect 353 163 359 197
rect 313 125 359 163
rect 313 91 319 125
rect 353 91 359 125
rect 313 53 359 91
rect 313 19 319 53
rect 353 19 359 53
rect 313 -19 359 19
rect 313 -53 319 -19
rect 353 -53 359 -19
rect 313 -91 359 -53
rect 313 -125 319 -91
rect 353 -125 359 -91
rect 313 -163 359 -125
rect 313 -197 319 -163
rect 353 -197 359 -163
rect 313 -235 359 -197
rect 313 -269 319 -235
rect 353 -269 359 -235
rect 313 -307 359 -269
rect 313 -341 319 -307
rect 353 -341 359 -307
rect 313 -379 359 -341
rect 313 -413 319 -379
rect 353 -413 359 -379
rect 313 -451 359 -413
rect 313 -485 319 -451
rect 353 -485 359 -451
rect 313 -500 359 -485
rect 409 485 455 500
rect 409 451 415 485
rect 449 451 455 485
rect 409 413 455 451
rect 409 379 415 413
rect 449 379 455 413
rect 409 341 455 379
rect 409 307 415 341
rect 449 307 455 341
rect 409 269 455 307
rect 409 235 415 269
rect 449 235 455 269
rect 409 197 455 235
rect 409 163 415 197
rect 449 163 455 197
rect 409 125 455 163
rect 409 91 415 125
rect 449 91 455 125
rect 409 53 455 91
rect 409 19 415 53
rect 449 19 455 53
rect 409 -19 455 19
rect 409 -53 415 -19
rect 449 -53 455 -19
rect 409 -91 455 -53
rect 409 -125 415 -91
rect 449 -125 455 -91
rect 409 -163 455 -125
rect 409 -197 415 -163
rect 449 -197 455 -163
rect 409 -235 455 -197
rect 409 -269 415 -235
rect 449 -269 455 -235
rect 409 -307 455 -269
rect 409 -341 415 -307
rect 449 -341 455 -307
rect 409 -379 455 -341
rect 409 -413 415 -379
rect 449 -413 455 -379
rect 409 -451 455 -413
rect 409 -485 415 -451
rect 449 -485 455 -451
rect 409 -500 455 -485
rect -413 -538 -355 -532
rect -413 -572 -401 -538
rect -367 -572 -355 -538
rect -413 -578 -355 -572
rect -221 -538 -163 -532
rect -221 -572 -209 -538
rect -175 -572 -163 -538
rect -221 -578 -163 -572
rect -29 -538 29 -532
rect -29 -572 -17 -538
rect 17 -572 29 -538
rect -29 -578 29 -572
rect 163 -538 221 -532
rect 163 -572 175 -538
rect 209 -572 221 -538
rect 163 -578 221 -572
rect 355 -538 413 -532
rect 355 -572 367 -538
rect 401 -572 413 -538
rect 355 -578 413 -572
<< properties >>
string FIXED_BBOX -546 -657 546 657
<< end >>
