magic
tech sky130A
magscale 1 2
timestamp 1635855079
<< error_p >>
rect -29 812 29 818
rect -29 778 -17 812
rect -29 772 29 778
rect -29 -778 29 -772
rect -29 -812 -17 -778
rect -29 -818 29 -812
<< pwell >>
rect -201 -940 201 940
<< nmoslvt >>
rect -15 -740 15 740
<< ndiff >>
rect -73 697 -15 740
rect -73 663 -61 697
rect -27 663 -15 697
rect -73 629 -15 663
rect -73 595 -61 629
rect -27 595 -15 629
rect -73 561 -15 595
rect -73 527 -61 561
rect -27 527 -15 561
rect -73 493 -15 527
rect -73 459 -61 493
rect -27 459 -15 493
rect -73 425 -15 459
rect -73 391 -61 425
rect -27 391 -15 425
rect -73 357 -15 391
rect -73 323 -61 357
rect -27 323 -15 357
rect -73 289 -15 323
rect -73 255 -61 289
rect -27 255 -15 289
rect -73 221 -15 255
rect -73 187 -61 221
rect -27 187 -15 221
rect -73 153 -15 187
rect -73 119 -61 153
rect -27 119 -15 153
rect -73 85 -15 119
rect -73 51 -61 85
rect -27 51 -15 85
rect -73 17 -15 51
rect -73 -17 -61 17
rect -27 -17 -15 17
rect -73 -51 -15 -17
rect -73 -85 -61 -51
rect -27 -85 -15 -51
rect -73 -119 -15 -85
rect -73 -153 -61 -119
rect -27 -153 -15 -119
rect -73 -187 -15 -153
rect -73 -221 -61 -187
rect -27 -221 -15 -187
rect -73 -255 -15 -221
rect -73 -289 -61 -255
rect -27 -289 -15 -255
rect -73 -323 -15 -289
rect -73 -357 -61 -323
rect -27 -357 -15 -323
rect -73 -391 -15 -357
rect -73 -425 -61 -391
rect -27 -425 -15 -391
rect -73 -459 -15 -425
rect -73 -493 -61 -459
rect -27 -493 -15 -459
rect -73 -527 -15 -493
rect -73 -561 -61 -527
rect -27 -561 -15 -527
rect -73 -595 -15 -561
rect -73 -629 -61 -595
rect -27 -629 -15 -595
rect -73 -663 -15 -629
rect -73 -697 -61 -663
rect -27 -697 -15 -663
rect -73 -740 -15 -697
rect 15 697 73 740
rect 15 663 27 697
rect 61 663 73 697
rect 15 629 73 663
rect 15 595 27 629
rect 61 595 73 629
rect 15 561 73 595
rect 15 527 27 561
rect 61 527 73 561
rect 15 493 73 527
rect 15 459 27 493
rect 61 459 73 493
rect 15 425 73 459
rect 15 391 27 425
rect 61 391 73 425
rect 15 357 73 391
rect 15 323 27 357
rect 61 323 73 357
rect 15 289 73 323
rect 15 255 27 289
rect 61 255 73 289
rect 15 221 73 255
rect 15 187 27 221
rect 61 187 73 221
rect 15 153 73 187
rect 15 119 27 153
rect 61 119 73 153
rect 15 85 73 119
rect 15 51 27 85
rect 61 51 73 85
rect 15 17 73 51
rect 15 -17 27 17
rect 61 -17 73 17
rect 15 -51 73 -17
rect 15 -85 27 -51
rect 61 -85 73 -51
rect 15 -119 73 -85
rect 15 -153 27 -119
rect 61 -153 73 -119
rect 15 -187 73 -153
rect 15 -221 27 -187
rect 61 -221 73 -187
rect 15 -255 73 -221
rect 15 -289 27 -255
rect 61 -289 73 -255
rect 15 -323 73 -289
rect 15 -357 27 -323
rect 61 -357 73 -323
rect 15 -391 73 -357
rect 15 -425 27 -391
rect 61 -425 73 -391
rect 15 -459 73 -425
rect 15 -493 27 -459
rect 61 -493 73 -459
rect 15 -527 73 -493
rect 15 -561 27 -527
rect 61 -561 73 -527
rect 15 -595 73 -561
rect 15 -629 27 -595
rect 61 -629 73 -595
rect 15 -663 73 -629
rect 15 -697 27 -663
rect 61 -697 73 -663
rect 15 -740 73 -697
<< ndiffc >>
rect -61 663 -27 697
rect -61 595 -27 629
rect -61 527 -27 561
rect -61 459 -27 493
rect -61 391 -27 425
rect -61 323 -27 357
rect -61 255 -27 289
rect -61 187 -27 221
rect -61 119 -27 153
rect -61 51 -27 85
rect -61 -17 -27 17
rect -61 -85 -27 -51
rect -61 -153 -27 -119
rect -61 -221 -27 -187
rect -61 -289 -27 -255
rect -61 -357 -27 -323
rect -61 -425 -27 -391
rect -61 -493 -27 -459
rect -61 -561 -27 -527
rect -61 -629 -27 -595
rect -61 -697 -27 -663
rect 27 663 61 697
rect 27 595 61 629
rect 27 527 61 561
rect 27 459 61 493
rect 27 391 61 425
rect 27 323 61 357
rect 27 255 61 289
rect 27 187 61 221
rect 27 119 61 153
rect 27 51 61 85
rect 27 -17 61 17
rect 27 -85 61 -51
rect 27 -153 61 -119
rect 27 -221 61 -187
rect 27 -289 61 -255
rect 27 -357 61 -323
rect 27 -425 61 -391
rect 27 -493 61 -459
rect 27 -561 61 -527
rect 27 -629 61 -595
rect 27 -697 61 -663
<< psubdiff >>
rect -175 880 -51 914
rect -17 880 17 914
rect 51 880 175 914
rect -175 799 -141 880
rect -175 731 -141 765
rect 141 799 175 880
rect -175 663 -141 697
rect -175 595 -141 629
rect -175 527 -141 561
rect -175 459 -141 493
rect -175 391 -141 425
rect -175 323 -141 357
rect -175 255 -141 289
rect -175 187 -141 221
rect -175 119 -141 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -175 -153 -141 -119
rect -175 -221 -141 -187
rect -175 -289 -141 -255
rect -175 -357 -141 -323
rect -175 -425 -141 -391
rect -175 -493 -141 -459
rect -175 -561 -141 -527
rect -175 -629 -141 -595
rect -175 -697 -141 -663
rect -175 -765 -141 -731
rect 141 731 175 765
rect 141 663 175 697
rect 141 595 175 629
rect 141 527 175 561
rect 141 459 175 493
rect 141 391 175 425
rect 141 323 175 357
rect 141 255 175 289
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
rect 141 -289 175 -255
rect 141 -357 175 -323
rect 141 -425 175 -391
rect 141 -493 175 -459
rect 141 -561 175 -527
rect 141 -629 175 -595
rect 141 -697 175 -663
rect -175 -880 -141 -799
rect 141 -765 175 -731
rect 141 -880 175 -799
rect -175 -914 -51 -880
rect -17 -914 17 -880
rect 51 -914 175 -880
<< psubdiffcont >>
rect -51 880 -17 914
rect 17 880 51 914
rect -175 765 -141 799
rect 141 765 175 799
rect -175 697 -141 731
rect -175 629 -141 663
rect -175 561 -141 595
rect -175 493 -141 527
rect -175 425 -141 459
rect -175 357 -141 391
rect -175 289 -141 323
rect -175 221 -141 255
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -175 -255 -141 -221
rect -175 -323 -141 -289
rect -175 -391 -141 -357
rect -175 -459 -141 -425
rect -175 -527 -141 -493
rect -175 -595 -141 -561
rect -175 -663 -141 -629
rect -175 -731 -141 -697
rect 141 697 175 731
rect 141 629 175 663
rect 141 561 175 595
rect 141 493 175 527
rect 141 425 175 459
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect 141 -459 175 -425
rect 141 -527 175 -493
rect 141 -595 175 -561
rect 141 -663 175 -629
rect 141 -731 175 -697
rect -175 -799 -141 -765
rect 141 -799 175 -765
rect -51 -914 -17 -880
rect 17 -914 51 -880
<< poly >>
rect -33 812 33 828
rect -33 778 -17 812
rect 17 778 33 812
rect -33 762 33 778
rect -15 740 15 762
rect -15 -762 15 -740
rect -33 -778 33 -762
rect -33 -812 -17 -778
rect 17 -812 33 -778
rect -33 -828 33 -812
<< polycont >>
rect -17 778 17 812
rect -17 -812 17 -778
<< locali >>
rect -175 880 -51 914
rect -17 880 17 914
rect 51 880 175 914
rect -175 799 -141 880
rect -33 778 -17 812
rect 17 778 33 812
rect 141 799 175 880
rect -175 731 -141 765
rect -175 663 -141 697
rect -175 595 -141 629
rect -175 527 -141 561
rect -175 459 -141 493
rect -175 391 -141 425
rect -175 323 -141 357
rect -175 255 -141 289
rect -175 187 -141 221
rect -175 119 -141 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -175 -153 -141 -119
rect -175 -221 -141 -187
rect -175 -289 -141 -255
rect -175 -357 -141 -323
rect -175 -425 -141 -391
rect -175 -493 -141 -459
rect -175 -561 -141 -527
rect -175 -629 -141 -595
rect -175 -697 -141 -663
rect -175 -765 -141 -731
rect -61 701 -27 744
rect -61 629 -27 663
rect -61 561 -27 595
rect -61 493 -27 523
rect -61 425 -27 451
rect -61 357 -27 379
rect -61 289 -27 307
rect -61 221 -27 235
rect -61 153 -27 163
rect -61 85 -27 91
rect -61 17 -27 19
rect -61 -19 -27 -17
rect -61 -91 -27 -85
rect -61 -163 -27 -153
rect -61 -235 -27 -221
rect -61 -307 -27 -289
rect -61 -379 -27 -357
rect -61 -451 -27 -425
rect -61 -523 -27 -493
rect -61 -595 -27 -561
rect -61 -663 -27 -629
rect -61 -744 -27 -701
rect 27 701 61 744
rect 27 629 61 663
rect 27 561 61 595
rect 27 493 61 523
rect 27 425 61 451
rect 27 357 61 379
rect 27 289 61 307
rect 27 221 61 235
rect 27 153 61 163
rect 27 85 61 91
rect 27 17 61 19
rect 27 -19 61 -17
rect 27 -91 61 -85
rect 27 -163 61 -153
rect 27 -235 61 -221
rect 27 -307 61 -289
rect 27 -379 61 -357
rect 27 -451 61 -425
rect 27 -523 61 -493
rect 27 -595 61 -561
rect 27 -663 61 -629
rect 27 -744 61 -701
rect 141 731 175 765
rect 141 663 175 697
rect 141 595 175 629
rect 141 527 175 561
rect 141 459 175 493
rect 141 391 175 425
rect 141 323 175 357
rect 141 255 175 289
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
rect 141 -289 175 -255
rect 141 -357 175 -323
rect 141 -425 175 -391
rect 141 -493 175 -459
rect 141 -561 175 -527
rect 141 -629 175 -595
rect 141 -697 175 -663
rect 141 -765 175 -731
rect -175 -880 -141 -799
rect -33 -812 -17 -778
rect 17 -812 33 -778
rect 141 -880 175 -799
rect -175 -914 -51 -880
rect -17 -914 17 -880
rect 51 -914 175 -880
<< viali >>
rect -17 778 17 812
rect -61 697 -27 701
rect -61 667 -27 697
rect -61 595 -27 629
rect -61 527 -27 557
rect -61 523 -27 527
rect -61 459 -27 485
rect -61 451 -27 459
rect -61 391 -27 413
rect -61 379 -27 391
rect -61 323 -27 341
rect -61 307 -27 323
rect -61 255 -27 269
rect -61 235 -27 255
rect -61 187 -27 197
rect -61 163 -27 187
rect -61 119 -27 125
rect -61 91 -27 119
rect -61 51 -27 53
rect -61 19 -27 51
rect -61 -51 -27 -19
rect -61 -53 -27 -51
rect -61 -119 -27 -91
rect -61 -125 -27 -119
rect -61 -187 -27 -163
rect -61 -197 -27 -187
rect -61 -255 -27 -235
rect -61 -269 -27 -255
rect -61 -323 -27 -307
rect -61 -341 -27 -323
rect -61 -391 -27 -379
rect -61 -413 -27 -391
rect -61 -459 -27 -451
rect -61 -485 -27 -459
rect -61 -527 -27 -523
rect -61 -557 -27 -527
rect -61 -629 -27 -595
rect -61 -697 -27 -667
rect -61 -701 -27 -697
rect 27 697 61 701
rect 27 667 61 697
rect 27 595 61 629
rect 27 527 61 557
rect 27 523 61 527
rect 27 459 61 485
rect 27 451 61 459
rect 27 391 61 413
rect 27 379 61 391
rect 27 323 61 341
rect 27 307 61 323
rect 27 255 61 269
rect 27 235 61 255
rect 27 187 61 197
rect 27 163 61 187
rect 27 119 61 125
rect 27 91 61 119
rect 27 51 61 53
rect 27 19 61 51
rect 27 -51 61 -19
rect 27 -53 61 -51
rect 27 -119 61 -91
rect 27 -125 61 -119
rect 27 -187 61 -163
rect 27 -197 61 -187
rect 27 -255 61 -235
rect 27 -269 61 -255
rect 27 -323 61 -307
rect 27 -341 61 -323
rect 27 -391 61 -379
rect 27 -413 61 -391
rect 27 -459 61 -451
rect 27 -485 61 -459
rect 27 -527 61 -523
rect 27 -557 61 -527
rect 27 -629 61 -595
rect 27 -697 61 -667
rect 27 -701 61 -697
rect -17 -812 17 -778
<< metal1 >>
rect -29 812 29 818
rect -29 778 -17 812
rect 17 778 29 812
rect -29 772 29 778
rect -67 701 -21 740
rect -67 667 -61 701
rect -27 667 -21 701
rect -67 629 -21 667
rect -67 595 -61 629
rect -27 595 -21 629
rect -67 557 -21 595
rect -67 523 -61 557
rect -27 523 -21 557
rect -67 485 -21 523
rect -67 451 -61 485
rect -27 451 -21 485
rect -67 413 -21 451
rect -67 379 -61 413
rect -27 379 -21 413
rect -67 341 -21 379
rect -67 307 -61 341
rect -27 307 -21 341
rect -67 269 -21 307
rect -67 235 -61 269
rect -27 235 -21 269
rect -67 197 -21 235
rect -67 163 -61 197
rect -27 163 -21 197
rect -67 125 -21 163
rect -67 91 -61 125
rect -27 91 -21 125
rect -67 53 -21 91
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -91 -21 -53
rect -67 -125 -61 -91
rect -27 -125 -21 -91
rect -67 -163 -21 -125
rect -67 -197 -61 -163
rect -27 -197 -21 -163
rect -67 -235 -21 -197
rect -67 -269 -61 -235
rect -27 -269 -21 -235
rect -67 -307 -21 -269
rect -67 -341 -61 -307
rect -27 -341 -21 -307
rect -67 -379 -21 -341
rect -67 -413 -61 -379
rect -27 -413 -21 -379
rect -67 -451 -21 -413
rect -67 -485 -61 -451
rect -27 -485 -21 -451
rect -67 -523 -21 -485
rect -67 -557 -61 -523
rect -27 -557 -21 -523
rect -67 -595 -21 -557
rect -67 -629 -61 -595
rect -27 -629 -21 -595
rect -67 -667 -21 -629
rect -67 -701 -61 -667
rect -27 -701 -21 -667
rect -67 -740 -21 -701
rect 21 701 67 740
rect 21 667 27 701
rect 61 667 67 701
rect 21 629 67 667
rect 21 595 27 629
rect 61 595 67 629
rect 21 557 67 595
rect 21 523 27 557
rect 61 523 67 557
rect 21 485 67 523
rect 21 451 27 485
rect 61 451 67 485
rect 21 413 67 451
rect 21 379 27 413
rect 61 379 67 413
rect 21 341 67 379
rect 21 307 27 341
rect 61 307 67 341
rect 21 269 67 307
rect 21 235 27 269
rect 61 235 67 269
rect 21 197 67 235
rect 21 163 27 197
rect 61 163 67 197
rect 21 125 67 163
rect 21 91 27 125
rect 61 91 67 125
rect 21 53 67 91
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -91 67 -53
rect 21 -125 27 -91
rect 61 -125 67 -91
rect 21 -163 67 -125
rect 21 -197 27 -163
rect 61 -197 67 -163
rect 21 -235 67 -197
rect 21 -269 27 -235
rect 61 -269 67 -235
rect 21 -307 67 -269
rect 21 -341 27 -307
rect 61 -341 67 -307
rect 21 -379 67 -341
rect 21 -413 27 -379
rect 61 -413 67 -379
rect 21 -451 67 -413
rect 21 -485 27 -451
rect 61 -485 67 -451
rect 21 -523 67 -485
rect 21 -557 27 -523
rect 61 -557 67 -523
rect 21 -595 67 -557
rect 21 -629 27 -595
rect 61 -629 67 -595
rect 21 -667 67 -629
rect 21 -701 27 -667
rect 61 -701 67 -667
rect 21 -740 67 -701
rect -29 -778 29 -772
rect -29 -812 -17 -778
rect 17 -812 29 -778
rect -29 -818 29 -812
<< properties >>
string FIXED_BBOX -158 -897 158 897
<< end >>
