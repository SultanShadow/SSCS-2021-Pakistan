magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< metal3 >>
rect -112892 277247 -106540 278506
rect -112892 272223 -111987 277247
rect -107523 272223 -106540 277247
rect -112892 48598 -106540 272223
rect -63902 48598 2036 48704
rect -112994 43994 2036 48598
rect -112994 43888 -47056 43994
<< via3 >>
rect -111987 272223 -107523 277247
<< metal4 >>
rect -112562 277253 -106746 278124
rect -112562 277247 -111953 277253
rect -107557 277247 -106746 277253
rect -112562 272223 -111987 277247
rect -107523 272223 -106746 277247
rect -112562 272217 -111953 272223
rect -107557 272217 -106746 272223
rect -112562 271196 -106746 272217
rect -65094 234571 -56226 237548
rect -65094 225055 -62403 234571
rect -58327 225055 -56226 234571
rect -65094 68696 -56226 225055
rect -43588 68696 4524 68716
rect -65094 68544 4524 68696
rect -65094 65030 4688 68544
rect -65094 64738 4524 65030
rect -65094 64448 156 64738
<< via4 >>
rect -111953 277247 -107557 277253
rect -111953 272223 -107557 277247
rect -111953 272217 -107557 272223
rect -62403 225055 -58327 234571
<< metal5 >>
rect -112006 277253 -107504 277264
rect -112006 272217 -111953 277253
rect -107557 272217 -107504 277253
rect -112006 272206 -107504 272217
rect -62546 234571 -58184 234660
rect -62546 225055 -62403 234571
rect -58327 225055 -58184 234571
rect -62546 224966 -58184 225055
use WITHOUT_IND  WITHOUT_IND_0
timestamp 1636132012
transform 1 0 16 0 1 0
box -16 0 143952 98786
use INDUCTOR_layout  INDUCTOR_layout_0
timestamp 1636132012
transform 1 0 -902970 0 1 -2981242
box 788000 2884000 1344000 3262000
<< end >>
