magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< nwell >>
rect -338 -338 338 338
<< pwell >>
rect -466 380 466 466
rect -466 -380 -380 380
rect 380 -380 466 380
rect -466 -466 466 -380
<< psubdiff >>
rect -440 406 -323 440
rect -289 406 -255 440
rect -221 406 -187 440
rect -153 406 -119 440
rect -85 406 -51 440
rect -17 406 17 440
rect 51 406 85 440
rect 119 406 153 440
rect 187 406 221 440
rect 255 406 289 440
rect 323 406 440 440
rect -440 323 -406 406
rect 406 323 440 406
rect -440 255 -406 289
rect -440 187 -406 221
rect -440 119 -406 153
rect -440 51 -406 85
rect -440 -17 -406 17
rect -440 -85 -406 -51
rect -440 -153 -406 -119
rect -440 -221 -406 -187
rect -440 -289 -406 -255
rect 406 255 440 289
rect 406 187 440 221
rect 406 119 440 153
rect 406 51 440 85
rect 406 -17 440 17
rect 406 -85 440 -51
rect 406 -153 440 -119
rect 406 -221 440 -187
rect 406 -289 440 -255
rect -440 -406 -406 -323
rect 406 -406 440 -323
rect -440 -440 -323 -406
rect -289 -440 -255 -406
rect -221 -440 -187 -406
rect -153 -440 -119 -406
rect -85 -440 -51 -406
rect -17 -440 17 -406
rect 51 -440 85 -406
rect 119 -440 153 -406
rect 187 -440 221 -406
rect 255 -440 289 -406
rect 323 -440 440 -406
<< nsubdiff >>
rect -302 268 -187 302
rect -153 268 -119 302
rect -85 268 -51 302
rect -17 268 17 302
rect 51 268 85 302
rect 119 268 153 302
rect 187 268 302 302
rect -302 187 -268 268
rect -302 119 -268 153
rect -302 51 -268 85
rect -302 -17 -268 17
rect -302 -85 -268 -51
rect -302 -153 -268 -119
rect -302 -268 -268 -187
rect 268 187 302 268
rect 268 119 302 153
rect 268 51 302 85
rect 268 -17 302 17
rect 268 -85 302 -51
rect 268 -153 302 -119
rect 268 -268 302 -187
rect -302 -302 -187 -268
rect -153 -302 -119 -268
rect -85 -302 -51 -268
rect -17 -302 17 -268
rect 51 -302 85 -268
rect 119 -302 153 -268
rect 187 -302 302 -268
<< psubdiffcont >>
rect -323 406 -289 440
rect -255 406 -221 440
rect -187 406 -153 440
rect -119 406 -85 440
rect -51 406 -17 440
rect 17 406 51 440
rect 85 406 119 440
rect 153 406 187 440
rect 221 406 255 440
rect 289 406 323 440
rect -440 289 -406 323
rect -440 221 -406 255
rect -440 153 -406 187
rect -440 85 -406 119
rect -440 17 -406 51
rect -440 -51 -406 -17
rect -440 -119 -406 -85
rect -440 -187 -406 -153
rect -440 -255 -406 -221
rect -440 -323 -406 -289
rect 406 289 440 323
rect 406 221 440 255
rect 406 153 440 187
rect 406 85 440 119
rect 406 17 440 51
rect 406 -51 440 -17
rect 406 -119 440 -85
rect 406 -187 440 -153
rect 406 -255 440 -221
rect 406 -323 440 -289
rect -323 -440 -289 -406
rect -255 -440 -221 -406
rect -187 -440 -153 -406
rect -119 -440 -85 -406
rect -51 -440 -17 -406
rect 17 -440 51 -406
rect 85 -440 119 -406
rect 153 -440 187 -406
rect 221 -440 255 -406
rect 289 -440 323 -406
<< nsubdiffcont >>
rect -187 268 -153 302
rect -119 268 -85 302
rect -51 268 -17 302
rect 17 268 51 302
rect 85 268 119 302
rect 153 268 187 302
rect -302 153 -268 187
rect -302 85 -268 119
rect -302 17 -268 51
rect -302 -51 -268 -17
rect -302 -119 -268 -85
rect -302 -187 -268 -153
rect 268 153 302 187
rect 268 85 302 119
rect 268 17 302 51
rect 268 -51 302 -17
rect 268 -119 302 -85
rect 268 -187 302 -153
rect -187 -302 -153 -268
rect -119 -302 -85 -268
rect -51 -302 -17 -268
rect 17 -302 51 -268
rect 85 -302 119 -268
rect 153 -302 187 -268
<< pdiode >>
rect -200 187 200 200
rect -200 -187 -187 187
rect 187 -187 200 187
rect -200 -200 200 -187
<< pdiodec >>
rect -187 -187 187 187
<< locali >>
rect -440 406 -323 440
rect -289 406 -255 440
rect -221 406 -187 440
rect -153 406 -119 440
rect -85 406 -51 440
rect -17 406 17 440
rect 51 406 85 440
rect 119 406 153 440
rect 187 406 221 440
rect 255 406 289 440
rect 323 406 440 440
rect -440 323 -406 406
rect 406 323 440 406
rect -440 255 -406 289
rect -440 187 -406 221
rect -440 119 -406 153
rect -440 51 -406 85
rect -440 -17 -406 17
rect -440 -85 -406 -51
rect -440 -153 -406 -119
rect -440 -221 -406 -187
rect -440 -289 -406 -255
rect -302 268 -187 302
rect -153 268 -119 302
rect -85 268 -51 302
rect -17 268 17 302
rect 51 268 85 302
rect 119 268 153 302
rect 187 268 302 302
rect -302 187 -268 268
rect -302 119 -268 153
rect -302 51 -268 85
rect -302 -17 -268 17
rect -302 -85 -268 -51
rect -302 -153 -268 -119
rect -302 -268 -268 -187
rect -204 187 204 188
rect -204 -187 -187 187
rect 187 -187 204 187
rect -204 -188 204 -187
rect 268 187 302 268
rect 268 119 302 153
rect 268 51 302 85
rect 268 -17 302 17
rect 268 -85 302 -51
rect 268 -153 302 -119
rect 268 -268 302 -187
rect -302 -302 -187 -268
rect -153 -302 -119 -268
rect -85 -302 -51 -268
rect -17 -302 17 -268
rect 51 -302 85 -268
rect 119 -302 153 -268
rect 187 -302 302 -268
rect 406 255 440 289
rect 406 187 440 221
rect 406 119 440 153
rect 406 51 440 85
rect 406 -17 440 17
rect 406 -85 440 -51
rect 406 -153 440 -119
rect 406 -221 440 -187
rect 406 -289 440 -255
rect -440 -406 -406 -323
rect 406 -406 440 -323
rect -440 -440 -323 -406
rect -289 -440 -255 -406
rect -221 -440 -187 -406
rect -153 -440 -119 -406
rect -85 -440 -51 -406
rect -17 -440 17 -406
rect 51 -440 85 -406
rect 119 -440 153 -406
rect 187 -440 221 -406
rect 255 -440 289 -406
rect 323 -440 440 -406
<< viali >>
rect -161 -161 161 161
<< metal1 >>
rect -200 161 200 194
rect -200 -161 -161 161
rect 161 -161 200 161
rect -200 -194 200 -161
<< properties >>
string FIXED_BBOX -284 -284 284 284
<< end >>
