magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< locali >>
rect 6239 21889 6632 22186
rect 9068 21889 9341 21898
rect 6239 21886 9341 21889
rect 6240 20081 9341 21886
rect 9068 12151 9341 20081
rect 8251 10317 9292 10790
rect 8251 7547 9663 10317
rect 21766 301 22279 324
rect 21710 288 22336 301
rect 7675 -812 8880 278
rect 21710 182 21789 288
rect 22255 182 22336 288
rect 21710 113 22336 182
rect 7675 -918 7758 -812
rect 8800 -918 8880 -812
rect 7675 -1008 8880 -918
<< viali >>
rect 21789 182 22255 288
rect 7758 -918 8800 -812
<< metal1 >>
rect 10100 20784 10686 22109
rect 10100 20604 10256 20784
rect 10564 20604 10686 20784
rect 10100 20465 10686 20604
rect 20916 20774 22367 20923
rect 20916 20594 21187 20774
rect 22135 20594 22367 20774
rect 16137 19908 16203 19932
rect 20916 19807 22367 20594
rect 20916 19653 22363 19807
rect 20916 19281 21030 19653
rect 22234 19281 22363 19653
rect 4746 11413 4769 11548
rect 18350 11430 18372 11611
rect 20916 7963 22363 19281
rect 20916 7832 22626 7963
rect 20916 7268 21111 7832
rect 22187 7268 22626 7832
rect 20916 7115 22626 7268
rect 24154 7527 25284 7716
rect 24154 7091 24444 7527
rect 25072 7091 25284 7527
rect 25714 7231 26132 7265
rect 24154 6862 25284 7091
rect 9299 6447 25286 6862
rect 9068 5733 9096 5740
rect 6847 3355 6851 3373
rect 14495 1810 14806 4002
rect 11512 1551 11518 1617
rect 7796 1379 13978 1473
rect 7796 1058 13373 1379
rect 10586 385 10590 455
rect 13282 -209 13373 1058
rect 13873 -209 13978 1379
rect 17168 192 17605 391
rect 21669 288 22340 386
rect 13282 -292 13978 -209
rect 21669 182 21789 288
rect 22255 182 22340 288
rect 21669 -704 22340 182
rect 23385 45 23833 52
rect 23385 13 23833 29
rect 17168 -707 22340 -704
rect 7675 -812 22340 -707
rect 7675 -918 7758 -812
rect 8800 -918 22340 -812
rect 7675 -1008 22340 -918
<< via1 >>
rect 10256 20604 10564 20784
rect 21187 20594 22135 20774
rect 21030 19281 22234 19653
rect 21111 7268 22187 7832
rect 24444 7091 25072 7527
rect 13373 -209 13873 1379
<< metal2 >>
rect 3161 21130 3210 21778
rect 20783 20916 22367 20923
rect 6644 20784 22367 20916
rect 6644 20604 10256 20784
rect 10564 20774 22367 20784
rect 10564 20604 21187 20774
rect 6644 20594 21187 20604
rect 22135 20594 22367 20774
rect 6644 20465 22367 20594
rect 16989 20059 17135 20076
rect 18489 19653 22363 19808
rect 18489 19281 21030 19653
rect 22234 19281 22363 19653
rect 18489 19142 22363 19281
rect 9900 16840 11015 17236
rect 9900 13264 10212 16840
rect 10748 13264 11015 16840
rect 9900 12902 11015 13264
rect 11647 13307 18207 13554
rect 11647 13011 14247 13307
rect 17183 13011 18207 13307
rect 11647 12869 18207 13011
rect 10511 9633 19534 9763
rect 10511 9257 18118 9633
rect 18974 9257 19534 9633
rect 10511 9115 19534 9257
rect 11424 7832 22630 7965
rect 11424 7268 21111 7832
rect 22187 7268 22630 7832
rect 11424 7115 22630 7268
rect 23139 7641 23744 7784
rect 23139 7345 23294 7641
rect 23590 7345 23744 7641
rect 23139 6948 23744 7345
rect 24154 7527 25284 7716
rect 24154 7091 24444 7527
rect 25072 7091 25284 7527
rect 24154 7021 25284 7091
rect 17187 2947 18219 2955
rect 12450 1979 19290 2947
rect 17187 1529 18219 1979
rect 13282 1379 13978 1473
rect 13282 1373 13373 1379
rect 13873 1373 13978 1379
rect 13282 -203 13355 1373
rect 13891 -203 13978 1373
rect 13282 -209 13373 -203
rect 13873 -209 13978 -203
rect 13282 -292 13978 -209
<< via2 >>
rect 10212 13264 10748 16840
rect 14247 13011 17183 13307
rect 18118 9257 18974 9633
rect 23294 7345 23590 7641
rect 24450 7121 25066 7497
rect 13355 -203 13373 1373
rect 13373 -203 13873 1373
rect 13873 -203 13891 1373
<< metal3 >>
rect 9899 16844 11015 17237
rect 9899 13260 10208 16844
rect 10752 13260 11015 16844
rect 9899 12902 11015 13260
rect 13560 13311 18058 13554
rect 13560 13007 14243 13311
rect 17187 13007 18058 13311
rect 13560 12869 18058 13007
rect 18012 9637 19175 9763
rect 18012 9253 18114 9637
rect 18978 9253 19175 9637
rect 18012 9115 19175 9253
rect 23139 7645 23744 7784
rect 23139 7341 23290 7645
rect 23594 7341 23744 7645
rect 23139 7203 23744 7341
rect 24154 7501 25284 7716
rect 24154 7117 24446 7501
rect 25070 7117 25284 7501
rect 24154 7021 25284 7117
rect 13282 1377 13978 1473
rect 13282 -207 13351 1377
rect 13895 -207 13978 1377
rect 13282 -292 13978 -207
<< via3 >>
rect 10208 16840 10752 16844
rect 10208 13264 10212 16840
rect 10212 13264 10748 16840
rect 10748 13264 10752 16840
rect 10208 13260 10752 13264
rect 14243 13307 17187 13311
rect 14243 13011 14247 13307
rect 14247 13011 17183 13307
rect 17183 13011 17187 13307
rect 14243 13007 17187 13011
rect 18114 9633 18978 9637
rect 18114 9257 18118 9633
rect 18118 9257 18974 9633
rect 18974 9257 18978 9633
rect 18114 9253 18978 9257
rect 23290 7641 23594 7645
rect 23290 7345 23294 7641
rect 23294 7345 23590 7641
rect 23590 7345 23594 7641
rect 23290 7341 23594 7345
rect 24446 7497 25070 7501
rect 24446 7121 24450 7497
rect 24450 7121 25066 7497
rect 25066 7121 25070 7497
rect 24446 7117 25070 7121
rect 13351 1373 13895 1377
rect 13351 -203 13355 1373
rect 13355 -203 13891 1373
rect 13891 -203 13895 1373
rect 13351 -207 13895 -203
<< metal4 >>
rect 9899 16844 11015 17237
rect 9899 13260 10208 16844
rect 10752 13260 11015 16844
rect 9899 12902 11015 13260
rect 13560 13311 18058 13554
rect 13560 13007 14243 13311
rect 17187 13007 18058 13311
rect 13560 12869 18058 13007
rect 18012 9637 19576 9763
rect 18012 9253 18114 9637
rect 18978 9253 19576 9637
rect 18012 9115 19576 9253
rect 23139 7645 23744 7784
rect 23139 7341 23290 7645
rect 23594 7341 23744 7645
rect 23139 7203 23744 7341
rect 24154 7501 25284 7716
rect 24154 7117 24446 7501
rect 25070 7117 25284 7501
rect 24154 7021 25284 7117
rect 13282 1377 13978 1473
rect 13282 1343 13351 1377
rect 13895 1343 13978 1377
rect 13282 -173 13345 1343
rect 13901 -173 13978 1343
rect 13282 -207 13351 -173
rect 13895 -207 13978 -173
rect 13282 -292 13978 -207
<< via4 >>
rect 14317 13041 14553 13277
rect 14637 13041 14873 13277
rect 14957 13041 15193 13277
rect 15277 13041 15513 13277
rect 15597 13041 15833 13277
rect 15917 13041 16153 13277
rect 16237 13041 16473 13277
rect 16557 13041 16793 13277
rect 16877 13041 17113 13277
rect 23324 7375 23560 7611
rect 24480 7191 24716 7427
rect 24800 7191 25036 7427
rect 13345 -173 13351 1343
rect 13351 -173 13895 1343
rect 13895 -173 13901 1343
<< metal5 >>
rect 13560 13277 18058 15016
rect 13560 13041 14317 13277
rect 14553 13041 14637 13277
rect 14873 13041 14957 13277
rect 15193 13041 15277 13277
rect 15513 13041 15597 13277
rect 15833 13041 15917 13277
rect 16153 13041 16237 13277
rect 16473 13041 16557 13277
rect 16793 13041 16877 13277
rect 17113 13041 18058 13277
rect 13560 12869 18058 13041
rect 18064 9115 19576 9763
rect 23139 7611 23744 8578
rect 23139 7375 23324 7611
rect 23560 7375 23744 7611
rect 23139 7203 23744 7375
rect 24154 7427 25284 7716
rect 24154 7191 24480 7427
rect 24716 7191 24800 7427
rect 25036 7191 25284 7427
rect 24154 6650 25284 7191
rect 13282 1343 15152 1473
rect 13282 -173 13345 1343
rect 13901 -173 15152 1343
rect 13282 -292 15152 -173
use PA_BUFF  PA_BUFF_0
timestamp 1636132012
transform 1 0 3802 0 -1 21092
box -641 -1212 6958 8136
use Switch  Switch_0
timestamp 1636132012
transform 1 0 10953 0 1 9891
box -6207 -129 7419 3455
use LNA_2ndstage  LNA_2ndstage_0
timestamp 1636132012
transform 1 0 20364 0 1 902
box -6280 -889 7501 7084
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1636132012
transform -1 0 22629 0 1 11359
box -3351 -3101 3373 3101
use LNA_Buff  LNA_Buff_0
timestamp 1636132012
transform -1 0 18309 0 1 18676
box -466 -5034 6978 1638
use LNA  LNA_0
timestamp 1636132012
transform 1 0 6847 0 1 2730
box -6847 -2730 6094 5235
<< labels >>
rlabel metal1 s 4747 11473 4747 11473 4 VSWN
port 1 nsew
rlabel metal1 s 18368 11505 18368 11505 4 VSWP
port 2 nsew
rlabel metal1 s 10685 21626 10685 21626 4 VDD
port 3 nsew
rlabel metal1 s 11517 1585 11517 1585 4 VBIAS1
port 4 nsew
rlabel metal1 s 9082 5739 9082 5739 4 VSS
port 5 nsew
rlabel metal1 s 6847 3362 6847 3362 4 VCASC1
port 6 nsew
rlabel metal1 s 10589 416 10589 416 4 VBIAS2
port 7 nsew
rlabel metal1 s 23636 16 23636 16 4 VBIAS3
port 8 nsew
rlabel metal1 s 25902 7253 25902 7253 4 VCASC2
port 9 nsew
rlabel metal2 s 17068 20074 17068 20074 4 RFOUTLNA
port 10 nsew
rlabel metal1 s 16171 19930 16171 19930 4 VBIAS4
port 11 nsew
rlabel metal2 s 3161 21423 3161 21423 4 RFOUTPA
port 12 nsew
<< end >>
