magic
tech sky130A
magscale 1 2
timestamp 1636132012
<< locali >>
rect -44 8214 9194 8270
rect -44 8212 5634 8214
rect -44 8210 3784 8212
rect -44 8208 1014 8210
rect -44 8198 90 8208
rect 232 8206 1014 8208
rect 232 8198 548 8206
rect 690 8198 1014 8206
rect 1156 8204 1936 8210
rect 1156 8198 1476 8204
rect 1618 8198 1936 8204
rect 2078 8208 2862 8210
rect 2078 8198 2398 8208
rect 2540 8198 2862 8208
rect 3004 8198 3324 8210
rect 3466 8198 3784 8210
rect 3926 8210 5634 8212
rect 3926 8206 4708 8210
rect 3926 8198 4246 8206
rect 4388 8198 4708 8206
rect 4850 8198 5168 8210
rect 5310 8198 5634 8210
rect 5776 8198 6096 8214
rect 6238 8212 9194 8214
rect 6238 8198 6556 8212
rect 6698 8210 7942 8212
rect 6698 8208 7482 8210
rect 6698 8198 7018 8208
rect 7160 8198 7482 8208
rect 7624 8198 7942 8210
rect 8084 8198 8404 8212
rect 8546 8198 8868 8212
rect 9010 8198 9194 8212
rect -52 -8038 88 -8028
rect 230 -8036 550 -8028
rect 692 -8036 1014 -8028
rect 1156 -8034 1478 -8028
rect 1620 -8034 1936 -8028
rect 2078 -8034 2400 -8028
rect 1156 -8036 2400 -8034
rect 2542 -8032 2862 -8028
rect 3004 -8032 3322 -8028
rect 2542 -8034 3322 -8032
rect 3464 -8034 3786 -8028
rect 3928 -8034 4250 -8028
rect 2542 -8036 4250 -8034
rect 4392 -8034 4712 -8028
rect 4854 -8034 5172 -8028
rect 5314 -8034 5636 -8028
rect 5778 -8032 6096 -8028
rect 6238 -8032 6558 -8028
rect 5778 -8034 6558 -8032
rect 4392 -8036 6558 -8034
rect 6700 -8032 7022 -8028
rect 7164 -8032 7484 -8028
rect 7626 -8032 7942 -8028
rect 6700 -8034 7942 -8032
rect 8084 -8034 8402 -8028
rect 8544 -8034 8868 -8028
rect 9010 -8034 9158 -8028
rect 6700 -8036 9158 -8034
rect 230 -8038 9158 -8036
rect -52 -8116 9158 -8038
<< metal1 >>
rect 120 8118 9114 8286
rect -166 8042 112 8072
rect -166 7990 -113 8042
rect -61 7990 -49 8042
rect 3 7990 112 8042
rect -166 7954 112 7990
rect 430 8037 572 8072
rect 430 7985 460 8037
rect 512 7985 572 8037
rect 430 7954 572 7985
rect 890 8055 1034 8068
rect 890 8003 940 8055
rect 992 8003 1034 8055
rect 890 7952 1034 8003
rect 1354 8047 1496 8074
rect 1354 7995 1388 8047
rect 1440 7995 1496 8047
rect 1354 7950 1496 7995
rect 1806 8039 1962 8074
rect 1806 7987 1836 8039
rect 1888 7987 1962 8039
rect 1806 7940 1962 7987
rect 2278 8049 2422 8074
rect 2278 7997 2304 8049
rect 2356 7997 2422 8049
rect 2278 7942 2422 7997
rect 2732 8049 2884 8078
rect 2732 7997 2764 8049
rect 2816 7997 2884 8049
rect 2732 7940 2884 7997
rect 3200 8045 3350 8080
rect 3200 7993 3232 8045
rect 3284 7993 3350 8045
rect 3200 7942 3350 7993
rect 3702 8025 3808 8084
rect 3702 7973 3734 8025
rect 3786 7973 3808 8025
rect 3702 7942 3808 7973
rect 4122 8041 4272 8084
rect 4122 7989 4164 8041
rect 4216 7989 4272 8041
rect 4122 7950 4272 7989
rect 4582 8049 4732 8078
rect 4582 7997 4616 8049
rect 4668 7997 4732 8049
rect 4582 7954 4732 7997
rect 5082 8035 5196 8084
rect 5082 7983 5096 8035
rect 5148 7983 5196 8035
rect 5082 7950 5196 7983
rect 5512 8033 5654 8086
rect 5512 7981 5542 8033
rect 5594 7981 5654 8033
rect 5512 7948 5654 7981
rect 5970 8055 6118 8084
rect 5970 8003 6024 8055
rect 6076 8003 6118 8055
rect 5970 7968 6118 8003
rect 6434 8049 6574 8086
rect 6434 7997 6468 8049
rect 6520 7997 6574 8049
rect 6434 7966 6574 7997
rect 6896 8049 7040 8082
rect 6896 7997 6926 8049
rect 6978 7997 7040 8049
rect 6896 7962 7040 7997
rect 7392 8043 7504 8070
rect 7392 7991 7418 8043
rect 7470 7991 7504 8043
rect 7392 7962 7504 7991
rect 7854 8051 7964 8066
rect 7854 7999 7878 8051
rect 7930 7999 7964 8051
rect 7854 7966 7964 7999
rect 8316 8061 8426 8074
rect 8316 8009 8342 8061
rect 8394 8009 8426 8061
rect 8316 7964 8426 8009
rect 8750 8049 8888 8072
rect 8750 7997 8768 8049
rect 8820 7997 8888 8049
rect 8750 7964 8888 7997
rect 204 -7831 316 -7790
rect 204 -7883 244 -7831
rect 296 -7883 316 -7831
rect 204 -7906 316 -7883
rect 666 -7817 788 -7788
rect 666 -7869 706 -7817
rect 758 -7869 788 -7817
rect 666 -7906 788 -7869
rect 1118 -7817 1242 -7786
rect 1118 -7869 1162 -7817
rect 1214 -7869 1242 -7817
rect 1118 -7916 1242 -7869
rect 1590 -7821 1708 -7780
rect 1590 -7873 1626 -7821
rect 1678 -7873 1708 -7821
rect 1590 -7916 1708 -7873
rect 2046 -7813 2166 -7782
rect 2046 -7865 2082 -7813
rect 2134 -7865 2166 -7813
rect 2046 -7916 2166 -7865
rect 2504 -7823 2632 -7776
rect 2504 -7875 2550 -7823
rect 2602 -7875 2632 -7823
rect 2504 -7916 2632 -7875
rect 2964 -7803 3092 -7770
rect 2964 -7855 3024 -7803
rect 3076 -7855 3092 -7803
rect 2964 -7918 3092 -7855
rect 3430 -7815 3558 -7774
rect 3430 -7867 3474 -7815
rect 3526 -7867 3558 -7815
rect 3430 -7918 3558 -7867
rect 3894 -7813 4018 -7770
rect 3894 -7865 3946 -7813
rect 3998 -7865 4018 -7813
rect 3894 -7920 4018 -7865
rect 4354 -7805 4484 -7768
rect 4354 -7857 4410 -7805
rect 4462 -7857 4484 -7805
rect 4354 -7916 4484 -7857
rect 4814 -7805 4942 -7760
rect 4814 -7857 4872 -7805
rect 4924 -7857 4942 -7805
rect 4814 -7918 4942 -7857
rect 5292 -7795 5434 -7766
rect 5292 -7847 5324 -7795
rect 5376 -7847 5434 -7795
rect 5292 -7902 5434 -7847
rect 5752 -7811 5898 -7764
rect 5752 -7863 5782 -7811
rect 5834 -7863 5898 -7811
rect 5752 -7920 5898 -7863
rect 6214 -7799 6362 -7768
rect 6214 -7851 6254 -7799
rect 6306 -7851 6362 -7799
rect 6214 -7902 6362 -7851
rect 6674 -7793 6824 -7764
rect 6674 -7845 6748 -7793
rect 6800 -7845 6824 -7793
rect 6674 -7906 6824 -7845
rect 7136 -7787 7290 -7766
rect 7136 -7839 7194 -7787
rect 7246 -7839 7290 -7787
rect 7136 -7920 7290 -7839
rect 7600 -7793 7744 -7772
rect 7600 -7845 7658 -7793
rect 7710 -7845 7744 -7793
rect 7600 -7902 7744 -7845
rect 8060 -7795 8216 -7768
rect 8060 -7847 8120 -7795
rect 8172 -7847 8216 -7795
rect 8060 -7900 8216 -7847
rect 8520 -7797 8670 -7778
rect 8520 -7849 8578 -7797
rect 8630 -7849 8670 -7797
rect 8520 -7902 8670 -7849
rect 8986 -7801 9138 -7762
rect 8986 -7853 9038 -7801
rect 9090 -7853 9138 -7801
rect 8986 -7906 9138 -7853
rect 114 -8222 9138 -7950
<< via1 >>
rect -113 7990 -61 8042
rect -49 7990 3 8042
rect 460 7985 512 8037
rect 940 8003 992 8055
rect 1388 7995 1440 8047
rect 1836 7987 1888 8039
rect 2304 7997 2356 8049
rect 2764 7997 2816 8049
rect 3232 7993 3284 8045
rect 3734 7973 3786 8025
rect 4164 7989 4216 8041
rect 4616 7997 4668 8049
rect 5096 7983 5148 8035
rect 5542 7981 5594 8033
rect 6024 8003 6076 8055
rect 6468 7997 6520 8049
rect 6926 7997 6978 8049
rect 7418 7991 7470 8043
rect 7878 7999 7930 8051
rect 8342 8009 8394 8061
rect 8768 7997 8820 8049
rect 244 -7883 296 -7831
rect 706 -7869 758 -7817
rect 1162 -7869 1214 -7817
rect 1626 -7873 1678 -7821
rect 2082 -7865 2134 -7813
rect 2550 -7875 2602 -7823
rect 3024 -7855 3076 -7803
rect 3474 -7867 3526 -7815
rect 3946 -7865 3998 -7813
rect 4410 -7857 4462 -7805
rect 4872 -7857 4924 -7805
rect 5324 -7847 5376 -7795
rect 5782 -7863 5834 -7811
rect 6254 -7851 6306 -7799
rect 6748 -7845 6800 -7793
rect 7194 -7839 7246 -7787
rect 7658 -7845 7710 -7793
rect 8120 -7847 8172 -7795
rect 8578 -7849 8630 -7797
rect 9038 -7853 9090 -7801
<< metal2 >>
rect 2278 8084 2884 8088
rect 4602 8086 5194 8088
rect 6026 8086 6576 8088
rect 3200 8084 3810 8086
rect 2278 8080 4274 8084
rect 4602 8080 7040 8086
rect -166 8072 572 8078
rect 2278 8074 7040 8080
rect 1398 8072 7040 8074
rect 7864 8082 8426 8086
rect 7864 8072 8890 8082
rect -166 8061 8890 8072
rect -166 8055 8342 8061
rect -166 8042 940 8055
rect -166 7990 -113 8042
rect -61 7990 -49 8042
rect 3 8037 940 8042
rect 3 7990 460 8037
rect -166 7985 460 7990
rect 512 8003 940 8037
rect 992 8049 6024 8055
rect 992 8047 2304 8049
rect 992 8003 1388 8047
rect 512 7995 1388 8003
rect 1440 8039 2304 8047
rect 1440 7995 1836 8039
rect 512 7987 1836 7995
rect 1888 7997 2304 8039
rect 2356 7997 2764 8049
rect 2816 8045 4616 8049
rect 2816 7997 3232 8045
rect 1888 7993 3232 7997
rect 3284 8041 4616 8045
rect 3284 8025 4164 8041
rect 3284 7993 3734 8025
rect 1888 7987 3734 7993
rect 512 7985 3734 7987
rect -166 7973 3734 7985
rect 3786 7989 4164 8025
rect 4216 7997 4616 8041
rect 4668 8035 6024 8049
rect 4668 7997 5096 8035
rect 4216 7989 5096 7997
rect 3786 7983 5096 7989
rect 5148 8033 6024 8035
rect 5148 7983 5542 8033
rect 3786 7981 5542 7983
rect 5594 8003 6024 8033
rect 6076 8051 8342 8055
rect 6076 8049 7878 8051
rect 6076 8003 6468 8049
rect 5594 7997 6468 8003
rect 6520 7997 6926 8049
rect 6978 8043 7878 8049
rect 6978 7997 7418 8043
rect 5594 7991 7418 7997
rect 7470 7999 7878 8043
rect 7930 8009 8342 8051
rect 8394 8049 8890 8061
rect 8394 8009 8768 8049
rect 7930 7999 8768 8009
rect 7470 7997 8768 7999
rect 8820 7997 8890 8049
rect 7470 7991 8890 7997
rect 5594 7981 8890 7991
rect 3786 7973 8890 7981
rect -166 7968 8890 7973
rect -166 7954 5656 7968
rect 6026 7964 8890 7968
rect 6432 7962 8426 7964
rect 6432 7960 7506 7962
rect 928 7952 5656 7954
rect 928 7950 4274 7952
rect 1398 7948 4274 7950
rect 5084 7948 5656 7952
rect 1398 7942 3810 7948
rect 1910 7940 2884 7942
rect 2278 7938 2884 7940
rect 3200 7938 3810 7942
rect 6212 -7762 6826 -7760
rect 4360 -7766 7290 -7762
rect 8522 -7764 9136 -7760
rect 8064 -7766 9136 -7764
rect 3892 -7768 9136 -7766
rect 3428 -7770 9136 -7768
rect 2962 -7774 9136 -7770
rect 2502 -7778 9136 -7774
rect 1588 -7782 9136 -7778
rect 1126 -7786 9136 -7782
rect 692 -7787 9136 -7786
rect 692 -7790 7194 -7787
rect -308 -7793 7194 -7790
rect -308 -7795 6748 -7793
rect -308 -7803 5324 -7795
rect -308 -7813 3024 -7803
rect -308 -7817 2082 -7813
rect -308 -7831 706 -7817
rect -308 -7883 244 -7831
rect 296 -7869 706 -7831
rect 758 -7869 1162 -7817
rect 1214 -7821 2082 -7817
rect 1214 -7869 1626 -7821
rect 296 -7873 1626 -7869
rect 1678 -7865 2082 -7821
rect 2134 -7823 3024 -7813
rect 2134 -7865 2550 -7823
rect 1678 -7873 2550 -7865
rect 296 -7875 2550 -7873
rect 2602 -7855 3024 -7823
rect 3076 -7805 5324 -7803
rect 3076 -7813 4410 -7805
rect 3076 -7815 3946 -7813
rect 3076 -7855 3474 -7815
rect 2602 -7867 3474 -7855
rect 3526 -7865 3946 -7815
rect 3998 -7857 4410 -7813
rect 4462 -7857 4872 -7805
rect 4924 -7847 5324 -7805
rect 5376 -7799 6748 -7795
rect 5376 -7811 6254 -7799
rect 5376 -7847 5782 -7811
rect 4924 -7857 5782 -7847
rect 3998 -7863 5782 -7857
rect 5834 -7851 6254 -7811
rect 6306 -7845 6748 -7799
rect 6800 -7839 7194 -7793
rect 7246 -7793 9136 -7787
rect 7246 -7839 7658 -7793
rect 6800 -7845 7658 -7839
rect 7710 -7795 9136 -7793
rect 7710 -7845 8120 -7795
rect 6306 -7847 8120 -7845
rect 8172 -7797 9136 -7795
rect 8172 -7847 8578 -7797
rect 6306 -7849 8578 -7847
rect 8630 -7801 9136 -7797
rect 8630 -7849 9038 -7801
rect 6306 -7851 9038 -7849
rect 5834 -7853 9038 -7851
rect 9090 -7853 9136 -7801
rect 5834 -7863 9136 -7853
rect 3998 -7865 9136 -7863
rect 3526 -7867 9136 -7865
rect 2602 -7875 9136 -7867
rect 296 -7883 9136 -7875
rect -308 -7906 9136 -7883
rect 692 -7916 9136 -7906
rect 2036 -7918 9136 -7916
rect 2502 -7920 9136 -7918
rect 3428 -7924 4018 -7920
rect 4360 -7922 9136 -7920
rect 4814 -7924 5900 -7922
rect 7132 -7924 9136 -7922
rect 4814 -7926 5438 -7924
use sky130_fd_pr__nfet_01v8_lvt_BPY4AF  sky130_fd_pr__nfet_01v8_lvt_BPY4AF_0
array 19 0 462 0 0 16420
timestamp 1636132012
transform 1 0 159 0 1 85
box -221 -8200 221 8200
<< labels >>
rlabel locali s -14 8224 -14 8224 4 B
port 1 nsew
rlabel metal1 s 242 8152 242 8152 4 G
port 2 nsew
rlabel metal2 s -142 8020 -142 8020 4 D
port 3 nsew
rlabel metal2 s -204 -7864 -204 -7864 4 S
port 4 nsew
<< end >>
