magic
tech sky130A
magscale 1 2
timestamp 1635855079
<< error_p >>
rect -6389 6350 -6329 12550
rect -6309 6350 -6249 12550
rect -70 6350 -10 12550
rect 10 6350 70 12550
rect 6249 6350 6309 12550
rect 6329 6350 6389 12550
rect -6389 50 -6329 6250
rect -6309 50 -6249 6250
rect -70 50 -10 6250
rect 10 50 70 6250
rect 6249 50 6309 6250
rect 6329 50 6389 6250
rect -6389 -6250 -6329 -50
rect -6309 -6250 -6249 -50
rect -70 -6250 -10 -50
rect 10 -6250 70 -50
rect 6249 -6250 6309 -50
rect 6329 -6250 6389 -50
rect -6389 -12550 -6329 -6350
rect -6309 -12550 -6249 -6350
rect -70 -12550 -10 -6350
rect 10 -12550 70 -6350
rect 6249 -12550 6309 -6350
rect 6329 -12550 6389 -6350
<< metal3 >>
rect -12628 12522 -6329 12550
rect -12628 12458 -6413 12522
rect -6349 12458 -6329 12522
rect -12628 12442 -6329 12458
rect -12628 12378 -6413 12442
rect -6349 12378 -6329 12442
rect -12628 12362 -6329 12378
rect -12628 12298 -6413 12362
rect -6349 12298 -6329 12362
rect -12628 12282 -6329 12298
rect -12628 12218 -6413 12282
rect -6349 12218 -6329 12282
rect -12628 12202 -6329 12218
rect -12628 12138 -6413 12202
rect -6349 12138 -6329 12202
rect -12628 12122 -6329 12138
rect -12628 12058 -6413 12122
rect -6349 12058 -6329 12122
rect -12628 12042 -6329 12058
rect -12628 11978 -6413 12042
rect -6349 11978 -6329 12042
rect -12628 11962 -6329 11978
rect -12628 11898 -6413 11962
rect -6349 11898 -6329 11962
rect -12628 11882 -6329 11898
rect -12628 11818 -6413 11882
rect -6349 11818 -6329 11882
rect -12628 11802 -6329 11818
rect -12628 11738 -6413 11802
rect -6349 11738 -6329 11802
rect -12628 11722 -6329 11738
rect -12628 11658 -6413 11722
rect -6349 11658 -6329 11722
rect -12628 11642 -6329 11658
rect -12628 11578 -6413 11642
rect -6349 11578 -6329 11642
rect -12628 11562 -6329 11578
rect -12628 11498 -6413 11562
rect -6349 11498 -6329 11562
rect -12628 11482 -6329 11498
rect -12628 11418 -6413 11482
rect -6349 11418 -6329 11482
rect -12628 11402 -6329 11418
rect -12628 11338 -6413 11402
rect -6349 11338 -6329 11402
rect -12628 11322 -6329 11338
rect -12628 11258 -6413 11322
rect -6349 11258 -6329 11322
rect -12628 11242 -6329 11258
rect -12628 11178 -6413 11242
rect -6349 11178 -6329 11242
rect -12628 11162 -6329 11178
rect -12628 11098 -6413 11162
rect -6349 11098 -6329 11162
rect -12628 11082 -6329 11098
rect -12628 11018 -6413 11082
rect -6349 11018 -6329 11082
rect -12628 11002 -6329 11018
rect -12628 10938 -6413 11002
rect -6349 10938 -6329 11002
rect -12628 10922 -6329 10938
rect -12628 10858 -6413 10922
rect -6349 10858 -6329 10922
rect -12628 10842 -6329 10858
rect -12628 10778 -6413 10842
rect -6349 10778 -6329 10842
rect -12628 10762 -6329 10778
rect -12628 10698 -6413 10762
rect -6349 10698 -6329 10762
rect -12628 10682 -6329 10698
rect -12628 10618 -6413 10682
rect -6349 10618 -6329 10682
rect -12628 10602 -6329 10618
rect -12628 10538 -6413 10602
rect -6349 10538 -6329 10602
rect -12628 10522 -6329 10538
rect -12628 10458 -6413 10522
rect -6349 10458 -6329 10522
rect -12628 10442 -6329 10458
rect -12628 10378 -6413 10442
rect -6349 10378 -6329 10442
rect -12628 10362 -6329 10378
rect -12628 10298 -6413 10362
rect -6349 10298 -6329 10362
rect -12628 10282 -6329 10298
rect -12628 10218 -6413 10282
rect -6349 10218 -6329 10282
rect -12628 10202 -6329 10218
rect -12628 10138 -6413 10202
rect -6349 10138 -6329 10202
rect -12628 10122 -6329 10138
rect -12628 10058 -6413 10122
rect -6349 10058 -6329 10122
rect -12628 10042 -6329 10058
rect -12628 9978 -6413 10042
rect -6349 9978 -6329 10042
rect -12628 9962 -6329 9978
rect -12628 9898 -6413 9962
rect -6349 9898 -6329 9962
rect -12628 9882 -6329 9898
rect -12628 9818 -6413 9882
rect -6349 9818 -6329 9882
rect -12628 9802 -6329 9818
rect -12628 9738 -6413 9802
rect -6349 9738 -6329 9802
rect -12628 9722 -6329 9738
rect -12628 9658 -6413 9722
rect -6349 9658 -6329 9722
rect -12628 9642 -6329 9658
rect -12628 9578 -6413 9642
rect -6349 9578 -6329 9642
rect -12628 9562 -6329 9578
rect -12628 9498 -6413 9562
rect -6349 9498 -6329 9562
rect -12628 9482 -6329 9498
rect -12628 9418 -6413 9482
rect -6349 9418 -6329 9482
rect -12628 9402 -6329 9418
rect -12628 9338 -6413 9402
rect -6349 9338 -6329 9402
rect -12628 9322 -6329 9338
rect -12628 9258 -6413 9322
rect -6349 9258 -6329 9322
rect -12628 9242 -6329 9258
rect -12628 9178 -6413 9242
rect -6349 9178 -6329 9242
rect -12628 9162 -6329 9178
rect -12628 9098 -6413 9162
rect -6349 9098 -6329 9162
rect -12628 9082 -6329 9098
rect -12628 9018 -6413 9082
rect -6349 9018 -6329 9082
rect -12628 9002 -6329 9018
rect -12628 8938 -6413 9002
rect -6349 8938 -6329 9002
rect -12628 8922 -6329 8938
rect -12628 8858 -6413 8922
rect -6349 8858 -6329 8922
rect -12628 8842 -6329 8858
rect -12628 8778 -6413 8842
rect -6349 8778 -6329 8842
rect -12628 8762 -6329 8778
rect -12628 8698 -6413 8762
rect -6349 8698 -6329 8762
rect -12628 8682 -6329 8698
rect -12628 8618 -6413 8682
rect -6349 8618 -6329 8682
rect -12628 8602 -6329 8618
rect -12628 8538 -6413 8602
rect -6349 8538 -6329 8602
rect -12628 8522 -6329 8538
rect -12628 8458 -6413 8522
rect -6349 8458 -6329 8522
rect -12628 8442 -6329 8458
rect -12628 8378 -6413 8442
rect -6349 8378 -6329 8442
rect -12628 8362 -6329 8378
rect -12628 8298 -6413 8362
rect -6349 8298 -6329 8362
rect -12628 8282 -6329 8298
rect -12628 8218 -6413 8282
rect -6349 8218 -6329 8282
rect -12628 8202 -6329 8218
rect -12628 8138 -6413 8202
rect -6349 8138 -6329 8202
rect -12628 8122 -6329 8138
rect -12628 8058 -6413 8122
rect -6349 8058 -6329 8122
rect -12628 8042 -6329 8058
rect -12628 7978 -6413 8042
rect -6349 7978 -6329 8042
rect -12628 7962 -6329 7978
rect -12628 7898 -6413 7962
rect -6349 7898 -6329 7962
rect -12628 7882 -6329 7898
rect -12628 7818 -6413 7882
rect -6349 7818 -6329 7882
rect -12628 7802 -6329 7818
rect -12628 7738 -6413 7802
rect -6349 7738 -6329 7802
rect -12628 7722 -6329 7738
rect -12628 7658 -6413 7722
rect -6349 7658 -6329 7722
rect -12628 7642 -6329 7658
rect -12628 7578 -6413 7642
rect -6349 7578 -6329 7642
rect -12628 7562 -6329 7578
rect -12628 7498 -6413 7562
rect -6349 7498 -6329 7562
rect -12628 7482 -6329 7498
rect -12628 7418 -6413 7482
rect -6349 7418 -6329 7482
rect -12628 7402 -6329 7418
rect -12628 7338 -6413 7402
rect -6349 7338 -6329 7402
rect -12628 7322 -6329 7338
rect -12628 7258 -6413 7322
rect -6349 7258 -6329 7322
rect -12628 7242 -6329 7258
rect -12628 7178 -6413 7242
rect -6349 7178 -6329 7242
rect -12628 7162 -6329 7178
rect -12628 7098 -6413 7162
rect -6349 7098 -6329 7162
rect -12628 7082 -6329 7098
rect -12628 7018 -6413 7082
rect -6349 7018 -6329 7082
rect -12628 7002 -6329 7018
rect -12628 6938 -6413 7002
rect -6349 6938 -6329 7002
rect -12628 6922 -6329 6938
rect -12628 6858 -6413 6922
rect -6349 6858 -6329 6922
rect -12628 6842 -6329 6858
rect -12628 6778 -6413 6842
rect -6349 6778 -6329 6842
rect -12628 6762 -6329 6778
rect -12628 6698 -6413 6762
rect -6349 6698 -6329 6762
rect -12628 6682 -6329 6698
rect -12628 6618 -6413 6682
rect -6349 6618 -6329 6682
rect -12628 6602 -6329 6618
rect -12628 6538 -6413 6602
rect -6349 6538 -6329 6602
rect -12628 6522 -6329 6538
rect -12628 6458 -6413 6522
rect -6349 6458 -6329 6522
rect -12628 6442 -6329 6458
rect -12628 6378 -6413 6442
rect -6349 6378 -6329 6442
rect -12628 6350 -6329 6378
rect -6309 12522 -10 12550
rect -6309 12458 -94 12522
rect -30 12458 -10 12522
rect -6309 12442 -10 12458
rect -6309 12378 -94 12442
rect -30 12378 -10 12442
rect -6309 12362 -10 12378
rect -6309 12298 -94 12362
rect -30 12298 -10 12362
rect -6309 12282 -10 12298
rect -6309 12218 -94 12282
rect -30 12218 -10 12282
rect -6309 12202 -10 12218
rect -6309 12138 -94 12202
rect -30 12138 -10 12202
rect -6309 12122 -10 12138
rect -6309 12058 -94 12122
rect -30 12058 -10 12122
rect -6309 12042 -10 12058
rect -6309 11978 -94 12042
rect -30 11978 -10 12042
rect -6309 11962 -10 11978
rect -6309 11898 -94 11962
rect -30 11898 -10 11962
rect -6309 11882 -10 11898
rect -6309 11818 -94 11882
rect -30 11818 -10 11882
rect -6309 11802 -10 11818
rect -6309 11738 -94 11802
rect -30 11738 -10 11802
rect -6309 11722 -10 11738
rect -6309 11658 -94 11722
rect -30 11658 -10 11722
rect -6309 11642 -10 11658
rect -6309 11578 -94 11642
rect -30 11578 -10 11642
rect -6309 11562 -10 11578
rect -6309 11498 -94 11562
rect -30 11498 -10 11562
rect -6309 11482 -10 11498
rect -6309 11418 -94 11482
rect -30 11418 -10 11482
rect -6309 11402 -10 11418
rect -6309 11338 -94 11402
rect -30 11338 -10 11402
rect -6309 11322 -10 11338
rect -6309 11258 -94 11322
rect -30 11258 -10 11322
rect -6309 11242 -10 11258
rect -6309 11178 -94 11242
rect -30 11178 -10 11242
rect -6309 11162 -10 11178
rect -6309 11098 -94 11162
rect -30 11098 -10 11162
rect -6309 11082 -10 11098
rect -6309 11018 -94 11082
rect -30 11018 -10 11082
rect -6309 11002 -10 11018
rect -6309 10938 -94 11002
rect -30 10938 -10 11002
rect -6309 10922 -10 10938
rect -6309 10858 -94 10922
rect -30 10858 -10 10922
rect -6309 10842 -10 10858
rect -6309 10778 -94 10842
rect -30 10778 -10 10842
rect -6309 10762 -10 10778
rect -6309 10698 -94 10762
rect -30 10698 -10 10762
rect -6309 10682 -10 10698
rect -6309 10618 -94 10682
rect -30 10618 -10 10682
rect -6309 10602 -10 10618
rect -6309 10538 -94 10602
rect -30 10538 -10 10602
rect -6309 10522 -10 10538
rect -6309 10458 -94 10522
rect -30 10458 -10 10522
rect -6309 10442 -10 10458
rect -6309 10378 -94 10442
rect -30 10378 -10 10442
rect -6309 10362 -10 10378
rect -6309 10298 -94 10362
rect -30 10298 -10 10362
rect -6309 10282 -10 10298
rect -6309 10218 -94 10282
rect -30 10218 -10 10282
rect -6309 10202 -10 10218
rect -6309 10138 -94 10202
rect -30 10138 -10 10202
rect -6309 10122 -10 10138
rect -6309 10058 -94 10122
rect -30 10058 -10 10122
rect -6309 10042 -10 10058
rect -6309 9978 -94 10042
rect -30 9978 -10 10042
rect -6309 9962 -10 9978
rect -6309 9898 -94 9962
rect -30 9898 -10 9962
rect -6309 9882 -10 9898
rect -6309 9818 -94 9882
rect -30 9818 -10 9882
rect -6309 9802 -10 9818
rect -6309 9738 -94 9802
rect -30 9738 -10 9802
rect -6309 9722 -10 9738
rect -6309 9658 -94 9722
rect -30 9658 -10 9722
rect -6309 9642 -10 9658
rect -6309 9578 -94 9642
rect -30 9578 -10 9642
rect -6309 9562 -10 9578
rect -6309 9498 -94 9562
rect -30 9498 -10 9562
rect -6309 9482 -10 9498
rect -6309 9418 -94 9482
rect -30 9418 -10 9482
rect -6309 9402 -10 9418
rect -6309 9338 -94 9402
rect -30 9338 -10 9402
rect -6309 9322 -10 9338
rect -6309 9258 -94 9322
rect -30 9258 -10 9322
rect -6309 9242 -10 9258
rect -6309 9178 -94 9242
rect -30 9178 -10 9242
rect -6309 9162 -10 9178
rect -6309 9098 -94 9162
rect -30 9098 -10 9162
rect -6309 9082 -10 9098
rect -6309 9018 -94 9082
rect -30 9018 -10 9082
rect -6309 9002 -10 9018
rect -6309 8938 -94 9002
rect -30 8938 -10 9002
rect -6309 8922 -10 8938
rect -6309 8858 -94 8922
rect -30 8858 -10 8922
rect -6309 8842 -10 8858
rect -6309 8778 -94 8842
rect -30 8778 -10 8842
rect -6309 8762 -10 8778
rect -6309 8698 -94 8762
rect -30 8698 -10 8762
rect -6309 8682 -10 8698
rect -6309 8618 -94 8682
rect -30 8618 -10 8682
rect -6309 8602 -10 8618
rect -6309 8538 -94 8602
rect -30 8538 -10 8602
rect -6309 8522 -10 8538
rect -6309 8458 -94 8522
rect -30 8458 -10 8522
rect -6309 8442 -10 8458
rect -6309 8378 -94 8442
rect -30 8378 -10 8442
rect -6309 8362 -10 8378
rect -6309 8298 -94 8362
rect -30 8298 -10 8362
rect -6309 8282 -10 8298
rect -6309 8218 -94 8282
rect -30 8218 -10 8282
rect -6309 8202 -10 8218
rect -6309 8138 -94 8202
rect -30 8138 -10 8202
rect -6309 8122 -10 8138
rect -6309 8058 -94 8122
rect -30 8058 -10 8122
rect -6309 8042 -10 8058
rect -6309 7978 -94 8042
rect -30 7978 -10 8042
rect -6309 7962 -10 7978
rect -6309 7898 -94 7962
rect -30 7898 -10 7962
rect -6309 7882 -10 7898
rect -6309 7818 -94 7882
rect -30 7818 -10 7882
rect -6309 7802 -10 7818
rect -6309 7738 -94 7802
rect -30 7738 -10 7802
rect -6309 7722 -10 7738
rect -6309 7658 -94 7722
rect -30 7658 -10 7722
rect -6309 7642 -10 7658
rect -6309 7578 -94 7642
rect -30 7578 -10 7642
rect -6309 7562 -10 7578
rect -6309 7498 -94 7562
rect -30 7498 -10 7562
rect -6309 7482 -10 7498
rect -6309 7418 -94 7482
rect -30 7418 -10 7482
rect -6309 7402 -10 7418
rect -6309 7338 -94 7402
rect -30 7338 -10 7402
rect -6309 7322 -10 7338
rect -6309 7258 -94 7322
rect -30 7258 -10 7322
rect -6309 7242 -10 7258
rect -6309 7178 -94 7242
rect -30 7178 -10 7242
rect -6309 7162 -10 7178
rect -6309 7098 -94 7162
rect -30 7098 -10 7162
rect -6309 7082 -10 7098
rect -6309 7018 -94 7082
rect -30 7018 -10 7082
rect -6309 7002 -10 7018
rect -6309 6938 -94 7002
rect -30 6938 -10 7002
rect -6309 6922 -10 6938
rect -6309 6858 -94 6922
rect -30 6858 -10 6922
rect -6309 6842 -10 6858
rect -6309 6778 -94 6842
rect -30 6778 -10 6842
rect -6309 6762 -10 6778
rect -6309 6698 -94 6762
rect -30 6698 -10 6762
rect -6309 6682 -10 6698
rect -6309 6618 -94 6682
rect -30 6618 -10 6682
rect -6309 6602 -10 6618
rect -6309 6538 -94 6602
rect -30 6538 -10 6602
rect -6309 6522 -10 6538
rect -6309 6458 -94 6522
rect -30 6458 -10 6522
rect -6309 6442 -10 6458
rect -6309 6378 -94 6442
rect -30 6378 -10 6442
rect -6309 6350 -10 6378
rect 10 12522 6309 12550
rect 10 12458 6225 12522
rect 6289 12458 6309 12522
rect 10 12442 6309 12458
rect 10 12378 6225 12442
rect 6289 12378 6309 12442
rect 10 12362 6309 12378
rect 10 12298 6225 12362
rect 6289 12298 6309 12362
rect 10 12282 6309 12298
rect 10 12218 6225 12282
rect 6289 12218 6309 12282
rect 10 12202 6309 12218
rect 10 12138 6225 12202
rect 6289 12138 6309 12202
rect 10 12122 6309 12138
rect 10 12058 6225 12122
rect 6289 12058 6309 12122
rect 10 12042 6309 12058
rect 10 11978 6225 12042
rect 6289 11978 6309 12042
rect 10 11962 6309 11978
rect 10 11898 6225 11962
rect 6289 11898 6309 11962
rect 10 11882 6309 11898
rect 10 11818 6225 11882
rect 6289 11818 6309 11882
rect 10 11802 6309 11818
rect 10 11738 6225 11802
rect 6289 11738 6309 11802
rect 10 11722 6309 11738
rect 10 11658 6225 11722
rect 6289 11658 6309 11722
rect 10 11642 6309 11658
rect 10 11578 6225 11642
rect 6289 11578 6309 11642
rect 10 11562 6309 11578
rect 10 11498 6225 11562
rect 6289 11498 6309 11562
rect 10 11482 6309 11498
rect 10 11418 6225 11482
rect 6289 11418 6309 11482
rect 10 11402 6309 11418
rect 10 11338 6225 11402
rect 6289 11338 6309 11402
rect 10 11322 6309 11338
rect 10 11258 6225 11322
rect 6289 11258 6309 11322
rect 10 11242 6309 11258
rect 10 11178 6225 11242
rect 6289 11178 6309 11242
rect 10 11162 6309 11178
rect 10 11098 6225 11162
rect 6289 11098 6309 11162
rect 10 11082 6309 11098
rect 10 11018 6225 11082
rect 6289 11018 6309 11082
rect 10 11002 6309 11018
rect 10 10938 6225 11002
rect 6289 10938 6309 11002
rect 10 10922 6309 10938
rect 10 10858 6225 10922
rect 6289 10858 6309 10922
rect 10 10842 6309 10858
rect 10 10778 6225 10842
rect 6289 10778 6309 10842
rect 10 10762 6309 10778
rect 10 10698 6225 10762
rect 6289 10698 6309 10762
rect 10 10682 6309 10698
rect 10 10618 6225 10682
rect 6289 10618 6309 10682
rect 10 10602 6309 10618
rect 10 10538 6225 10602
rect 6289 10538 6309 10602
rect 10 10522 6309 10538
rect 10 10458 6225 10522
rect 6289 10458 6309 10522
rect 10 10442 6309 10458
rect 10 10378 6225 10442
rect 6289 10378 6309 10442
rect 10 10362 6309 10378
rect 10 10298 6225 10362
rect 6289 10298 6309 10362
rect 10 10282 6309 10298
rect 10 10218 6225 10282
rect 6289 10218 6309 10282
rect 10 10202 6309 10218
rect 10 10138 6225 10202
rect 6289 10138 6309 10202
rect 10 10122 6309 10138
rect 10 10058 6225 10122
rect 6289 10058 6309 10122
rect 10 10042 6309 10058
rect 10 9978 6225 10042
rect 6289 9978 6309 10042
rect 10 9962 6309 9978
rect 10 9898 6225 9962
rect 6289 9898 6309 9962
rect 10 9882 6309 9898
rect 10 9818 6225 9882
rect 6289 9818 6309 9882
rect 10 9802 6309 9818
rect 10 9738 6225 9802
rect 6289 9738 6309 9802
rect 10 9722 6309 9738
rect 10 9658 6225 9722
rect 6289 9658 6309 9722
rect 10 9642 6309 9658
rect 10 9578 6225 9642
rect 6289 9578 6309 9642
rect 10 9562 6309 9578
rect 10 9498 6225 9562
rect 6289 9498 6309 9562
rect 10 9482 6309 9498
rect 10 9418 6225 9482
rect 6289 9418 6309 9482
rect 10 9402 6309 9418
rect 10 9338 6225 9402
rect 6289 9338 6309 9402
rect 10 9322 6309 9338
rect 10 9258 6225 9322
rect 6289 9258 6309 9322
rect 10 9242 6309 9258
rect 10 9178 6225 9242
rect 6289 9178 6309 9242
rect 10 9162 6309 9178
rect 10 9098 6225 9162
rect 6289 9098 6309 9162
rect 10 9082 6309 9098
rect 10 9018 6225 9082
rect 6289 9018 6309 9082
rect 10 9002 6309 9018
rect 10 8938 6225 9002
rect 6289 8938 6309 9002
rect 10 8922 6309 8938
rect 10 8858 6225 8922
rect 6289 8858 6309 8922
rect 10 8842 6309 8858
rect 10 8778 6225 8842
rect 6289 8778 6309 8842
rect 10 8762 6309 8778
rect 10 8698 6225 8762
rect 6289 8698 6309 8762
rect 10 8682 6309 8698
rect 10 8618 6225 8682
rect 6289 8618 6309 8682
rect 10 8602 6309 8618
rect 10 8538 6225 8602
rect 6289 8538 6309 8602
rect 10 8522 6309 8538
rect 10 8458 6225 8522
rect 6289 8458 6309 8522
rect 10 8442 6309 8458
rect 10 8378 6225 8442
rect 6289 8378 6309 8442
rect 10 8362 6309 8378
rect 10 8298 6225 8362
rect 6289 8298 6309 8362
rect 10 8282 6309 8298
rect 10 8218 6225 8282
rect 6289 8218 6309 8282
rect 10 8202 6309 8218
rect 10 8138 6225 8202
rect 6289 8138 6309 8202
rect 10 8122 6309 8138
rect 10 8058 6225 8122
rect 6289 8058 6309 8122
rect 10 8042 6309 8058
rect 10 7978 6225 8042
rect 6289 7978 6309 8042
rect 10 7962 6309 7978
rect 10 7898 6225 7962
rect 6289 7898 6309 7962
rect 10 7882 6309 7898
rect 10 7818 6225 7882
rect 6289 7818 6309 7882
rect 10 7802 6309 7818
rect 10 7738 6225 7802
rect 6289 7738 6309 7802
rect 10 7722 6309 7738
rect 10 7658 6225 7722
rect 6289 7658 6309 7722
rect 10 7642 6309 7658
rect 10 7578 6225 7642
rect 6289 7578 6309 7642
rect 10 7562 6309 7578
rect 10 7498 6225 7562
rect 6289 7498 6309 7562
rect 10 7482 6309 7498
rect 10 7418 6225 7482
rect 6289 7418 6309 7482
rect 10 7402 6309 7418
rect 10 7338 6225 7402
rect 6289 7338 6309 7402
rect 10 7322 6309 7338
rect 10 7258 6225 7322
rect 6289 7258 6309 7322
rect 10 7242 6309 7258
rect 10 7178 6225 7242
rect 6289 7178 6309 7242
rect 10 7162 6309 7178
rect 10 7098 6225 7162
rect 6289 7098 6309 7162
rect 10 7082 6309 7098
rect 10 7018 6225 7082
rect 6289 7018 6309 7082
rect 10 7002 6309 7018
rect 10 6938 6225 7002
rect 6289 6938 6309 7002
rect 10 6922 6309 6938
rect 10 6858 6225 6922
rect 6289 6858 6309 6922
rect 10 6842 6309 6858
rect 10 6778 6225 6842
rect 6289 6778 6309 6842
rect 10 6762 6309 6778
rect 10 6698 6225 6762
rect 6289 6698 6309 6762
rect 10 6682 6309 6698
rect 10 6618 6225 6682
rect 6289 6618 6309 6682
rect 10 6602 6309 6618
rect 10 6538 6225 6602
rect 6289 6538 6309 6602
rect 10 6522 6309 6538
rect 10 6458 6225 6522
rect 6289 6458 6309 6522
rect 10 6442 6309 6458
rect 10 6378 6225 6442
rect 6289 6378 6309 6442
rect 10 6350 6309 6378
rect 6329 12522 12628 12550
rect 6329 12458 12544 12522
rect 12608 12458 12628 12522
rect 6329 12442 12628 12458
rect 6329 12378 12544 12442
rect 12608 12378 12628 12442
rect 6329 12362 12628 12378
rect 6329 12298 12544 12362
rect 12608 12298 12628 12362
rect 6329 12282 12628 12298
rect 6329 12218 12544 12282
rect 12608 12218 12628 12282
rect 6329 12202 12628 12218
rect 6329 12138 12544 12202
rect 12608 12138 12628 12202
rect 6329 12122 12628 12138
rect 6329 12058 12544 12122
rect 12608 12058 12628 12122
rect 6329 12042 12628 12058
rect 6329 11978 12544 12042
rect 12608 11978 12628 12042
rect 6329 11962 12628 11978
rect 6329 11898 12544 11962
rect 12608 11898 12628 11962
rect 6329 11882 12628 11898
rect 6329 11818 12544 11882
rect 12608 11818 12628 11882
rect 6329 11802 12628 11818
rect 6329 11738 12544 11802
rect 12608 11738 12628 11802
rect 6329 11722 12628 11738
rect 6329 11658 12544 11722
rect 12608 11658 12628 11722
rect 6329 11642 12628 11658
rect 6329 11578 12544 11642
rect 12608 11578 12628 11642
rect 6329 11562 12628 11578
rect 6329 11498 12544 11562
rect 12608 11498 12628 11562
rect 6329 11482 12628 11498
rect 6329 11418 12544 11482
rect 12608 11418 12628 11482
rect 6329 11402 12628 11418
rect 6329 11338 12544 11402
rect 12608 11338 12628 11402
rect 6329 11322 12628 11338
rect 6329 11258 12544 11322
rect 12608 11258 12628 11322
rect 6329 11242 12628 11258
rect 6329 11178 12544 11242
rect 12608 11178 12628 11242
rect 6329 11162 12628 11178
rect 6329 11098 12544 11162
rect 12608 11098 12628 11162
rect 6329 11082 12628 11098
rect 6329 11018 12544 11082
rect 12608 11018 12628 11082
rect 6329 11002 12628 11018
rect 6329 10938 12544 11002
rect 12608 10938 12628 11002
rect 6329 10922 12628 10938
rect 6329 10858 12544 10922
rect 12608 10858 12628 10922
rect 6329 10842 12628 10858
rect 6329 10778 12544 10842
rect 12608 10778 12628 10842
rect 6329 10762 12628 10778
rect 6329 10698 12544 10762
rect 12608 10698 12628 10762
rect 6329 10682 12628 10698
rect 6329 10618 12544 10682
rect 12608 10618 12628 10682
rect 6329 10602 12628 10618
rect 6329 10538 12544 10602
rect 12608 10538 12628 10602
rect 6329 10522 12628 10538
rect 6329 10458 12544 10522
rect 12608 10458 12628 10522
rect 6329 10442 12628 10458
rect 6329 10378 12544 10442
rect 12608 10378 12628 10442
rect 6329 10362 12628 10378
rect 6329 10298 12544 10362
rect 12608 10298 12628 10362
rect 6329 10282 12628 10298
rect 6329 10218 12544 10282
rect 12608 10218 12628 10282
rect 6329 10202 12628 10218
rect 6329 10138 12544 10202
rect 12608 10138 12628 10202
rect 6329 10122 12628 10138
rect 6329 10058 12544 10122
rect 12608 10058 12628 10122
rect 6329 10042 12628 10058
rect 6329 9978 12544 10042
rect 12608 9978 12628 10042
rect 6329 9962 12628 9978
rect 6329 9898 12544 9962
rect 12608 9898 12628 9962
rect 6329 9882 12628 9898
rect 6329 9818 12544 9882
rect 12608 9818 12628 9882
rect 6329 9802 12628 9818
rect 6329 9738 12544 9802
rect 12608 9738 12628 9802
rect 6329 9722 12628 9738
rect 6329 9658 12544 9722
rect 12608 9658 12628 9722
rect 6329 9642 12628 9658
rect 6329 9578 12544 9642
rect 12608 9578 12628 9642
rect 6329 9562 12628 9578
rect 6329 9498 12544 9562
rect 12608 9498 12628 9562
rect 6329 9482 12628 9498
rect 6329 9418 12544 9482
rect 12608 9418 12628 9482
rect 6329 9402 12628 9418
rect 6329 9338 12544 9402
rect 12608 9338 12628 9402
rect 6329 9322 12628 9338
rect 6329 9258 12544 9322
rect 12608 9258 12628 9322
rect 6329 9242 12628 9258
rect 6329 9178 12544 9242
rect 12608 9178 12628 9242
rect 6329 9162 12628 9178
rect 6329 9098 12544 9162
rect 12608 9098 12628 9162
rect 6329 9082 12628 9098
rect 6329 9018 12544 9082
rect 12608 9018 12628 9082
rect 6329 9002 12628 9018
rect 6329 8938 12544 9002
rect 12608 8938 12628 9002
rect 6329 8922 12628 8938
rect 6329 8858 12544 8922
rect 12608 8858 12628 8922
rect 6329 8842 12628 8858
rect 6329 8778 12544 8842
rect 12608 8778 12628 8842
rect 6329 8762 12628 8778
rect 6329 8698 12544 8762
rect 12608 8698 12628 8762
rect 6329 8682 12628 8698
rect 6329 8618 12544 8682
rect 12608 8618 12628 8682
rect 6329 8602 12628 8618
rect 6329 8538 12544 8602
rect 12608 8538 12628 8602
rect 6329 8522 12628 8538
rect 6329 8458 12544 8522
rect 12608 8458 12628 8522
rect 6329 8442 12628 8458
rect 6329 8378 12544 8442
rect 12608 8378 12628 8442
rect 6329 8362 12628 8378
rect 6329 8298 12544 8362
rect 12608 8298 12628 8362
rect 6329 8282 12628 8298
rect 6329 8218 12544 8282
rect 12608 8218 12628 8282
rect 6329 8202 12628 8218
rect 6329 8138 12544 8202
rect 12608 8138 12628 8202
rect 6329 8122 12628 8138
rect 6329 8058 12544 8122
rect 12608 8058 12628 8122
rect 6329 8042 12628 8058
rect 6329 7978 12544 8042
rect 12608 7978 12628 8042
rect 6329 7962 12628 7978
rect 6329 7898 12544 7962
rect 12608 7898 12628 7962
rect 6329 7882 12628 7898
rect 6329 7818 12544 7882
rect 12608 7818 12628 7882
rect 6329 7802 12628 7818
rect 6329 7738 12544 7802
rect 12608 7738 12628 7802
rect 6329 7722 12628 7738
rect 6329 7658 12544 7722
rect 12608 7658 12628 7722
rect 6329 7642 12628 7658
rect 6329 7578 12544 7642
rect 12608 7578 12628 7642
rect 6329 7562 12628 7578
rect 6329 7498 12544 7562
rect 12608 7498 12628 7562
rect 6329 7482 12628 7498
rect 6329 7418 12544 7482
rect 12608 7418 12628 7482
rect 6329 7402 12628 7418
rect 6329 7338 12544 7402
rect 12608 7338 12628 7402
rect 6329 7322 12628 7338
rect 6329 7258 12544 7322
rect 12608 7258 12628 7322
rect 6329 7242 12628 7258
rect 6329 7178 12544 7242
rect 12608 7178 12628 7242
rect 6329 7162 12628 7178
rect 6329 7098 12544 7162
rect 12608 7098 12628 7162
rect 6329 7082 12628 7098
rect 6329 7018 12544 7082
rect 12608 7018 12628 7082
rect 6329 7002 12628 7018
rect 6329 6938 12544 7002
rect 12608 6938 12628 7002
rect 6329 6922 12628 6938
rect 6329 6858 12544 6922
rect 12608 6858 12628 6922
rect 6329 6842 12628 6858
rect 6329 6778 12544 6842
rect 12608 6778 12628 6842
rect 6329 6762 12628 6778
rect 6329 6698 12544 6762
rect 12608 6698 12628 6762
rect 6329 6682 12628 6698
rect 6329 6618 12544 6682
rect 12608 6618 12628 6682
rect 6329 6602 12628 6618
rect 6329 6538 12544 6602
rect 12608 6538 12628 6602
rect 6329 6522 12628 6538
rect 6329 6458 12544 6522
rect 12608 6458 12628 6522
rect 6329 6442 12628 6458
rect 6329 6378 12544 6442
rect 12608 6378 12628 6442
rect 6329 6350 12628 6378
rect -12628 6222 -6329 6250
rect -12628 6158 -6413 6222
rect -6349 6158 -6329 6222
rect -12628 6142 -6329 6158
rect -12628 6078 -6413 6142
rect -6349 6078 -6329 6142
rect -12628 6062 -6329 6078
rect -12628 5998 -6413 6062
rect -6349 5998 -6329 6062
rect -12628 5982 -6329 5998
rect -12628 5918 -6413 5982
rect -6349 5918 -6329 5982
rect -12628 5902 -6329 5918
rect -12628 5838 -6413 5902
rect -6349 5838 -6329 5902
rect -12628 5822 -6329 5838
rect -12628 5758 -6413 5822
rect -6349 5758 -6329 5822
rect -12628 5742 -6329 5758
rect -12628 5678 -6413 5742
rect -6349 5678 -6329 5742
rect -12628 5662 -6329 5678
rect -12628 5598 -6413 5662
rect -6349 5598 -6329 5662
rect -12628 5582 -6329 5598
rect -12628 5518 -6413 5582
rect -6349 5518 -6329 5582
rect -12628 5502 -6329 5518
rect -12628 5438 -6413 5502
rect -6349 5438 -6329 5502
rect -12628 5422 -6329 5438
rect -12628 5358 -6413 5422
rect -6349 5358 -6329 5422
rect -12628 5342 -6329 5358
rect -12628 5278 -6413 5342
rect -6349 5278 -6329 5342
rect -12628 5262 -6329 5278
rect -12628 5198 -6413 5262
rect -6349 5198 -6329 5262
rect -12628 5182 -6329 5198
rect -12628 5118 -6413 5182
rect -6349 5118 -6329 5182
rect -12628 5102 -6329 5118
rect -12628 5038 -6413 5102
rect -6349 5038 -6329 5102
rect -12628 5022 -6329 5038
rect -12628 4958 -6413 5022
rect -6349 4958 -6329 5022
rect -12628 4942 -6329 4958
rect -12628 4878 -6413 4942
rect -6349 4878 -6329 4942
rect -12628 4862 -6329 4878
rect -12628 4798 -6413 4862
rect -6349 4798 -6329 4862
rect -12628 4782 -6329 4798
rect -12628 4718 -6413 4782
rect -6349 4718 -6329 4782
rect -12628 4702 -6329 4718
rect -12628 4638 -6413 4702
rect -6349 4638 -6329 4702
rect -12628 4622 -6329 4638
rect -12628 4558 -6413 4622
rect -6349 4558 -6329 4622
rect -12628 4542 -6329 4558
rect -12628 4478 -6413 4542
rect -6349 4478 -6329 4542
rect -12628 4462 -6329 4478
rect -12628 4398 -6413 4462
rect -6349 4398 -6329 4462
rect -12628 4382 -6329 4398
rect -12628 4318 -6413 4382
rect -6349 4318 -6329 4382
rect -12628 4302 -6329 4318
rect -12628 4238 -6413 4302
rect -6349 4238 -6329 4302
rect -12628 4222 -6329 4238
rect -12628 4158 -6413 4222
rect -6349 4158 -6329 4222
rect -12628 4142 -6329 4158
rect -12628 4078 -6413 4142
rect -6349 4078 -6329 4142
rect -12628 4062 -6329 4078
rect -12628 3998 -6413 4062
rect -6349 3998 -6329 4062
rect -12628 3982 -6329 3998
rect -12628 3918 -6413 3982
rect -6349 3918 -6329 3982
rect -12628 3902 -6329 3918
rect -12628 3838 -6413 3902
rect -6349 3838 -6329 3902
rect -12628 3822 -6329 3838
rect -12628 3758 -6413 3822
rect -6349 3758 -6329 3822
rect -12628 3742 -6329 3758
rect -12628 3678 -6413 3742
rect -6349 3678 -6329 3742
rect -12628 3662 -6329 3678
rect -12628 3598 -6413 3662
rect -6349 3598 -6329 3662
rect -12628 3582 -6329 3598
rect -12628 3518 -6413 3582
rect -6349 3518 -6329 3582
rect -12628 3502 -6329 3518
rect -12628 3438 -6413 3502
rect -6349 3438 -6329 3502
rect -12628 3422 -6329 3438
rect -12628 3358 -6413 3422
rect -6349 3358 -6329 3422
rect -12628 3342 -6329 3358
rect -12628 3278 -6413 3342
rect -6349 3278 -6329 3342
rect -12628 3262 -6329 3278
rect -12628 3198 -6413 3262
rect -6349 3198 -6329 3262
rect -12628 3182 -6329 3198
rect -12628 3118 -6413 3182
rect -6349 3118 -6329 3182
rect -12628 3102 -6329 3118
rect -12628 3038 -6413 3102
rect -6349 3038 -6329 3102
rect -12628 3022 -6329 3038
rect -12628 2958 -6413 3022
rect -6349 2958 -6329 3022
rect -12628 2942 -6329 2958
rect -12628 2878 -6413 2942
rect -6349 2878 -6329 2942
rect -12628 2862 -6329 2878
rect -12628 2798 -6413 2862
rect -6349 2798 -6329 2862
rect -12628 2782 -6329 2798
rect -12628 2718 -6413 2782
rect -6349 2718 -6329 2782
rect -12628 2702 -6329 2718
rect -12628 2638 -6413 2702
rect -6349 2638 -6329 2702
rect -12628 2622 -6329 2638
rect -12628 2558 -6413 2622
rect -6349 2558 -6329 2622
rect -12628 2542 -6329 2558
rect -12628 2478 -6413 2542
rect -6349 2478 -6329 2542
rect -12628 2462 -6329 2478
rect -12628 2398 -6413 2462
rect -6349 2398 -6329 2462
rect -12628 2382 -6329 2398
rect -12628 2318 -6413 2382
rect -6349 2318 -6329 2382
rect -12628 2302 -6329 2318
rect -12628 2238 -6413 2302
rect -6349 2238 -6329 2302
rect -12628 2222 -6329 2238
rect -12628 2158 -6413 2222
rect -6349 2158 -6329 2222
rect -12628 2142 -6329 2158
rect -12628 2078 -6413 2142
rect -6349 2078 -6329 2142
rect -12628 2062 -6329 2078
rect -12628 1998 -6413 2062
rect -6349 1998 -6329 2062
rect -12628 1982 -6329 1998
rect -12628 1918 -6413 1982
rect -6349 1918 -6329 1982
rect -12628 1902 -6329 1918
rect -12628 1838 -6413 1902
rect -6349 1838 -6329 1902
rect -12628 1822 -6329 1838
rect -12628 1758 -6413 1822
rect -6349 1758 -6329 1822
rect -12628 1742 -6329 1758
rect -12628 1678 -6413 1742
rect -6349 1678 -6329 1742
rect -12628 1662 -6329 1678
rect -12628 1598 -6413 1662
rect -6349 1598 -6329 1662
rect -12628 1582 -6329 1598
rect -12628 1518 -6413 1582
rect -6349 1518 -6329 1582
rect -12628 1502 -6329 1518
rect -12628 1438 -6413 1502
rect -6349 1438 -6329 1502
rect -12628 1422 -6329 1438
rect -12628 1358 -6413 1422
rect -6349 1358 -6329 1422
rect -12628 1342 -6329 1358
rect -12628 1278 -6413 1342
rect -6349 1278 -6329 1342
rect -12628 1262 -6329 1278
rect -12628 1198 -6413 1262
rect -6349 1198 -6329 1262
rect -12628 1182 -6329 1198
rect -12628 1118 -6413 1182
rect -6349 1118 -6329 1182
rect -12628 1102 -6329 1118
rect -12628 1038 -6413 1102
rect -6349 1038 -6329 1102
rect -12628 1022 -6329 1038
rect -12628 958 -6413 1022
rect -6349 958 -6329 1022
rect -12628 942 -6329 958
rect -12628 878 -6413 942
rect -6349 878 -6329 942
rect -12628 862 -6329 878
rect -12628 798 -6413 862
rect -6349 798 -6329 862
rect -12628 782 -6329 798
rect -12628 718 -6413 782
rect -6349 718 -6329 782
rect -12628 702 -6329 718
rect -12628 638 -6413 702
rect -6349 638 -6329 702
rect -12628 622 -6329 638
rect -12628 558 -6413 622
rect -6349 558 -6329 622
rect -12628 542 -6329 558
rect -12628 478 -6413 542
rect -6349 478 -6329 542
rect -12628 462 -6329 478
rect -12628 398 -6413 462
rect -6349 398 -6329 462
rect -12628 382 -6329 398
rect -12628 318 -6413 382
rect -6349 318 -6329 382
rect -12628 302 -6329 318
rect -12628 238 -6413 302
rect -6349 238 -6329 302
rect -12628 222 -6329 238
rect -12628 158 -6413 222
rect -6349 158 -6329 222
rect -12628 142 -6329 158
rect -12628 78 -6413 142
rect -6349 78 -6329 142
rect -12628 50 -6329 78
rect -6309 6222 -10 6250
rect -6309 6158 -94 6222
rect -30 6158 -10 6222
rect -6309 6142 -10 6158
rect -6309 6078 -94 6142
rect -30 6078 -10 6142
rect -6309 6062 -10 6078
rect -6309 5998 -94 6062
rect -30 5998 -10 6062
rect -6309 5982 -10 5998
rect -6309 5918 -94 5982
rect -30 5918 -10 5982
rect -6309 5902 -10 5918
rect -6309 5838 -94 5902
rect -30 5838 -10 5902
rect -6309 5822 -10 5838
rect -6309 5758 -94 5822
rect -30 5758 -10 5822
rect -6309 5742 -10 5758
rect -6309 5678 -94 5742
rect -30 5678 -10 5742
rect -6309 5662 -10 5678
rect -6309 5598 -94 5662
rect -30 5598 -10 5662
rect -6309 5582 -10 5598
rect -6309 5518 -94 5582
rect -30 5518 -10 5582
rect -6309 5502 -10 5518
rect -6309 5438 -94 5502
rect -30 5438 -10 5502
rect -6309 5422 -10 5438
rect -6309 5358 -94 5422
rect -30 5358 -10 5422
rect -6309 5342 -10 5358
rect -6309 5278 -94 5342
rect -30 5278 -10 5342
rect -6309 5262 -10 5278
rect -6309 5198 -94 5262
rect -30 5198 -10 5262
rect -6309 5182 -10 5198
rect -6309 5118 -94 5182
rect -30 5118 -10 5182
rect -6309 5102 -10 5118
rect -6309 5038 -94 5102
rect -30 5038 -10 5102
rect -6309 5022 -10 5038
rect -6309 4958 -94 5022
rect -30 4958 -10 5022
rect -6309 4942 -10 4958
rect -6309 4878 -94 4942
rect -30 4878 -10 4942
rect -6309 4862 -10 4878
rect -6309 4798 -94 4862
rect -30 4798 -10 4862
rect -6309 4782 -10 4798
rect -6309 4718 -94 4782
rect -30 4718 -10 4782
rect -6309 4702 -10 4718
rect -6309 4638 -94 4702
rect -30 4638 -10 4702
rect -6309 4622 -10 4638
rect -6309 4558 -94 4622
rect -30 4558 -10 4622
rect -6309 4542 -10 4558
rect -6309 4478 -94 4542
rect -30 4478 -10 4542
rect -6309 4462 -10 4478
rect -6309 4398 -94 4462
rect -30 4398 -10 4462
rect -6309 4382 -10 4398
rect -6309 4318 -94 4382
rect -30 4318 -10 4382
rect -6309 4302 -10 4318
rect -6309 4238 -94 4302
rect -30 4238 -10 4302
rect -6309 4222 -10 4238
rect -6309 4158 -94 4222
rect -30 4158 -10 4222
rect -6309 4142 -10 4158
rect -6309 4078 -94 4142
rect -30 4078 -10 4142
rect -6309 4062 -10 4078
rect -6309 3998 -94 4062
rect -30 3998 -10 4062
rect -6309 3982 -10 3998
rect -6309 3918 -94 3982
rect -30 3918 -10 3982
rect -6309 3902 -10 3918
rect -6309 3838 -94 3902
rect -30 3838 -10 3902
rect -6309 3822 -10 3838
rect -6309 3758 -94 3822
rect -30 3758 -10 3822
rect -6309 3742 -10 3758
rect -6309 3678 -94 3742
rect -30 3678 -10 3742
rect -6309 3662 -10 3678
rect -6309 3598 -94 3662
rect -30 3598 -10 3662
rect -6309 3582 -10 3598
rect -6309 3518 -94 3582
rect -30 3518 -10 3582
rect -6309 3502 -10 3518
rect -6309 3438 -94 3502
rect -30 3438 -10 3502
rect -6309 3422 -10 3438
rect -6309 3358 -94 3422
rect -30 3358 -10 3422
rect -6309 3342 -10 3358
rect -6309 3278 -94 3342
rect -30 3278 -10 3342
rect -6309 3262 -10 3278
rect -6309 3198 -94 3262
rect -30 3198 -10 3262
rect -6309 3182 -10 3198
rect -6309 3118 -94 3182
rect -30 3118 -10 3182
rect -6309 3102 -10 3118
rect -6309 3038 -94 3102
rect -30 3038 -10 3102
rect -6309 3022 -10 3038
rect -6309 2958 -94 3022
rect -30 2958 -10 3022
rect -6309 2942 -10 2958
rect -6309 2878 -94 2942
rect -30 2878 -10 2942
rect -6309 2862 -10 2878
rect -6309 2798 -94 2862
rect -30 2798 -10 2862
rect -6309 2782 -10 2798
rect -6309 2718 -94 2782
rect -30 2718 -10 2782
rect -6309 2702 -10 2718
rect -6309 2638 -94 2702
rect -30 2638 -10 2702
rect -6309 2622 -10 2638
rect -6309 2558 -94 2622
rect -30 2558 -10 2622
rect -6309 2542 -10 2558
rect -6309 2478 -94 2542
rect -30 2478 -10 2542
rect -6309 2462 -10 2478
rect -6309 2398 -94 2462
rect -30 2398 -10 2462
rect -6309 2382 -10 2398
rect -6309 2318 -94 2382
rect -30 2318 -10 2382
rect -6309 2302 -10 2318
rect -6309 2238 -94 2302
rect -30 2238 -10 2302
rect -6309 2222 -10 2238
rect -6309 2158 -94 2222
rect -30 2158 -10 2222
rect -6309 2142 -10 2158
rect -6309 2078 -94 2142
rect -30 2078 -10 2142
rect -6309 2062 -10 2078
rect -6309 1998 -94 2062
rect -30 1998 -10 2062
rect -6309 1982 -10 1998
rect -6309 1918 -94 1982
rect -30 1918 -10 1982
rect -6309 1902 -10 1918
rect -6309 1838 -94 1902
rect -30 1838 -10 1902
rect -6309 1822 -10 1838
rect -6309 1758 -94 1822
rect -30 1758 -10 1822
rect -6309 1742 -10 1758
rect -6309 1678 -94 1742
rect -30 1678 -10 1742
rect -6309 1662 -10 1678
rect -6309 1598 -94 1662
rect -30 1598 -10 1662
rect -6309 1582 -10 1598
rect -6309 1518 -94 1582
rect -30 1518 -10 1582
rect -6309 1502 -10 1518
rect -6309 1438 -94 1502
rect -30 1438 -10 1502
rect -6309 1422 -10 1438
rect -6309 1358 -94 1422
rect -30 1358 -10 1422
rect -6309 1342 -10 1358
rect -6309 1278 -94 1342
rect -30 1278 -10 1342
rect -6309 1262 -10 1278
rect -6309 1198 -94 1262
rect -30 1198 -10 1262
rect -6309 1182 -10 1198
rect -6309 1118 -94 1182
rect -30 1118 -10 1182
rect -6309 1102 -10 1118
rect -6309 1038 -94 1102
rect -30 1038 -10 1102
rect -6309 1022 -10 1038
rect -6309 958 -94 1022
rect -30 958 -10 1022
rect -6309 942 -10 958
rect -6309 878 -94 942
rect -30 878 -10 942
rect -6309 862 -10 878
rect -6309 798 -94 862
rect -30 798 -10 862
rect -6309 782 -10 798
rect -6309 718 -94 782
rect -30 718 -10 782
rect -6309 702 -10 718
rect -6309 638 -94 702
rect -30 638 -10 702
rect -6309 622 -10 638
rect -6309 558 -94 622
rect -30 558 -10 622
rect -6309 542 -10 558
rect -6309 478 -94 542
rect -30 478 -10 542
rect -6309 462 -10 478
rect -6309 398 -94 462
rect -30 398 -10 462
rect -6309 382 -10 398
rect -6309 318 -94 382
rect -30 318 -10 382
rect -6309 302 -10 318
rect -6309 238 -94 302
rect -30 238 -10 302
rect -6309 222 -10 238
rect -6309 158 -94 222
rect -30 158 -10 222
rect -6309 142 -10 158
rect -6309 78 -94 142
rect -30 78 -10 142
rect -6309 50 -10 78
rect 10 6222 6309 6250
rect 10 6158 6225 6222
rect 6289 6158 6309 6222
rect 10 6142 6309 6158
rect 10 6078 6225 6142
rect 6289 6078 6309 6142
rect 10 6062 6309 6078
rect 10 5998 6225 6062
rect 6289 5998 6309 6062
rect 10 5982 6309 5998
rect 10 5918 6225 5982
rect 6289 5918 6309 5982
rect 10 5902 6309 5918
rect 10 5838 6225 5902
rect 6289 5838 6309 5902
rect 10 5822 6309 5838
rect 10 5758 6225 5822
rect 6289 5758 6309 5822
rect 10 5742 6309 5758
rect 10 5678 6225 5742
rect 6289 5678 6309 5742
rect 10 5662 6309 5678
rect 10 5598 6225 5662
rect 6289 5598 6309 5662
rect 10 5582 6309 5598
rect 10 5518 6225 5582
rect 6289 5518 6309 5582
rect 10 5502 6309 5518
rect 10 5438 6225 5502
rect 6289 5438 6309 5502
rect 10 5422 6309 5438
rect 10 5358 6225 5422
rect 6289 5358 6309 5422
rect 10 5342 6309 5358
rect 10 5278 6225 5342
rect 6289 5278 6309 5342
rect 10 5262 6309 5278
rect 10 5198 6225 5262
rect 6289 5198 6309 5262
rect 10 5182 6309 5198
rect 10 5118 6225 5182
rect 6289 5118 6309 5182
rect 10 5102 6309 5118
rect 10 5038 6225 5102
rect 6289 5038 6309 5102
rect 10 5022 6309 5038
rect 10 4958 6225 5022
rect 6289 4958 6309 5022
rect 10 4942 6309 4958
rect 10 4878 6225 4942
rect 6289 4878 6309 4942
rect 10 4862 6309 4878
rect 10 4798 6225 4862
rect 6289 4798 6309 4862
rect 10 4782 6309 4798
rect 10 4718 6225 4782
rect 6289 4718 6309 4782
rect 10 4702 6309 4718
rect 10 4638 6225 4702
rect 6289 4638 6309 4702
rect 10 4622 6309 4638
rect 10 4558 6225 4622
rect 6289 4558 6309 4622
rect 10 4542 6309 4558
rect 10 4478 6225 4542
rect 6289 4478 6309 4542
rect 10 4462 6309 4478
rect 10 4398 6225 4462
rect 6289 4398 6309 4462
rect 10 4382 6309 4398
rect 10 4318 6225 4382
rect 6289 4318 6309 4382
rect 10 4302 6309 4318
rect 10 4238 6225 4302
rect 6289 4238 6309 4302
rect 10 4222 6309 4238
rect 10 4158 6225 4222
rect 6289 4158 6309 4222
rect 10 4142 6309 4158
rect 10 4078 6225 4142
rect 6289 4078 6309 4142
rect 10 4062 6309 4078
rect 10 3998 6225 4062
rect 6289 3998 6309 4062
rect 10 3982 6309 3998
rect 10 3918 6225 3982
rect 6289 3918 6309 3982
rect 10 3902 6309 3918
rect 10 3838 6225 3902
rect 6289 3838 6309 3902
rect 10 3822 6309 3838
rect 10 3758 6225 3822
rect 6289 3758 6309 3822
rect 10 3742 6309 3758
rect 10 3678 6225 3742
rect 6289 3678 6309 3742
rect 10 3662 6309 3678
rect 10 3598 6225 3662
rect 6289 3598 6309 3662
rect 10 3582 6309 3598
rect 10 3518 6225 3582
rect 6289 3518 6309 3582
rect 10 3502 6309 3518
rect 10 3438 6225 3502
rect 6289 3438 6309 3502
rect 10 3422 6309 3438
rect 10 3358 6225 3422
rect 6289 3358 6309 3422
rect 10 3342 6309 3358
rect 10 3278 6225 3342
rect 6289 3278 6309 3342
rect 10 3262 6309 3278
rect 10 3198 6225 3262
rect 6289 3198 6309 3262
rect 10 3182 6309 3198
rect 10 3118 6225 3182
rect 6289 3118 6309 3182
rect 10 3102 6309 3118
rect 10 3038 6225 3102
rect 6289 3038 6309 3102
rect 10 3022 6309 3038
rect 10 2958 6225 3022
rect 6289 2958 6309 3022
rect 10 2942 6309 2958
rect 10 2878 6225 2942
rect 6289 2878 6309 2942
rect 10 2862 6309 2878
rect 10 2798 6225 2862
rect 6289 2798 6309 2862
rect 10 2782 6309 2798
rect 10 2718 6225 2782
rect 6289 2718 6309 2782
rect 10 2702 6309 2718
rect 10 2638 6225 2702
rect 6289 2638 6309 2702
rect 10 2622 6309 2638
rect 10 2558 6225 2622
rect 6289 2558 6309 2622
rect 10 2542 6309 2558
rect 10 2478 6225 2542
rect 6289 2478 6309 2542
rect 10 2462 6309 2478
rect 10 2398 6225 2462
rect 6289 2398 6309 2462
rect 10 2382 6309 2398
rect 10 2318 6225 2382
rect 6289 2318 6309 2382
rect 10 2302 6309 2318
rect 10 2238 6225 2302
rect 6289 2238 6309 2302
rect 10 2222 6309 2238
rect 10 2158 6225 2222
rect 6289 2158 6309 2222
rect 10 2142 6309 2158
rect 10 2078 6225 2142
rect 6289 2078 6309 2142
rect 10 2062 6309 2078
rect 10 1998 6225 2062
rect 6289 1998 6309 2062
rect 10 1982 6309 1998
rect 10 1918 6225 1982
rect 6289 1918 6309 1982
rect 10 1902 6309 1918
rect 10 1838 6225 1902
rect 6289 1838 6309 1902
rect 10 1822 6309 1838
rect 10 1758 6225 1822
rect 6289 1758 6309 1822
rect 10 1742 6309 1758
rect 10 1678 6225 1742
rect 6289 1678 6309 1742
rect 10 1662 6309 1678
rect 10 1598 6225 1662
rect 6289 1598 6309 1662
rect 10 1582 6309 1598
rect 10 1518 6225 1582
rect 6289 1518 6309 1582
rect 10 1502 6309 1518
rect 10 1438 6225 1502
rect 6289 1438 6309 1502
rect 10 1422 6309 1438
rect 10 1358 6225 1422
rect 6289 1358 6309 1422
rect 10 1342 6309 1358
rect 10 1278 6225 1342
rect 6289 1278 6309 1342
rect 10 1262 6309 1278
rect 10 1198 6225 1262
rect 6289 1198 6309 1262
rect 10 1182 6309 1198
rect 10 1118 6225 1182
rect 6289 1118 6309 1182
rect 10 1102 6309 1118
rect 10 1038 6225 1102
rect 6289 1038 6309 1102
rect 10 1022 6309 1038
rect 10 958 6225 1022
rect 6289 958 6309 1022
rect 10 942 6309 958
rect 10 878 6225 942
rect 6289 878 6309 942
rect 10 862 6309 878
rect 10 798 6225 862
rect 6289 798 6309 862
rect 10 782 6309 798
rect 10 718 6225 782
rect 6289 718 6309 782
rect 10 702 6309 718
rect 10 638 6225 702
rect 6289 638 6309 702
rect 10 622 6309 638
rect 10 558 6225 622
rect 6289 558 6309 622
rect 10 542 6309 558
rect 10 478 6225 542
rect 6289 478 6309 542
rect 10 462 6309 478
rect 10 398 6225 462
rect 6289 398 6309 462
rect 10 382 6309 398
rect 10 318 6225 382
rect 6289 318 6309 382
rect 10 302 6309 318
rect 10 238 6225 302
rect 6289 238 6309 302
rect 10 222 6309 238
rect 10 158 6225 222
rect 6289 158 6309 222
rect 10 142 6309 158
rect 10 78 6225 142
rect 6289 78 6309 142
rect 10 50 6309 78
rect 6329 6222 12628 6250
rect 6329 6158 12544 6222
rect 12608 6158 12628 6222
rect 6329 6142 12628 6158
rect 6329 6078 12544 6142
rect 12608 6078 12628 6142
rect 6329 6062 12628 6078
rect 6329 5998 12544 6062
rect 12608 5998 12628 6062
rect 6329 5982 12628 5998
rect 6329 5918 12544 5982
rect 12608 5918 12628 5982
rect 6329 5902 12628 5918
rect 6329 5838 12544 5902
rect 12608 5838 12628 5902
rect 6329 5822 12628 5838
rect 6329 5758 12544 5822
rect 12608 5758 12628 5822
rect 6329 5742 12628 5758
rect 6329 5678 12544 5742
rect 12608 5678 12628 5742
rect 6329 5662 12628 5678
rect 6329 5598 12544 5662
rect 12608 5598 12628 5662
rect 6329 5582 12628 5598
rect 6329 5518 12544 5582
rect 12608 5518 12628 5582
rect 6329 5502 12628 5518
rect 6329 5438 12544 5502
rect 12608 5438 12628 5502
rect 6329 5422 12628 5438
rect 6329 5358 12544 5422
rect 12608 5358 12628 5422
rect 6329 5342 12628 5358
rect 6329 5278 12544 5342
rect 12608 5278 12628 5342
rect 6329 5262 12628 5278
rect 6329 5198 12544 5262
rect 12608 5198 12628 5262
rect 6329 5182 12628 5198
rect 6329 5118 12544 5182
rect 12608 5118 12628 5182
rect 6329 5102 12628 5118
rect 6329 5038 12544 5102
rect 12608 5038 12628 5102
rect 6329 5022 12628 5038
rect 6329 4958 12544 5022
rect 12608 4958 12628 5022
rect 6329 4942 12628 4958
rect 6329 4878 12544 4942
rect 12608 4878 12628 4942
rect 6329 4862 12628 4878
rect 6329 4798 12544 4862
rect 12608 4798 12628 4862
rect 6329 4782 12628 4798
rect 6329 4718 12544 4782
rect 12608 4718 12628 4782
rect 6329 4702 12628 4718
rect 6329 4638 12544 4702
rect 12608 4638 12628 4702
rect 6329 4622 12628 4638
rect 6329 4558 12544 4622
rect 12608 4558 12628 4622
rect 6329 4542 12628 4558
rect 6329 4478 12544 4542
rect 12608 4478 12628 4542
rect 6329 4462 12628 4478
rect 6329 4398 12544 4462
rect 12608 4398 12628 4462
rect 6329 4382 12628 4398
rect 6329 4318 12544 4382
rect 12608 4318 12628 4382
rect 6329 4302 12628 4318
rect 6329 4238 12544 4302
rect 12608 4238 12628 4302
rect 6329 4222 12628 4238
rect 6329 4158 12544 4222
rect 12608 4158 12628 4222
rect 6329 4142 12628 4158
rect 6329 4078 12544 4142
rect 12608 4078 12628 4142
rect 6329 4062 12628 4078
rect 6329 3998 12544 4062
rect 12608 3998 12628 4062
rect 6329 3982 12628 3998
rect 6329 3918 12544 3982
rect 12608 3918 12628 3982
rect 6329 3902 12628 3918
rect 6329 3838 12544 3902
rect 12608 3838 12628 3902
rect 6329 3822 12628 3838
rect 6329 3758 12544 3822
rect 12608 3758 12628 3822
rect 6329 3742 12628 3758
rect 6329 3678 12544 3742
rect 12608 3678 12628 3742
rect 6329 3662 12628 3678
rect 6329 3598 12544 3662
rect 12608 3598 12628 3662
rect 6329 3582 12628 3598
rect 6329 3518 12544 3582
rect 12608 3518 12628 3582
rect 6329 3502 12628 3518
rect 6329 3438 12544 3502
rect 12608 3438 12628 3502
rect 6329 3422 12628 3438
rect 6329 3358 12544 3422
rect 12608 3358 12628 3422
rect 6329 3342 12628 3358
rect 6329 3278 12544 3342
rect 12608 3278 12628 3342
rect 6329 3262 12628 3278
rect 6329 3198 12544 3262
rect 12608 3198 12628 3262
rect 6329 3182 12628 3198
rect 6329 3118 12544 3182
rect 12608 3118 12628 3182
rect 6329 3102 12628 3118
rect 6329 3038 12544 3102
rect 12608 3038 12628 3102
rect 6329 3022 12628 3038
rect 6329 2958 12544 3022
rect 12608 2958 12628 3022
rect 6329 2942 12628 2958
rect 6329 2878 12544 2942
rect 12608 2878 12628 2942
rect 6329 2862 12628 2878
rect 6329 2798 12544 2862
rect 12608 2798 12628 2862
rect 6329 2782 12628 2798
rect 6329 2718 12544 2782
rect 12608 2718 12628 2782
rect 6329 2702 12628 2718
rect 6329 2638 12544 2702
rect 12608 2638 12628 2702
rect 6329 2622 12628 2638
rect 6329 2558 12544 2622
rect 12608 2558 12628 2622
rect 6329 2542 12628 2558
rect 6329 2478 12544 2542
rect 12608 2478 12628 2542
rect 6329 2462 12628 2478
rect 6329 2398 12544 2462
rect 12608 2398 12628 2462
rect 6329 2382 12628 2398
rect 6329 2318 12544 2382
rect 12608 2318 12628 2382
rect 6329 2302 12628 2318
rect 6329 2238 12544 2302
rect 12608 2238 12628 2302
rect 6329 2222 12628 2238
rect 6329 2158 12544 2222
rect 12608 2158 12628 2222
rect 6329 2142 12628 2158
rect 6329 2078 12544 2142
rect 12608 2078 12628 2142
rect 6329 2062 12628 2078
rect 6329 1998 12544 2062
rect 12608 1998 12628 2062
rect 6329 1982 12628 1998
rect 6329 1918 12544 1982
rect 12608 1918 12628 1982
rect 6329 1902 12628 1918
rect 6329 1838 12544 1902
rect 12608 1838 12628 1902
rect 6329 1822 12628 1838
rect 6329 1758 12544 1822
rect 12608 1758 12628 1822
rect 6329 1742 12628 1758
rect 6329 1678 12544 1742
rect 12608 1678 12628 1742
rect 6329 1662 12628 1678
rect 6329 1598 12544 1662
rect 12608 1598 12628 1662
rect 6329 1582 12628 1598
rect 6329 1518 12544 1582
rect 12608 1518 12628 1582
rect 6329 1502 12628 1518
rect 6329 1438 12544 1502
rect 12608 1438 12628 1502
rect 6329 1422 12628 1438
rect 6329 1358 12544 1422
rect 12608 1358 12628 1422
rect 6329 1342 12628 1358
rect 6329 1278 12544 1342
rect 12608 1278 12628 1342
rect 6329 1262 12628 1278
rect 6329 1198 12544 1262
rect 12608 1198 12628 1262
rect 6329 1182 12628 1198
rect 6329 1118 12544 1182
rect 12608 1118 12628 1182
rect 6329 1102 12628 1118
rect 6329 1038 12544 1102
rect 12608 1038 12628 1102
rect 6329 1022 12628 1038
rect 6329 958 12544 1022
rect 12608 958 12628 1022
rect 6329 942 12628 958
rect 6329 878 12544 942
rect 12608 878 12628 942
rect 6329 862 12628 878
rect 6329 798 12544 862
rect 12608 798 12628 862
rect 6329 782 12628 798
rect 6329 718 12544 782
rect 12608 718 12628 782
rect 6329 702 12628 718
rect 6329 638 12544 702
rect 12608 638 12628 702
rect 6329 622 12628 638
rect 6329 558 12544 622
rect 12608 558 12628 622
rect 6329 542 12628 558
rect 6329 478 12544 542
rect 12608 478 12628 542
rect 6329 462 12628 478
rect 6329 398 12544 462
rect 12608 398 12628 462
rect 6329 382 12628 398
rect 6329 318 12544 382
rect 12608 318 12628 382
rect 6329 302 12628 318
rect 6329 238 12544 302
rect 12608 238 12628 302
rect 6329 222 12628 238
rect 6329 158 12544 222
rect 12608 158 12628 222
rect 6329 142 12628 158
rect 6329 78 12544 142
rect 12608 78 12628 142
rect 6329 50 12628 78
rect -12628 -78 -6329 -50
rect -12628 -142 -6413 -78
rect -6349 -142 -6329 -78
rect -12628 -158 -6329 -142
rect -12628 -222 -6413 -158
rect -6349 -222 -6329 -158
rect -12628 -238 -6329 -222
rect -12628 -302 -6413 -238
rect -6349 -302 -6329 -238
rect -12628 -318 -6329 -302
rect -12628 -382 -6413 -318
rect -6349 -382 -6329 -318
rect -12628 -398 -6329 -382
rect -12628 -462 -6413 -398
rect -6349 -462 -6329 -398
rect -12628 -478 -6329 -462
rect -12628 -542 -6413 -478
rect -6349 -542 -6329 -478
rect -12628 -558 -6329 -542
rect -12628 -622 -6413 -558
rect -6349 -622 -6329 -558
rect -12628 -638 -6329 -622
rect -12628 -702 -6413 -638
rect -6349 -702 -6329 -638
rect -12628 -718 -6329 -702
rect -12628 -782 -6413 -718
rect -6349 -782 -6329 -718
rect -12628 -798 -6329 -782
rect -12628 -862 -6413 -798
rect -6349 -862 -6329 -798
rect -12628 -878 -6329 -862
rect -12628 -942 -6413 -878
rect -6349 -942 -6329 -878
rect -12628 -958 -6329 -942
rect -12628 -1022 -6413 -958
rect -6349 -1022 -6329 -958
rect -12628 -1038 -6329 -1022
rect -12628 -1102 -6413 -1038
rect -6349 -1102 -6329 -1038
rect -12628 -1118 -6329 -1102
rect -12628 -1182 -6413 -1118
rect -6349 -1182 -6329 -1118
rect -12628 -1198 -6329 -1182
rect -12628 -1262 -6413 -1198
rect -6349 -1262 -6329 -1198
rect -12628 -1278 -6329 -1262
rect -12628 -1342 -6413 -1278
rect -6349 -1342 -6329 -1278
rect -12628 -1358 -6329 -1342
rect -12628 -1422 -6413 -1358
rect -6349 -1422 -6329 -1358
rect -12628 -1438 -6329 -1422
rect -12628 -1502 -6413 -1438
rect -6349 -1502 -6329 -1438
rect -12628 -1518 -6329 -1502
rect -12628 -1582 -6413 -1518
rect -6349 -1582 -6329 -1518
rect -12628 -1598 -6329 -1582
rect -12628 -1662 -6413 -1598
rect -6349 -1662 -6329 -1598
rect -12628 -1678 -6329 -1662
rect -12628 -1742 -6413 -1678
rect -6349 -1742 -6329 -1678
rect -12628 -1758 -6329 -1742
rect -12628 -1822 -6413 -1758
rect -6349 -1822 -6329 -1758
rect -12628 -1838 -6329 -1822
rect -12628 -1902 -6413 -1838
rect -6349 -1902 -6329 -1838
rect -12628 -1918 -6329 -1902
rect -12628 -1982 -6413 -1918
rect -6349 -1982 -6329 -1918
rect -12628 -1998 -6329 -1982
rect -12628 -2062 -6413 -1998
rect -6349 -2062 -6329 -1998
rect -12628 -2078 -6329 -2062
rect -12628 -2142 -6413 -2078
rect -6349 -2142 -6329 -2078
rect -12628 -2158 -6329 -2142
rect -12628 -2222 -6413 -2158
rect -6349 -2222 -6329 -2158
rect -12628 -2238 -6329 -2222
rect -12628 -2302 -6413 -2238
rect -6349 -2302 -6329 -2238
rect -12628 -2318 -6329 -2302
rect -12628 -2382 -6413 -2318
rect -6349 -2382 -6329 -2318
rect -12628 -2398 -6329 -2382
rect -12628 -2462 -6413 -2398
rect -6349 -2462 -6329 -2398
rect -12628 -2478 -6329 -2462
rect -12628 -2542 -6413 -2478
rect -6349 -2542 -6329 -2478
rect -12628 -2558 -6329 -2542
rect -12628 -2622 -6413 -2558
rect -6349 -2622 -6329 -2558
rect -12628 -2638 -6329 -2622
rect -12628 -2702 -6413 -2638
rect -6349 -2702 -6329 -2638
rect -12628 -2718 -6329 -2702
rect -12628 -2782 -6413 -2718
rect -6349 -2782 -6329 -2718
rect -12628 -2798 -6329 -2782
rect -12628 -2862 -6413 -2798
rect -6349 -2862 -6329 -2798
rect -12628 -2878 -6329 -2862
rect -12628 -2942 -6413 -2878
rect -6349 -2942 -6329 -2878
rect -12628 -2958 -6329 -2942
rect -12628 -3022 -6413 -2958
rect -6349 -3022 -6329 -2958
rect -12628 -3038 -6329 -3022
rect -12628 -3102 -6413 -3038
rect -6349 -3102 -6329 -3038
rect -12628 -3118 -6329 -3102
rect -12628 -3182 -6413 -3118
rect -6349 -3182 -6329 -3118
rect -12628 -3198 -6329 -3182
rect -12628 -3262 -6413 -3198
rect -6349 -3262 -6329 -3198
rect -12628 -3278 -6329 -3262
rect -12628 -3342 -6413 -3278
rect -6349 -3342 -6329 -3278
rect -12628 -3358 -6329 -3342
rect -12628 -3422 -6413 -3358
rect -6349 -3422 -6329 -3358
rect -12628 -3438 -6329 -3422
rect -12628 -3502 -6413 -3438
rect -6349 -3502 -6329 -3438
rect -12628 -3518 -6329 -3502
rect -12628 -3582 -6413 -3518
rect -6349 -3582 -6329 -3518
rect -12628 -3598 -6329 -3582
rect -12628 -3662 -6413 -3598
rect -6349 -3662 -6329 -3598
rect -12628 -3678 -6329 -3662
rect -12628 -3742 -6413 -3678
rect -6349 -3742 -6329 -3678
rect -12628 -3758 -6329 -3742
rect -12628 -3822 -6413 -3758
rect -6349 -3822 -6329 -3758
rect -12628 -3838 -6329 -3822
rect -12628 -3902 -6413 -3838
rect -6349 -3902 -6329 -3838
rect -12628 -3918 -6329 -3902
rect -12628 -3982 -6413 -3918
rect -6349 -3982 -6329 -3918
rect -12628 -3998 -6329 -3982
rect -12628 -4062 -6413 -3998
rect -6349 -4062 -6329 -3998
rect -12628 -4078 -6329 -4062
rect -12628 -4142 -6413 -4078
rect -6349 -4142 -6329 -4078
rect -12628 -4158 -6329 -4142
rect -12628 -4222 -6413 -4158
rect -6349 -4222 -6329 -4158
rect -12628 -4238 -6329 -4222
rect -12628 -4302 -6413 -4238
rect -6349 -4302 -6329 -4238
rect -12628 -4318 -6329 -4302
rect -12628 -4382 -6413 -4318
rect -6349 -4382 -6329 -4318
rect -12628 -4398 -6329 -4382
rect -12628 -4462 -6413 -4398
rect -6349 -4462 -6329 -4398
rect -12628 -4478 -6329 -4462
rect -12628 -4542 -6413 -4478
rect -6349 -4542 -6329 -4478
rect -12628 -4558 -6329 -4542
rect -12628 -4622 -6413 -4558
rect -6349 -4622 -6329 -4558
rect -12628 -4638 -6329 -4622
rect -12628 -4702 -6413 -4638
rect -6349 -4702 -6329 -4638
rect -12628 -4718 -6329 -4702
rect -12628 -4782 -6413 -4718
rect -6349 -4782 -6329 -4718
rect -12628 -4798 -6329 -4782
rect -12628 -4862 -6413 -4798
rect -6349 -4862 -6329 -4798
rect -12628 -4878 -6329 -4862
rect -12628 -4942 -6413 -4878
rect -6349 -4942 -6329 -4878
rect -12628 -4958 -6329 -4942
rect -12628 -5022 -6413 -4958
rect -6349 -5022 -6329 -4958
rect -12628 -5038 -6329 -5022
rect -12628 -5102 -6413 -5038
rect -6349 -5102 -6329 -5038
rect -12628 -5118 -6329 -5102
rect -12628 -5182 -6413 -5118
rect -6349 -5182 -6329 -5118
rect -12628 -5198 -6329 -5182
rect -12628 -5262 -6413 -5198
rect -6349 -5262 -6329 -5198
rect -12628 -5278 -6329 -5262
rect -12628 -5342 -6413 -5278
rect -6349 -5342 -6329 -5278
rect -12628 -5358 -6329 -5342
rect -12628 -5422 -6413 -5358
rect -6349 -5422 -6329 -5358
rect -12628 -5438 -6329 -5422
rect -12628 -5502 -6413 -5438
rect -6349 -5502 -6329 -5438
rect -12628 -5518 -6329 -5502
rect -12628 -5582 -6413 -5518
rect -6349 -5582 -6329 -5518
rect -12628 -5598 -6329 -5582
rect -12628 -5662 -6413 -5598
rect -6349 -5662 -6329 -5598
rect -12628 -5678 -6329 -5662
rect -12628 -5742 -6413 -5678
rect -6349 -5742 -6329 -5678
rect -12628 -5758 -6329 -5742
rect -12628 -5822 -6413 -5758
rect -6349 -5822 -6329 -5758
rect -12628 -5838 -6329 -5822
rect -12628 -5902 -6413 -5838
rect -6349 -5902 -6329 -5838
rect -12628 -5918 -6329 -5902
rect -12628 -5982 -6413 -5918
rect -6349 -5982 -6329 -5918
rect -12628 -5998 -6329 -5982
rect -12628 -6062 -6413 -5998
rect -6349 -6062 -6329 -5998
rect -12628 -6078 -6329 -6062
rect -12628 -6142 -6413 -6078
rect -6349 -6142 -6329 -6078
rect -12628 -6158 -6329 -6142
rect -12628 -6222 -6413 -6158
rect -6349 -6222 -6329 -6158
rect -12628 -6250 -6329 -6222
rect -6309 -78 -10 -50
rect -6309 -142 -94 -78
rect -30 -142 -10 -78
rect -6309 -158 -10 -142
rect -6309 -222 -94 -158
rect -30 -222 -10 -158
rect -6309 -238 -10 -222
rect -6309 -302 -94 -238
rect -30 -302 -10 -238
rect -6309 -318 -10 -302
rect -6309 -382 -94 -318
rect -30 -382 -10 -318
rect -6309 -398 -10 -382
rect -6309 -462 -94 -398
rect -30 -462 -10 -398
rect -6309 -478 -10 -462
rect -6309 -542 -94 -478
rect -30 -542 -10 -478
rect -6309 -558 -10 -542
rect -6309 -622 -94 -558
rect -30 -622 -10 -558
rect -6309 -638 -10 -622
rect -6309 -702 -94 -638
rect -30 -702 -10 -638
rect -6309 -718 -10 -702
rect -6309 -782 -94 -718
rect -30 -782 -10 -718
rect -6309 -798 -10 -782
rect -6309 -862 -94 -798
rect -30 -862 -10 -798
rect -6309 -878 -10 -862
rect -6309 -942 -94 -878
rect -30 -942 -10 -878
rect -6309 -958 -10 -942
rect -6309 -1022 -94 -958
rect -30 -1022 -10 -958
rect -6309 -1038 -10 -1022
rect -6309 -1102 -94 -1038
rect -30 -1102 -10 -1038
rect -6309 -1118 -10 -1102
rect -6309 -1182 -94 -1118
rect -30 -1182 -10 -1118
rect -6309 -1198 -10 -1182
rect -6309 -1262 -94 -1198
rect -30 -1262 -10 -1198
rect -6309 -1278 -10 -1262
rect -6309 -1342 -94 -1278
rect -30 -1342 -10 -1278
rect -6309 -1358 -10 -1342
rect -6309 -1422 -94 -1358
rect -30 -1422 -10 -1358
rect -6309 -1438 -10 -1422
rect -6309 -1502 -94 -1438
rect -30 -1502 -10 -1438
rect -6309 -1518 -10 -1502
rect -6309 -1582 -94 -1518
rect -30 -1582 -10 -1518
rect -6309 -1598 -10 -1582
rect -6309 -1662 -94 -1598
rect -30 -1662 -10 -1598
rect -6309 -1678 -10 -1662
rect -6309 -1742 -94 -1678
rect -30 -1742 -10 -1678
rect -6309 -1758 -10 -1742
rect -6309 -1822 -94 -1758
rect -30 -1822 -10 -1758
rect -6309 -1838 -10 -1822
rect -6309 -1902 -94 -1838
rect -30 -1902 -10 -1838
rect -6309 -1918 -10 -1902
rect -6309 -1982 -94 -1918
rect -30 -1982 -10 -1918
rect -6309 -1998 -10 -1982
rect -6309 -2062 -94 -1998
rect -30 -2062 -10 -1998
rect -6309 -2078 -10 -2062
rect -6309 -2142 -94 -2078
rect -30 -2142 -10 -2078
rect -6309 -2158 -10 -2142
rect -6309 -2222 -94 -2158
rect -30 -2222 -10 -2158
rect -6309 -2238 -10 -2222
rect -6309 -2302 -94 -2238
rect -30 -2302 -10 -2238
rect -6309 -2318 -10 -2302
rect -6309 -2382 -94 -2318
rect -30 -2382 -10 -2318
rect -6309 -2398 -10 -2382
rect -6309 -2462 -94 -2398
rect -30 -2462 -10 -2398
rect -6309 -2478 -10 -2462
rect -6309 -2542 -94 -2478
rect -30 -2542 -10 -2478
rect -6309 -2558 -10 -2542
rect -6309 -2622 -94 -2558
rect -30 -2622 -10 -2558
rect -6309 -2638 -10 -2622
rect -6309 -2702 -94 -2638
rect -30 -2702 -10 -2638
rect -6309 -2718 -10 -2702
rect -6309 -2782 -94 -2718
rect -30 -2782 -10 -2718
rect -6309 -2798 -10 -2782
rect -6309 -2862 -94 -2798
rect -30 -2862 -10 -2798
rect -6309 -2878 -10 -2862
rect -6309 -2942 -94 -2878
rect -30 -2942 -10 -2878
rect -6309 -2958 -10 -2942
rect -6309 -3022 -94 -2958
rect -30 -3022 -10 -2958
rect -6309 -3038 -10 -3022
rect -6309 -3102 -94 -3038
rect -30 -3102 -10 -3038
rect -6309 -3118 -10 -3102
rect -6309 -3182 -94 -3118
rect -30 -3182 -10 -3118
rect -6309 -3198 -10 -3182
rect -6309 -3262 -94 -3198
rect -30 -3262 -10 -3198
rect -6309 -3278 -10 -3262
rect -6309 -3342 -94 -3278
rect -30 -3342 -10 -3278
rect -6309 -3358 -10 -3342
rect -6309 -3422 -94 -3358
rect -30 -3422 -10 -3358
rect -6309 -3438 -10 -3422
rect -6309 -3502 -94 -3438
rect -30 -3502 -10 -3438
rect -6309 -3518 -10 -3502
rect -6309 -3582 -94 -3518
rect -30 -3582 -10 -3518
rect -6309 -3598 -10 -3582
rect -6309 -3662 -94 -3598
rect -30 -3662 -10 -3598
rect -6309 -3678 -10 -3662
rect -6309 -3742 -94 -3678
rect -30 -3742 -10 -3678
rect -6309 -3758 -10 -3742
rect -6309 -3822 -94 -3758
rect -30 -3822 -10 -3758
rect -6309 -3838 -10 -3822
rect -6309 -3902 -94 -3838
rect -30 -3902 -10 -3838
rect -6309 -3918 -10 -3902
rect -6309 -3982 -94 -3918
rect -30 -3982 -10 -3918
rect -6309 -3998 -10 -3982
rect -6309 -4062 -94 -3998
rect -30 -4062 -10 -3998
rect -6309 -4078 -10 -4062
rect -6309 -4142 -94 -4078
rect -30 -4142 -10 -4078
rect -6309 -4158 -10 -4142
rect -6309 -4222 -94 -4158
rect -30 -4222 -10 -4158
rect -6309 -4238 -10 -4222
rect -6309 -4302 -94 -4238
rect -30 -4302 -10 -4238
rect -6309 -4318 -10 -4302
rect -6309 -4382 -94 -4318
rect -30 -4382 -10 -4318
rect -6309 -4398 -10 -4382
rect -6309 -4462 -94 -4398
rect -30 -4462 -10 -4398
rect -6309 -4478 -10 -4462
rect -6309 -4542 -94 -4478
rect -30 -4542 -10 -4478
rect -6309 -4558 -10 -4542
rect -6309 -4622 -94 -4558
rect -30 -4622 -10 -4558
rect -6309 -4638 -10 -4622
rect -6309 -4702 -94 -4638
rect -30 -4702 -10 -4638
rect -6309 -4718 -10 -4702
rect -6309 -4782 -94 -4718
rect -30 -4782 -10 -4718
rect -6309 -4798 -10 -4782
rect -6309 -4862 -94 -4798
rect -30 -4862 -10 -4798
rect -6309 -4878 -10 -4862
rect -6309 -4942 -94 -4878
rect -30 -4942 -10 -4878
rect -6309 -4958 -10 -4942
rect -6309 -5022 -94 -4958
rect -30 -5022 -10 -4958
rect -6309 -5038 -10 -5022
rect -6309 -5102 -94 -5038
rect -30 -5102 -10 -5038
rect -6309 -5118 -10 -5102
rect -6309 -5182 -94 -5118
rect -30 -5182 -10 -5118
rect -6309 -5198 -10 -5182
rect -6309 -5262 -94 -5198
rect -30 -5262 -10 -5198
rect -6309 -5278 -10 -5262
rect -6309 -5342 -94 -5278
rect -30 -5342 -10 -5278
rect -6309 -5358 -10 -5342
rect -6309 -5422 -94 -5358
rect -30 -5422 -10 -5358
rect -6309 -5438 -10 -5422
rect -6309 -5502 -94 -5438
rect -30 -5502 -10 -5438
rect -6309 -5518 -10 -5502
rect -6309 -5582 -94 -5518
rect -30 -5582 -10 -5518
rect -6309 -5598 -10 -5582
rect -6309 -5662 -94 -5598
rect -30 -5662 -10 -5598
rect -6309 -5678 -10 -5662
rect -6309 -5742 -94 -5678
rect -30 -5742 -10 -5678
rect -6309 -5758 -10 -5742
rect -6309 -5822 -94 -5758
rect -30 -5822 -10 -5758
rect -6309 -5838 -10 -5822
rect -6309 -5902 -94 -5838
rect -30 -5902 -10 -5838
rect -6309 -5918 -10 -5902
rect -6309 -5982 -94 -5918
rect -30 -5982 -10 -5918
rect -6309 -5998 -10 -5982
rect -6309 -6062 -94 -5998
rect -30 -6062 -10 -5998
rect -6309 -6078 -10 -6062
rect -6309 -6142 -94 -6078
rect -30 -6142 -10 -6078
rect -6309 -6158 -10 -6142
rect -6309 -6222 -94 -6158
rect -30 -6222 -10 -6158
rect -6309 -6250 -10 -6222
rect 10 -78 6309 -50
rect 10 -142 6225 -78
rect 6289 -142 6309 -78
rect 10 -158 6309 -142
rect 10 -222 6225 -158
rect 6289 -222 6309 -158
rect 10 -238 6309 -222
rect 10 -302 6225 -238
rect 6289 -302 6309 -238
rect 10 -318 6309 -302
rect 10 -382 6225 -318
rect 6289 -382 6309 -318
rect 10 -398 6309 -382
rect 10 -462 6225 -398
rect 6289 -462 6309 -398
rect 10 -478 6309 -462
rect 10 -542 6225 -478
rect 6289 -542 6309 -478
rect 10 -558 6309 -542
rect 10 -622 6225 -558
rect 6289 -622 6309 -558
rect 10 -638 6309 -622
rect 10 -702 6225 -638
rect 6289 -702 6309 -638
rect 10 -718 6309 -702
rect 10 -782 6225 -718
rect 6289 -782 6309 -718
rect 10 -798 6309 -782
rect 10 -862 6225 -798
rect 6289 -862 6309 -798
rect 10 -878 6309 -862
rect 10 -942 6225 -878
rect 6289 -942 6309 -878
rect 10 -958 6309 -942
rect 10 -1022 6225 -958
rect 6289 -1022 6309 -958
rect 10 -1038 6309 -1022
rect 10 -1102 6225 -1038
rect 6289 -1102 6309 -1038
rect 10 -1118 6309 -1102
rect 10 -1182 6225 -1118
rect 6289 -1182 6309 -1118
rect 10 -1198 6309 -1182
rect 10 -1262 6225 -1198
rect 6289 -1262 6309 -1198
rect 10 -1278 6309 -1262
rect 10 -1342 6225 -1278
rect 6289 -1342 6309 -1278
rect 10 -1358 6309 -1342
rect 10 -1422 6225 -1358
rect 6289 -1422 6309 -1358
rect 10 -1438 6309 -1422
rect 10 -1502 6225 -1438
rect 6289 -1502 6309 -1438
rect 10 -1518 6309 -1502
rect 10 -1582 6225 -1518
rect 6289 -1582 6309 -1518
rect 10 -1598 6309 -1582
rect 10 -1662 6225 -1598
rect 6289 -1662 6309 -1598
rect 10 -1678 6309 -1662
rect 10 -1742 6225 -1678
rect 6289 -1742 6309 -1678
rect 10 -1758 6309 -1742
rect 10 -1822 6225 -1758
rect 6289 -1822 6309 -1758
rect 10 -1838 6309 -1822
rect 10 -1902 6225 -1838
rect 6289 -1902 6309 -1838
rect 10 -1918 6309 -1902
rect 10 -1982 6225 -1918
rect 6289 -1982 6309 -1918
rect 10 -1998 6309 -1982
rect 10 -2062 6225 -1998
rect 6289 -2062 6309 -1998
rect 10 -2078 6309 -2062
rect 10 -2142 6225 -2078
rect 6289 -2142 6309 -2078
rect 10 -2158 6309 -2142
rect 10 -2222 6225 -2158
rect 6289 -2222 6309 -2158
rect 10 -2238 6309 -2222
rect 10 -2302 6225 -2238
rect 6289 -2302 6309 -2238
rect 10 -2318 6309 -2302
rect 10 -2382 6225 -2318
rect 6289 -2382 6309 -2318
rect 10 -2398 6309 -2382
rect 10 -2462 6225 -2398
rect 6289 -2462 6309 -2398
rect 10 -2478 6309 -2462
rect 10 -2542 6225 -2478
rect 6289 -2542 6309 -2478
rect 10 -2558 6309 -2542
rect 10 -2622 6225 -2558
rect 6289 -2622 6309 -2558
rect 10 -2638 6309 -2622
rect 10 -2702 6225 -2638
rect 6289 -2702 6309 -2638
rect 10 -2718 6309 -2702
rect 10 -2782 6225 -2718
rect 6289 -2782 6309 -2718
rect 10 -2798 6309 -2782
rect 10 -2862 6225 -2798
rect 6289 -2862 6309 -2798
rect 10 -2878 6309 -2862
rect 10 -2942 6225 -2878
rect 6289 -2942 6309 -2878
rect 10 -2958 6309 -2942
rect 10 -3022 6225 -2958
rect 6289 -3022 6309 -2958
rect 10 -3038 6309 -3022
rect 10 -3102 6225 -3038
rect 6289 -3102 6309 -3038
rect 10 -3118 6309 -3102
rect 10 -3182 6225 -3118
rect 6289 -3182 6309 -3118
rect 10 -3198 6309 -3182
rect 10 -3262 6225 -3198
rect 6289 -3262 6309 -3198
rect 10 -3278 6309 -3262
rect 10 -3342 6225 -3278
rect 6289 -3342 6309 -3278
rect 10 -3358 6309 -3342
rect 10 -3422 6225 -3358
rect 6289 -3422 6309 -3358
rect 10 -3438 6309 -3422
rect 10 -3502 6225 -3438
rect 6289 -3502 6309 -3438
rect 10 -3518 6309 -3502
rect 10 -3582 6225 -3518
rect 6289 -3582 6309 -3518
rect 10 -3598 6309 -3582
rect 10 -3662 6225 -3598
rect 6289 -3662 6309 -3598
rect 10 -3678 6309 -3662
rect 10 -3742 6225 -3678
rect 6289 -3742 6309 -3678
rect 10 -3758 6309 -3742
rect 10 -3822 6225 -3758
rect 6289 -3822 6309 -3758
rect 10 -3838 6309 -3822
rect 10 -3902 6225 -3838
rect 6289 -3902 6309 -3838
rect 10 -3918 6309 -3902
rect 10 -3982 6225 -3918
rect 6289 -3982 6309 -3918
rect 10 -3998 6309 -3982
rect 10 -4062 6225 -3998
rect 6289 -4062 6309 -3998
rect 10 -4078 6309 -4062
rect 10 -4142 6225 -4078
rect 6289 -4142 6309 -4078
rect 10 -4158 6309 -4142
rect 10 -4222 6225 -4158
rect 6289 -4222 6309 -4158
rect 10 -4238 6309 -4222
rect 10 -4302 6225 -4238
rect 6289 -4302 6309 -4238
rect 10 -4318 6309 -4302
rect 10 -4382 6225 -4318
rect 6289 -4382 6309 -4318
rect 10 -4398 6309 -4382
rect 10 -4462 6225 -4398
rect 6289 -4462 6309 -4398
rect 10 -4478 6309 -4462
rect 10 -4542 6225 -4478
rect 6289 -4542 6309 -4478
rect 10 -4558 6309 -4542
rect 10 -4622 6225 -4558
rect 6289 -4622 6309 -4558
rect 10 -4638 6309 -4622
rect 10 -4702 6225 -4638
rect 6289 -4702 6309 -4638
rect 10 -4718 6309 -4702
rect 10 -4782 6225 -4718
rect 6289 -4782 6309 -4718
rect 10 -4798 6309 -4782
rect 10 -4862 6225 -4798
rect 6289 -4862 6309 -4798
rect 10 -4878 6309 -4862
rect 10 -4942 6225 -4878
rect 6289 -4942 6309 -4878
rect 10 -4958 6309 -4942
rect 10 -5022 6225 -4958
rect 6289 -5022 6309 -4958
rect 10 -5038 6309 -5022
rect 10 -5102 6225 -5038
rect 6289 -5102 6309 -5038
rect 10 -5118 6309 -5102
rect 10 -5182 6225 -5118
rect 6289 -5182 6309 -5118
rect 10 -5198 6309 -5182
rect 10 -5262 6225 -5198
rect 6289 -5262 6309 -5198
rect 10 -5278 6309 -5262
rect 10 -5342 6225 -5278
rect 6289 -5342 6309 -5278
rect 10 -5358 6309 -5342
rect 10 -5422 6225 -5358
rect 6289 -5422 6309 -5358
rect 10 -5438 6309 -5422
rect 10 -5502 6225 -5438
rect 6289 -5502 6309 -5438
rect 10 -5518 6309 -5502
rect 10 -5582 6225 -5518
rect 6289 -5582 6309 -5518
rect 10 -5598 6309 -5582
rect 10 -5662 6225 -5598
rect 6289 -5662 6309 -5598
rect 10 -5678 6309 -5662
rect 10 -5742 6225 -5678
rect 6289 -5742 6309 -5678
rect 10 -5758 6309 -5742
rect 10 -5822 6225 -5758
rect 6289 -5822 6309 -5758
rect 10 -5838 6309 -5822
rect 10 -5902 6225 -5838
rect 6289 -5902 6309 -5838
rect 10 -5918 6309 -5902
rect 10 -5982 6225 -5918
rect 6289 -5982 6309 -5918
rect 10 -5998 6309 -5982
rect 10 -6062 6225 -5998
rect 6289 -6062 6309 -5998
rect 10 -6078 6309 -6062
rect 10 -6142 6225 -6078
rect 6289 -6142 6309 -6078
rect 10 -6158 6309 -6142
rect 10 -6222 6225 -6158
rect 6289 -6222 6309 -6158
rect 10 -6250 6309 -6222
rect 6329 -78 12628 -50
rect 6329 -142 12544 -78
rect 12608 -142 12628 -78
rect 6329 -158 12628 -142
rect 6329 -222 12544 -158
rect 12608 -222 12628 -158
rect 6329 -238 12628 -222
rect 6329 -302 12544 -238
rect 12608 -302 12628 -238
rect 6329 -318 12628 -302
rect 6329 -382 12544 -318
rect 12608 -382 12628 -318
rect 6329 -398 12628 -382
rect 6329 -462 12544 -398
rect 12608 -462 12628 -398
rect 6329 -478 12628 -462
rect 6329 -542 12544 -478
rect 12608 -542 12628 -478
rect 6329 -558 12628 -542
rect 6329 -622 12544 -558
rect 12608 -622 12628 -558
rect 6329 -638 12628 -622
rect 6329 -702 12544 -638
rect 12608 -702 12628 -638
rect 6329 -718 12628 -702
rect 6329 -782 12544 -718
rect 12608 -782 12628 -718
rect 6329 -798 12628 -782
rect 6329 -862 12544 -798
rect 12608 -862 12628 -798
rect 6329 -878 12628 -862
rect 6329 -942 12544 -878
rect 12608 -942 12628 -878
rect 6329 -958 12628 -942
rect 6329 -1022 12544 -958
rect 12608 -1022 12628 -958
rect 6329 -1038 12628 -1022
rect 6329 -1102 12544 -1038
rect 12608 -1102 12628 -1038
rect 6329 -1118 12628 -1102
rect 6329 -1182 12544 -1118
rect 12608 -1182 12628 -1118
rect 6329 -1198 12628 -1182
rect 6329 -1262 12544 -1198
rect 12608 -1262 12628 -1198
rect 6329 -1278 12628 -1262
rect 6329 -1342 12544 -1278
rect 12608 -1342 12628 -1278
rect 6329 -1358 12628 -1342
rect 6329 -1422 12544 -1358
rect 12608 -1422 12628 -1358
rect 6329 -1438 12628 -1422
rect 6329 -1502 12544 -1438
rect 12608 -1502 12628 -1438
rect 6329 -1518 12628 -1502
rect 6329 -1582 12544 -1518
rect 12608 -1582 12628 -1518
rect 6329 -1598 12628 -1582
rect 6329 -1662 12544 -1598
rect 12608 -1662 12628 -1598
rect 6329 -1678 12628 -1662
rect 6329 -1742 12544 -1678
rect 12608 -1742 12628 -1678
rect 6329 -1758 12628 -1742
rect 6329 -1822 12544 -1758
rect 12608 -1822 12628 -1758
rect 6329 -1838 12628 -1822
rect 6329 -1902 12544 -1838
rect 12608 -1902 12628 -1838
rect 6329 -1918 12628 -1902
rect 6329 -1982 12544 -1918
rect 12608 -1982 12628 -1918
rect 6329 -1998 12628 -1982
rect 6329 -2062 12544 -1998
rect 12608 -2062 12628 -1998
rect 6329 -2078 12628 -2062
rect 6329 -2142 12544 -2078
rect 12608 -2142 12628 -2078
rect 6329 -2158 12628 -2142
rect 6329 -2222 12544 -2158
rect 12608 -2222 12628 -2158
rect 6329 -2238 12628 -2222
rect 6329 -2302 12544 -2238
rect 12608 -2302 12628 -2238
rect 6329 -2318 12628 -2302
rect 6329 -2382 12544 -2318
rect 12608 -2382 12628 -2318
rect 6329 -2398 12628 -2382
rect 6329 -2462 12544 -2398
rect 12608 -2462 12628 -2398
rect 6329 -2478 12628 -2462
rect 6329 -2542 12544 -2478
rect 12608 -2542 12628 -2478
rect 6329 -2558 12628 -2542
rect 6329 -2622 12544 -2558
rect 12608 -2622 12628 -2558
rect 6329 -2638 12628 -2622
rect 6329 -2702 12544 -2638
rect 12608 -2702 12628 -2638
rect 6329 -2718 12628 -2702
rect 6329 -2782 12544 -2718
rect 12608 -2782 12628 -2718
rect 6329 -2798 12628 -2782
rect 6329 -2862 12544 -2798
rect 12608 -2862 12628 -2798
rect 6329 -2878 12628 -2862
rect 6329 -2942 12544 -2878
rect 12608 -2942 12628 -2878
rect 6329 -2958 12628 -2942
rect 6329 -3022 12544 -2958
rect 12608 -3022 12628 -2958
rect 6329 -3038 12628 -3022
rect 6329 -3102 12544 -3038
rect 12608 -3102 12628 -3038
rect 6329 -3118 12628 -3102
rect 6329 -3182 12544 -3118
rect 12608 -3182 12628 -3118
rect 6329 -3198 12628 -3182
rect 6329 -3262 12544 -3198
rect 12608 -3262 12628 -3198
rect 6329 -3278 12628 -3262
rect 6329 -3342 12544 -3278
rect 12608 -3342 12628 -3278
rect 6329 -3358 12628 -3342
rect 6329 -3422 12544 -3358
rect 12608 -3422 12628 -3358
rect 6329 -3438 12628 -3422
rect 6329 -3502 12544 -3438
rect 12608 -3502 12628 -3438
rect 6329 -3518 12628 -3502
rect 6329 -3582 12544 -3518
rect 12608 -3582 12628 -3518
rect 6329 -3598 12628 -3582
rect 6329 -3662 12544 -3598
rect 12608 -3662 12628 -3598
rect 6329 -3678 12628 -3662
rect 6329 -3742 12544 -3678
rect 12608 -3742 12628 -3678
rect 6329 -3758 12628 -3742
rect 6329 -3822 12544 -3758
rect 12608 -3822 12628 -3758
rect 6329 -3838 12628 -3822
rect 6329 -3902 12544 -3838
rect 12608 -3902 12628 -3838
rect 6329 -3918 12628 -3902
rect 6329 -3982 12544 -3918
rect 12608 -3982 12628 -3918
rect 6329 -3998 12628 -3982
rect 6329 -4062 12544 -3998
rect 12608 -4062 12628 -3998
rect 6329 -4078 12628 -4062
rect 6329 -4142 12544 -4078
rect 12608 -4142 12628 -4078
rect 6329 -4158 12628 -4142
rect 6329 -4222 12544 -4158
rect 12608 -4222 12628 -4158
rect 6329 -4238 12628 -4222
rect 6329 -4302 12544 -4238
rect 12608 -4302 12628 -4238
rect 6329 -4318 12628 -4302
rect 6329 -4382 12544 -4318
rect 12608 -4382 12628 -4318
rect 6329 -4398 12628 -4382
rect 6329 -4462 12544 -4398
rect 12608 -4462 12628 -4398
rect 6329 -4478 12628 -4462
rect 6329 -4542 12544 -4478
rect 12608 -4542 12628 -4478
rect 6329 -4558 12628 -4542
rect 6329 -4622 12544 -4558
rect 12608 -4622 12628 -4558
rect 6329 -4638 12628 -4622
rect 6329 -4702 12544 -4638
rect 12608 -4702 12628 -4638
rect 6329 -4718 12628 -4702
rect 6329 -4782 12544 -4718
rect 12608 -4782 12628 -4718
rect 6329 -4798 12628 -4782
rect 6329 -4862 12544 -4798
rect 12608 -4862 12628 -4798
rect 6329 -4878 12628 -4862
rect 6329 -4942 12544 -4878
rect 12608 -4942 12628 -4878
rect 6329 -4958 12628 -4942
rect 6329 -5022 12544 -4958
rect 12608 -5022 12628 -4958
rect 6329 -5038 12628 -5022
rect 6329 -5102 12544 -5038
rect 12608 -5102 12628 -5038
rect 6329 -5118 12628 -5102
rect 6329 -5182 12544 -5118
rect 12608 -5182 12628 -5118
rect 6329 -5198 12628 -5182
rect 6329 -5262 12544 -5198
rect 12608 -5262 12628 -5198
rect 6329 -5278 12628 -5262
rect 6329 -5342 12544 -5278
rect 12608 -5342 12628 -5278
rect 6329 -5358 12628 -5342
rect 6329 -5422 12544 -5358
rect 12608 -5422 12628 -5358
rect 6329 -5438 12628 -5422
rect 6329 -5502 12544 -5438
rect 12608 -5502 12628 -5438
rect 6329 -5518 12628 -5502
rect 6329 -5582 12544 -5518
rect 12608 -5582 12628 -5518
rect 6329 -5598 12628 -5582
rect 6329 -5662 12544 -5598
rect 12608 -5662 12628 -5598
rect 6329 -5678 12628 -5662
rect 6329 -5742 12544 -5678
rect 12608 -5742 12628 -5678
rect 6329 -5758 12628 -5742
rect 6329 -5822 12544 -5758
rect 12608 -5822 12628 -5758
rect 6329 -5838 12628 -5822
rect 6329 -5902 12544 -5838
rect 12608 -5902 12628 -5838
rect 6329 -5918 12628 -5902
rect 6329 -5982 12544 -5918
rect 12608 -5982 12628 -5918
rect 6329 -5998 12628 -5982
rect 6329 -6062 12544 -5998
rect 12608 -6062 12628 -5998
rect 6329 -6078 12628 -6062
rect 6329 -6142 12544 -6078
rect 12608 -6142 12628 -6078
rect 6329 -6158 12628 -6142
rect 6329 -6222 12544 -6158
rect 12608 -6222 12628 -6158
rect 6329 -6250 12628 -6222
rect -12628 -6378 -6329 -6350
rect -12628 -6442 -6413 -6378
rect -6349 -6442 -6329 -6378
rect -12628 -6458 -6329 -6442
rect -12628 -6522 -6413 -6458
rect -6349 -6522 -6329 -6458
rect -12628 -6538 -6329 -6522
rect -12628 -6602 -6413 -6538
rect -6349 -6602 -6329 -6538
rect -12628 -6618 -6329 -6602
rect -12628 -6682 -6413 -6618
rect -6349 -6682 -6329 -6618
rect -12628 -6698 -6329 -6682
rect -12628 -6762 -6413 -6698
rect -6349 -6762 -6329 -6698
rect -12628 -6778 -6329 -6762
rect -12628 -6842 -6413 -6778
rect -6349 -6842 -6329 -6778
rect -12628 -6858 -6329 -6842
rect -12628 -6922 -6413 -6858
rect -6349 -6922 -6329 -6858
rect -12628 -6938 -6329 -6922
rect -12628 -7002 -6413 -6938
rect -6349 -7002 -6329 -6938
rect -12628 -7018 -6329 -7002
rect -12628 -7082 -6413 -7018
rect -6349 -7082 -6329 -7018
rect -12628 -7098 -6329 -7082
rect -12628 -7162 -6413 -7098
rect -6349 -7162 -6329 -7098
rect -12628 -7178 -6329 -7162
rect -12628 -7242 -6413 -7178
rect -6349 -7242 -6329 -7178
rect -12628 -7258 -6329 -7242
rect -12628 -7322 -6413 -7258
rect -6349 -7322 -6329 -7258
rect -12628 -7338 -6329 -7322
rect -12628 -7402 -6413 -7338
rect -6349 -7402 -6329 -7338
rect -12628 -7418 -6329 -7402
rect -12628 -7482 -6413 -7418
rect -6349 -7482 -6329 -7418
rect -12628 -7498 -6329 -7482
rect -12628 -7562 -6413 -7498
rect -6349 -7562 -6329 -7498
rect -12628 -7578 -6329 -7562
rect -12628 -7642 -6413 -7578
rect -6349 -7642 -6329 -7578
rect -12628 -7658 -6329 -7642
rect -12628 -7722 -6413 -7658
rect -6349 -7722 -6329 -7658
rect -12628 -7738 -6329 -7722
rect -12628 -7802 -6413 -7738
rect -6349 -7802 -6329 -7738
rect -12628 -7818 -6329 -7802
rect -12628 -7882 -6413 -7818
rect -6349 -7882 -6329 -7818
rect -12628 -7898 -6329 -7882
rect -12628 -7962 -6413 -7898
rect -6349 -7962 -6329 -7898
rect -12628 -7978 -6329 -7962
rect -12628 -8042 -6413 -7978
rect -6349 -8042 -6329 -7978
rect -12628 -8058 -6329 -8042
rect -12628 -8122 -6413 -8058
rect -6349 -8122 -6329 -8058
rect -12628 -8138 -6329 -8122
rect -12628 -8202 -6413 -8138
rect -6349 -8202 -6329 -8138
rect -12628 -8218 -6329 -8202
rect -12628 -8282 -6413 -8218
rect -6349 -8282 -6329 -8218
rect -12628 -8298 -6329 -8282
rect -12628 -8362 -6413 -8298
rect -6349 -8362 -6329 -8298
rect -12628 -8378 -6329 -8362
rect -12628 -8442 -6413 -8378
rect -6349 -8442 -6329 -8378
rect -12628 -8458 -6329 -8442
rect -12628 -8522 -6413 -8458
rect -6349 -8522 -6329 -8458
rect -12628 -8538 -6329 -8522
rect -12628 -8602 -6413 -8538
rect -6349 -8602 -6329 -8538
rect -12628 -8618 -6329 -8602
rect -12628 -8682 -6413 -8618
rect -6349 -8682 -6329 -8618
rect -12628 -8698 -6329 -8682
rect -12628 -8762 -6413 -8698
rect -6349 -8762 -6329 -8698
rect -12628 -8778 -6329 -8762
rect -12628 -8842 -6413 -8778
rect -6349 -8842 -6329 -8778
rect -12628 -8858 -6329 -8842
rect -12628 -8922 -6413 -8858
rect -6349 -8922 -6329 -8858
rect -12628 -8938 -6329 -8922
rect -12628 -9002 -6413 -8938
rect -6349 -9002 -6329 -8938
rect -12628 -9018 -6329 -9002
rect -12628 -9082 -6413 -9018
rect -6349 -9082 -6329 -9018
rect -12628 -9098 -6329 -9082
rect -12628 -9162 -6413 -9098
rect -6349 -9162 -6329 -9098
rect -12628 -9178 -6329 -9162
rect -12628 -9242 -6413 -9178
rect -6349 -9242 -6329 -9178
rect -12628 -9258 -6329 -9242
rect -12628 -9322 -6413 -9258
rect -6349 -9322 -6329 -9258
rect -12628 -9338 -6329 -9322
rect -12628 -9402 -6413 -9338
rect -6349 -9402 -6329 -9338
rect -12628 -9418 -6329 -9402
rect -12628 -9482 -6413 -9418
rect -6349 -9482 -6329 -9418
rect -12628 -9498 -6329 -9482
rect -12628 -9562 -6413 -9498
rect -6349 -9562 -6329 -9498
rect -12628 -9578 -6329 -9562
rect -12628 -9642 -6413 -9578
rect -6349 -9642 -6329 -9578
rect -12628 -9658 -6329 -9642
rect -12628 -9722 -6413 -9658
rect -6349 -9722 -6329 -9658
rect -12628 -9738 -6329 -9722
rect -12628 -9802 -6413 -9738
rect -6349 -9802 -6329 -9738
rect -12628 -9818 -6329 -9802
rect -12628 -9882 -6413 -9818
rect -6349 -9882 -6329 -9818
rect -12628 -9898 -6329 -9882
rect -12628 -9962 -6413 -9898
rect -6349 -9962 -6329 -9898
rect -12628 -9978 -6329 -9962
rect -12628 -10042 -6413 -9978
rect -6349 -10042 -6329 -9978
rect -12628 -10058 -6329 -10042
rect -12628 -10122 -6413 -10058
rect -6349 -10122 -6329 -10058
rect -12628 -10138 -6329 -10122
rect -12628 -10202 -6413 -10138
rect -6349 -10202 -6329 -10138
rect -12628 -10218 -6329 -10202
rect -12628 -10282 -6413 -10218
rect -6349 -10282 -6329 -10218
rect -12628 -10298 -6329 -10282
rect -12628 -10362 -6413 -10298
rect -6349 -10362 -6329 -10298
rect -12628 -10378 -6329 -10362
rect -12628 -10442 -6413 -10378
rect -6349 -10442 -6329 -10378
rect -12628 -10458 -6329 -10442
rect -12628 -10522 -6413 -10458
rect -6349 -10522 -6329 -10458
rect -12628 -10538 -6329 -10522
rect -12628 -10602 -6413 -10538
rect -6349 -10602 -6329 -10538
rect -12628 -10618 -6329 -10602
rect -12628 -10682 -6413 -10618
rect -6349 -10682 -6329 -10618
rect -12628 -10698 -6329 -10682
rect -12628 -10762 -6413 -10698
rect -6349 -10762 -6329 -10698
rect -12628 -10778 -6329 -10762
rect -12628 -10842 -6413 -10778
rect -6349 -10842 -6329 -10778
rect -12628 -10858 -6329 -10842
rect -12628 -10922 -6413 -10858
rect -6349 -10922 -6329 -10858
rect -12628 -10938 -6329 -10922
rect -12628 -11002 -6413 -10938
rect -6349 -11002 -6329 -10938
rect -12628 -11018 -6329 -11002
rect -12628 -11082 -6413 -11018
rect -6349 -11082 -6329 -11018
rect -12628 -11098 -6329 -11082
rect -12628 -11162 -6413 -11098
rect -6349 -11162 -6329 -11098
rect -12628 -11178 -6329 -11162
rect -12628 -11242 -6413 -11178
rect -6349 -11242 -6329 -11178
rect -12628 -11258 -6329 -11242
rect -12628 -11322 -6413 -11258
rect -6349 -11322 -6329 -11258
rect -12628 -11338 -6329 -11322
rect -12628 -11402 -6413 -11338
rect -6349 -11402 -6329 -11338
rect -12628 -11418 -6329 -11402
rect -12628 -11482 -6413 -11418
rect -6349 -11482 -6329 -11418
rect -12628 -11498 -6329 -11482
rect -12628 -11562 -6413 -11498
rect -6349 -11562 -6329 -11498
rect -12628 -11578 -6329 -11562
rect -12628 -11642 -6413 -11578
rect -6349 -11642 -6329 -11578
rect -12628 -11658 -6329 -11642
rect -12628 -11722 -6413 -11658
rect -6349 -11722 -6329 -11658
rect -12628 -11738 -6329 -11722
rect -12628 -11802 -6413 -11738
rect -6349 -11802 -6329 -11738
rect -12628 -11818 -6329 -11802
rect -12628 -11882 -6413 -11818
rect -6349 -11882 -6329 -11818
rect -12628 -11898 -6329 -11882
rect -12628 -11962 -6413 -11898
rect -6349 -11962 -6329 -11898
rect -12628 -11978 -6329 -11962
rect -12628 -12042 -6413 -11978
rect -6349 -12042 -6329 -11978
rect -12628 -12058 -6329 -12042
rect -12628 -12122 -6413 -12058
rect -6349 -12122 -6329 -12058
rect -12628 -12138 -6329 -12122
rect -12628 -12202 -6413 -12138
rect -6349 -12202 -6329 -12138
rect -12628 -12218 -6329 -12202
rect -12628 -12282 -6413 -12218
rect -6349 -12282 -6329 -12218
rect -12628 -12298 -6329 -12282
rect -12628 -12362 -6413 -12298
rect -6349 -12362 -6329 -12298
rect -12628 -12378 -6329 -12362
rect -12628 -12442 -6413 -12378
rect -6349 -12442 -6329 -12378
rect -12628 -12458 -6329 -12442
rect -12628 -12522 -6413 -12458
rect -6349 -12522 -6329 -12458
rect -12628 -12550 -6329 -12522
rect -6309 -6378 -10 -6350
rect -6309 -6442 -94 -6378
rect -30 -6442 -10 -6378
rect -6309 -6458 -10 -6442
rect -6309 -6522 -94 -6458
rect -30 -6522 -10 -6458
rect -6309 -6538 -10 -6522
rect -6309 -6602 -94 -6538
rect -30 -6602 -10 -6538
rect -6309 -6618 -10 -6602
rect -6309 -6682 -94 -6618
rect -30 -6682 -10 -6618
rect -6309 -6698 -10 -6682
rect -6309 -6762 -94 -6698
rect -30 -6762 -10 -6698
rect -6309 -6778 -10 -6762
rect -6309 -6842 -94 -6778
rect -30 -6842 -10 -6778
rect -6309 -6858 -10 -6842
rect -6309 -6922 -94 -6858
rect -30 -6922 -10 -6858
rect -6309 -6938 -10 -6922
rect -6309 -7002 -94 -6938
rect -30 -7002 -10 -6938
rect -6309 -7018 -10 -7002
rect -6309 -7082 -94 -7018
rect -30 -7082 -10 -7018
rect -6309 -7098 -10 -7082
rect -6309 -7162 -94 -7098
rect -30 -7162 -10 -7098
rect -6309 -7178 -10 -7162
rect -6309 -7242 -94 -7178
rect -30 -7242 -10 -7178
rect -6309 -7258 -10 -7242
rect -6309 -7322 -94 -7258
rect -30 -7322 -10 -7258
rect -6309 -7338 -10 -7322
rect -6309 -7402 -94 -7338
rect -30 -7402 -10 -7338
rect -6309 -7418 -10 -7402
rect -6309 -7482 -94 -7418
rect -30 -7482 -10 -7418
rect -6309 -7498 -10 -7482
rect -6309 -7562 -94 -7498
rect -30 -7562 -10 -7498
rect -6309 -7578 -10 -7562
rect -6309 -7642 -94 -7578
rect -30 -7642 -10 -7578
rect -6309 -7658 -10 -7642
rect -6309 -7722 -94 -7658
rect -30 -7722 -10 -7658
rect -6309 -7738 -10 -7722
rect -6309 -7802 -94 -7738
rect -30 -7802 -10 -7738
rect -6309 -7818 -10 -7802
rect -6309 -7882 -94 -7818
rect -30 -7882 -10 -7818
rect -6309 -7898 -10 -7882
rect -6309 -7962 -94 -7898
rect -30 -7962 -10 -7898
rect -6309 -7978 -10 -7962
rect -6309 -8042 -94 -7978
rect -30 -8042 -10 -7978
rect -6309 -8058 -10 -8042
rect -6309 -8122 -94 -8058
rect -30 -8122 -10 -8058
rect -6309 -8138 -10 -8122
rect -6309 -8202 -94 -8138
rect -30 -8202 -10 -8138
rect -6309 -8218 -10 -8202
rect -6309 -8282 -94 -8218
rect -30 -8282 -10 -8218
rect -6309 -8298 -10 -8282
rect -6309 -8362 -94 -8298
rect -30 -8362 -10 -8298
rect -6309 -8378 -10 -8362
rect -6309 -8442 -94 -8378
rect -30 -8442 -10 -8378
rect -6309 -8458 -10 -8442
rect -6309 -8522 -94 -8458
rect -30 -8522 -10 -8458
rect -6309 -8538 -10 -8522
rect -6309 -8602 -94 -8538
rect -30 -8602 -10 -8538
rect -6309 -8618 -10 -8602
rect -6309 -8682 -94 -8618
rect -30 -8682 -10 -8618
rect -6309 -8698 -10 -8682
rect -6309 -8762 -94 -8698
rect -30 -8762 -10 -8698
rect -6309 -8778 -10 -8762
rect -6309 -8842 -94 -8778
rect -30 -8842 -10 -8778
rect -6309 -8858 -10 -8842
rect -6309 -8922 -94 -8858
rect -30 -8922 -10 -8858
rect -6309 -8938 -10 -8922
rect -6309 -9002 -94 -8938
rect -30 -9002 -10 -8938
rect -6309 -9018 -10 -9002
rect -6309 -9082 -94 -9018
rect -30 -9082 -10 -9018
rect -6309 -9098 -10 -9082
rect -6309 -9162 -94 -9098
rect -30 -9162 -10 -9098
rect -6309 -9178 -10 -9162
rect -6309 -9242 -94 -9178
rect -30 -9242 -10 -9178
rect -6309 -9258 -10 -9242
rect -6309 -9322 -94 -9258
rect -30 -9322 -10 -9258
rect -6309 -9338 -10 -9322
rect -6309 -9402 -94 -9338
rect -30 -9402 -10 -9338
rect -6309 -9418 -10 -9402
rect -6309 -9482 -94 -9418
rect -30 -9482 -10 -9418
rect -6309 -9498 -10 -9482
rect -6309 -9562 -94 -9498
rect -30 -9562 -10 -9498
rect -6309 -9578 -10 -9562
rect -6309 -9642 -94 -9578
rect -30 -9642 -10 -9578
rect -6309 -9658 -10 -9642
rect -6309 -9722 -94 -9658
rect -30 -9722 -10 -9658
rect -6309 -9738 -10 -9722
rect -6309 -9802 -94 -9738
rect -30 -9802 -10 -9738
rect -6309 -9818 -10 -9802
rect -6309 -9882 -94 -9818
rect -30 -9882 -10 -9818
rect -6309 -9898 -10 -9882
rect -6309 -9962 -94 -9898
rect -30 -9962 -10 -9898
rect -6309 -9978 -10 -9962
rect -6309 -10042 -94 -9978
rect -30 -10042 -10 -9978
rect -6309 -10058 -10 -10042
rect -6309 -10122 -94 -10058
rect -30 -10122 -10 -10058
rect -6309 -10138 -10 -10122
rect -6309 -10202 -94 -10138
rect -30 -10202 -10 -10138
rect -6309 -10218 -10 -10202
rect -6309 -10282 -94 -10218
rect -30 -10282 -10 -10218
rect -6309 -10298 -10 -10282
rect -6309 -10362 -94 -10298
rect -30 -10362 -10 -10298
rect -6309 -10378 -10 -10362
rect -6309 -10442 -94 -10378
rect -30 -10442 -10 -10378
rect -6309 -10458 -10 -10442
rect -6309 -10522 -94 -10458
rect -30 -10522 -10 -10458
rect -6309 -10538 -10 -10522
rect -6309 -10602 -94 -10538
rect -30 -10602 -10 -10538
rect -6309 -10618 -10 -10602
rect -6309 -10682 -94 -10618
rect -30 -10682 -10 -10618
rect -6309 -10698 -10 -10682
rect -6309 -10762 -94 -10698
rect -30 -10762 -10 -10698
rect -6309 -10778 -10 -10762
rect -6309 -10842 -94 -10778
rect -30 -10842 -10 -10778
rect -6309 -10858 -10 -10842
rect -6309 -10922 -94 -10858
rect -30 -10922 -10 -10858
rect -6309 -10938 -10 -10922
rect -6309 -11002 -94 -10938
rect -30 -11002 -10 -10938
rect -6309 -11018 -10 -11002
rect -6309 -11082 -94 -11018
rect -30 -11082 -10 -11018
rect -6309 -11098 -10 -11082
rect -6309 -11162 -94 -11098
rect -30 -11162 -10 -11098
rect -6309 -11178 -10 -11162
rect -6309 -11242 -94 -11178
rect -30 -11242 -10 -11178
rect -6309 -11258 -10 -11242
rect -6309 -11322 -94 -11258
rect -30 -11322 -10 -11258
rect -6309 -11338 -10 -11322
rect -6309 -11402 -94 -11338
rect -30 -11402 -10 -11338
rect -6309 -11418 -10 -11402
rect -6309 -11482 -94 -11418
rect -30 -11482 -10 -11418
rect -6309 -11498 -10 -11482
rect -6309 -11562 -94 -11498
rect -30 -11562 -10 -11498
rect -6309 -11578 -10 -11562
rect -6309 -11642 -94 -11578
rect -30 -11642 -10 -11578
rect -6309 -11658 -10 -11642
rect -6309 -11722 -94 -11658
rect -30 -11722 -10 -11658
rect -6309 -11738 -10 -11722
rect -6309 -11802 -94 -11738
rect -30 -11802 -10 -11738
rect -6309 -11818 -10 -11802
rect -6309 -11882 -94 -11818
rect -30 -11882 -10 -11818
rect -6309 -11898 -10 -11882
rect -6309 -11962 -94 -11898
rect -30 -11962 -10 -11898
rect -6309 -11978 -10 -11962
rect -6309 -12042 -94 -11978
rect -30 -12042 -10 -11978
rect -6309 -12058 -10 -12042
rect -6309 -12122 -94 -12058
rect -30 -12122 -10 -12058
rect -6309 -12138 -10 -12122
rect -6309 -12202 -94 -12138
rect -30 -12202 -10 -12138
rect -6309 -12218 -10 -12202
rect -6309 -12282 -94 -12218
rect -30 -12282 -10 -12218
rect -6309 -12298 -10 -12282
rect -6309 -12362 -94 -12298
rect -30 -12362 -10 -12298
rect -6309 -12378 -10 -12362
rect -6309 -12442 -94 -12378
rect -30 -12442 -10 -12378
rect -6309 -12458 -10 -12442
rect -6309 -12522 -94 -12458
rect -30 -12522 -10 -12458
rect -6309 -12550 -10 -12522
rect 10 -6378 6309 -6350
rect 10 -6442 6225 -6378
rect 6289 -6442 6309 -6378
rect 10 -6458 6309 -6442
rect 10 -6522 6225 -6458
rect 6289 -6522 6309 -6458
rect 10 -6538 6309 -6522
rect 10 -6602 6225 -6538
rect 6289 -6602 6309 -6538
rect 10 -6618 6309 -6602
rect 10 -6682 6225 -6618
rect 6289 -6682 6309 -6618
rect 10 -6698 6309 -6682
rect 10 -6762 6225 -6698
rect 6289 -6762 6309 -6698
rect 10 -6778 6309 -6762
rect 10 -6842 6225 -6778
rect 6289 -6842 6309 -6778
rect 10 -6858 6309 -6842
rect 10 -6922 6225 -6858
rect 6289 -6922 6309 -6858
rect 10 -6938 6309 -6922
rect 10 -7002 6225 -6938
rect 6289 -7002 6309 -6938
rect 10 -7018 6309 -7002
rect 10 -7082 6225 -7018
rect 6289 -7082 6309 -7018
rect 10 -7098 6309 -7082
rect 10 -7162 6225 -7098
rect 6289 -7162 6309 -7098
rect 10 -7178 6309 -7162
rect 10 -7242 6225 -7178
rect 6289 -7242 6309 -7178
rect 10 -7258 6309 -7242
rect 10 -7322 6225 -7258
rect 6289 -7322 6309 -7258
rect 10 -7338 6309 -7322
rect 10 -7402 6225 -7338
rect 6289 -7402 6309 -7338
rect 10 -7418 6309 -7402
rect 10 -7482 6225 -7418
rect 6289 -7482 6309 -7418
rect 10 -7498 6309 -7482
rect 10 -7562 6225 -7498
rect 6289 -7562 6309 -7498
rect 10 -7578 6309 -7562
rect 10 -7642 6225 -7578
rect 6289 -7642 6309 -7578
rect 10 -7658 6309 -7642
rect 10 -7722 6225 -7658
rect 6289 -7722 6309 -7658
rect 10 -7738 6309 -7722
rect 10 -7802 6225 -7738
rect 6289 -7802 6309 -7738
rect 10 -7818 6309 -7802
rect 10 -7882 6225 -7818
rect 6289 -7882 6309 -7818
rect 10 -7898 6309 -7882
rect 10 -7962 6225 -7898
rect 6289 -7962 6309 -7898
rect 10 -7978 6309 -7962
rect 10 -8042 6225 -7978
rect 6289 -8042 6309 -7978
rect 10 -8058 6309 -8042
rect 10 -8122 6225 -8058
rect 6289 -8122 6309 -8058
rect 10 -8138 6309 -8122
rect 10 -8202 6225 -8138
rect 6289 -8202 6309 -8138
rect 10 -8218 6309 -8202
rect 10 -8282 6225 -8218
rect 6289 -8282 6309 -8218
rect 10 -8298 6309 -8282
rect 10 -8362 6225 -8298
rect 6289 -8362 6309 -8298
rect 10 -8378 6309 -8362
rect 10 -8442 6225 -8378
rect 6289 -8442 6309 -8378
rect 10 -8458 6309 -8442
rect 10 -8522 6225 -8458
rect 6289 -8522 6309 -8458
rect 10 -8538 6309 -8522
rect 10 -8602 6225 -8538
rect 6289 -8602 6309 -8538
rect 10 -8618 6309 -8602
rect 10 -8682 6225 -8618
rect 6289 -8682 6309 -8618
rect 10 -8698 6309 -8682
rect 10 -8762 6225 -8698
rect 6289 -8762 6309 -8698
rect 10 -8778 6309 -8762
rect 10 -8842 6225 -8778
rect 6289 -8842 6309 -8778
rect 10 -8858 6309 -8842
rect 10 -8922 6225 -8858
rect 6289 -8922 6309 -8858
rect 10 -8938 6309 -8922
rect 10 -9002 6225 -8938
rect 6289 -9002 6309 -8938
rect 10 -9018 6309 -9002
rect 10 -9082 6225 -9018
rect 6289 -9082 6309 -9018
rect 10 -9098 6309 -9082
rect 10 -9162 6225 -9098
rect 6289 -9162 6309 -9098
rect 10 -9178 6309 -9162
rect 10 -9242 6225 -9178
rect 6289 -9242 6309 -9178
rect 10 -9258 6309 -9242
rect 10 -9322 6225 -9258
rect 6289 -9322 6309 -9258
rect 10 -9338 6309 -9322
rect 10 -9402 6225 -9338
rect 6289 -9402 6309 -9338
rect 10 -9418 6309 -9402
rect 10 -9482 6225 -9418
rect 6289 -9482 6309 -9418
rect 10 -9498 6309 -9482
rect 10 -9562 6225 -9498
rect 6289 -9562 6309 -9498
rect 10 -9578 6309 -9562
rect 10 -9642 6225 -9578
rect 6289 -9642 6309 -9578
rect 10 -9658 6309 -9642
rect 10 -9722 6225 -9658
rect 6289 -9722 6309 -9658
rect 10 -9738 6309 -9722
rect 10 -9802 6225 -9738
rect 6289 -9802 6309 -9738
rect 10 -9818 6309 -9802
rect 10 -9882 6225 -9818
rect 6289 -9882 6309 -9818
rect 10 -9898 6309 -9882
rect 10 -9962 6225 -9898
rect 6289 -9962 6309 -9898
rect 10 -9978 6309 -9962
rect 10 -10042 6225 -9978
rect 6289 -10042 6309 -9978
rect 10 -10058 6309 -10042
rect 10 -10122 6225 -10058
rect 6289 -10122 6309 -10058
rect 10 -10138 6309 -10122
rect 10 -10202 6225 -10138
rect 6289 -10202 6309 -10138
rect 10 -10218 6309 -10202
rect 10 -10282 6225 -10218
rect 6289 -10282 6309 -10218
rect 10 -10298 6309 -10282
rect 10 -10362 6225 -10298
rect 6289 -10362 6309 -10298
rect 10 -10378 6309 -10362
rect 10 -10442 6225 -10378
rect 6289 -10442 6309 -10378
rect 10 -10458 6309 -10442
rect 10 -10522 6225 -10458
rect 6289 -10522 6309 -10458
rect 10 -10538 6309 -10522
rect 10 -10602 6225 -10538
rect 6289 -10602 6309 -10538
rect 10 -10618 6309 -10602
rect 10 -10682 6225 -10618
rect 6289 -10682 6309 -10618
rect 10 -10698 6309 -10682
rect 10 -10762 6225 -10698
rect 6289 -10762 6309 -10698
rect 10 -10778 6309 -10762
rect 10 -10842 6225 -10778
rect 6289 -10842 6309 -10778
rect 10 -10858 6309 -10842
rect 10 -10922 6225 -10858
rect 6289 -10922 6309 -10858
rect 10 -10938 6309 -10922
rect 10 -11002 6225 -10938
rect 6289 -11002 6309 -10938
rect 10 -11018 6309 -11002
rect 10 -11082 6225 -11018
rect 6289 -11082 6309 -11018
rect 10 -11098 6309 -11082
rect 10 -11162 6225 -11098
rect 6289 -11162 6309 -11098
rect 10 -11178 6309 -11162
rect 10 -11242 6225 -11178
rect 6289 -11242 6309 -11178
rect 10 -11258 6309 -11242
rect 10 -11322 6225 -11258
rect 6289 -11322 6309 -11258
rect 10 -11338 6309 -11322
rect 10 -11402 6225 -11338
rect 6289 -11402 6309 -11338
rect 10 -11418 6309 -11402
rect 10 -11482 6225 -11418
rect 6289 -11482 6309 -11418
rect 10 -11498 6309 -11482
rect 10 -11562 6225 -11498
rect 6289 -11562 6309 -11498
rect 10 -11578 6309 -11562
rect 10 -11642 6225 -11578
rect 6289 -11642 6309 -11578
rect 10 -11658 6309 -11642
rect 10 -11722 6225 -11658
rect 6289 -11722 6309 -11658
rect 10 -11738 6309 -11722
rect 10 -11802 6225 -11738
rect 6289 -11802 6309 -11738
rect 10 -11818 6309 -11802
rect 10 -11882 6225 -11818
rect 6289 -11882 6309 -11818
rect 10 -11898 6309 -11882
rect 10 -11962 6225 -11898
rect 6289 -11962 6309 -11898
rect 10 -11978 6309 -11962
rect 10 -12042 6225 -11978
rect 6289 -12042 6309 -11978
rect 10 -12058 6309 -12042
rect 10 -12122 6225 -12058
rect 6289 -12122 6309 -12058
rect 10 -12138 6309 -12122
rect 10 -12202 6225 -12138
rect 6289 -12202 6309 -12138
rect 10 -12218 6309 -12202
rect 10 -12282 6225 -12218
rect 6289 -12282 6309 -12218
rect 10 -12298 6309 -12282
rect 10 -12362 6225 -12298
rect 6289 -12362 6309 -12298
rect 10 -12378 6309 -12362
rect 10 -12442 6225 -12378
rect 6289 -12442 6309 -12378
rect 10 -12458 6309 -12442
rect 10 -12522 6225 -12458
rect 6289 -12522 6309 -12458
rect 10 -12550 6309 -12522
rect 6329 -6378 12628 -6350
rect 6329 -6442 12544 -6378
rect 12608 -6442 12628 -6378
rect 6329 -6458 12628 -6442
rect 6329 -6522 12544 -6458
rect 12608 -6522 12628 -6458
rect 6329 -6538 12628 -6522
rect 6329 -6602 12544 -6538
rect 12608 -6602 12628 -6538
rect 6329 -6618 12628 -6602
rect 6329 -6682 12544 -6618
rect 12608 -6682 12628 -6618
rect 6329 -6698 12628 -6682
rect 6329 -6762 12544 -6698
rect 12608 -6762 12628 -6698
rect 6329 -6778 12628 -6762
rect 6329 -6842 12544 -6778
rect 12608 -6842 12628 -6778
rect 6329 -6858 12628 -6842
rect 6329 -6922 12544 -6858
rect 12608 -6922 12628 -6858
rect 6329 -6938 12628 -6922
rect 6329 -7002 12544 -6938
rect 12608 -7002 12628 -6938
rect 6329 -7018 12628 -7002
rect 6329 -7082 12544 -7018
rect 12608 -7082 12628 -7018
rect 6329 -7098 12628 -7082
rect 6329 -7162 12544 -7098
rect 12608 -7162 12628 -7098
rect 6329 -7178 12628 -7162
rect 6329 -7242 12544 -7178
rect 12608 -7242 12628 -7178
rect 6329 -7258 12628 -7242
rect 6329 -7322 12544 -7258
rect 12608 -7322 12628 -7258
rect 6329 -7338 12628 -7322
rect 6329 -7402 12544 -7338
rect 12608 -7402 12628 -7338
rect 6329 -7418 12628 -7402
rect 6329 -7482 12544 -7418
rect 12608 -7482 12628 -7418
rect 6329 -7498 12628 -7482
rect 6329 -7562 12544 -7498
rect 12608 -7562 12628 -7498
rect 6329 -7578 12628 -7562
rect 6329 -7642 12544 -7578
rect 12608 -7642 12628 -7578
rect 6329 -7658 12628 -7642
rect 6329 -7722 12544 -7658
rect 12608 -7722 12628 -7658
rect 6329 -7738 12628 -7722
rect 6329 -7802 12544 -7738
rect 12608 -7802 12628 -7738
rect 6329 -7818 12628 -7802
rect 6329 -7882 12544 -7818
rect 12608 -7882 12628 -7818
rect 6329 -7898 12628 -7882
rect 6329 -7962 12544 -7898
rect 12608 -7962 12628 -7898
rect 6329 -7978 12628 -7962
rect 6329 -8042 12544 -7978
rect 12608 -8042 12628 -7978
rect 6329 -8058 12628 -8042
rect 6329 -8122 12544 -8058
rect 12608 -8122 12628 -8058
rect 6329 -8138 12628 -8122
rect 6329 -8202 12544 -8138
rect 12608 -8202 12628 -8138
rect 6329 -8218 12628 -8202
rect 6329 -8282 12544 -8218
rect 12608 -8282 12628 -8218
rect 6329 -8298 12628 -8282
rect 6329 -8362 12544 -8298
rect 12608 -8362 12628 -8298
rect 6329 -8378 12628 -8362
rect 6329 -8442 12544 -8378
rect 12608 -8442 12628 -8378
rect 6329 -8458 12628 -8442
rect 6329 -8522 12544 -8458
rect 12608 -8522 12628 -8458
rect 6329 -8538 12628 -8522
rect 6329 -8602 12544 -8538
rect 12608 -8602 12628 -8538
rect 6329 -8618 12628 -8602
rect 6329 -8682 12544 -8618
rect 12608 -8682 12628 -8618
rect 6329 -8698 12628 -8682
rect 6329 -8762 12544 -8698
rect 12608 -8762 12628 -8698
rect 6329 -8778 12628 -8762
rect 6329 -8842 12544 -8778
rect 12608 -8842 12628 -8778
rect 6329 -8858 12628 -8842
rect 6329 -8922 12544 -8858
rect 12608 -8922 12628 -8858
rect 6329 -8938 12628 -8922
rect 6329 -9002 12544 -8938
rect 12608 -9002 12628 -8938
rect 6329 -9018 12628 -9002
rect 6329 -9082 12544 -9018
rect 12608 -9082 12628 -9018
rect 6329 -9098 12628 -9082
rect 6329 -9162 12544 -9098
rect 12608 -9162 12628 -9098
rect 6329 -9178 12628 -9162
rect 6329 -9242 12544 -9178
rect 12608 -9242 12628 -9178
rect 6329 -9258 12628 -9242
rect 6329 -9322 12544 -9258
rect 12608 -9322 12628 -9258
rect 6329 -9338 12628 -9322
rect 6329 -9402 12544 -9338
rect 12608 -9402 12628 -9338
rect 6329 -9418 12628 -9402
rect 6329 -9482 12544 -9418
rect 12608 -9482 12628 -9418
rect 6329 -9498 12628 -9482
rect 6329 -9562 12544 -9498
rect 12608 -9562 12628 -9498
rect 6329 -9578 12628 -9562
rect 6329 -9642 12544 -9578
rect 12608 -9642 12628 -9578
rect 6329 -9658 12628 -9642
rect 6329 -9722 12544 -9658
rect 12608 -9722 12628 -9658
rect 6329 -9738 12628 -9722
rect 6329 -9802 12544 -9738
rect 12608 -9802 12628 -9738
rect 6329 -9818 12628 -9802
rect 6329 -9882 12544 -9818
rect 12608 -9882 12628 -9818
rect 6329 -9898 12628 -9882
rect 6329 -9962 12544 -9898
rect 12608 -9962 12628 -9898
rect 6329 -9978 12628 -9962
rect 6329 -10042 12544 -9978
rect 12608 -10042 12628 -9978
rect 6329 -10058 12628 -10042
rect 6329 -10122 12544 -10058
rect 12608 -10122 12628 -10058
rect 6329 -10138 12628 -10122
rect 6329 -10202 12544 -10138
rect 12608 -10202 12628 -10138
rect 6329 -10218 12628 -10202
rect 6329 -10282 12544 -10218
rect 12608 -10282 12628 -10218
rect 6329 -10298 12628 -10282
rect 6329 -10362 12544 -10298
rect 12608 -10362 12628 -10298
rect 6329 -10378 12628 -10362
rect 6329 -10442 12544 -10378
rect 12608 -10442 12628 -10378
rect 6329 -10458 12628 -10442
rect 6329 -10522 12544 -10458
rect 12608 -10522 12628 -10458
rect 6329 -10538 12628 -10522
rect 6329 -10602 12544 -10538
rect 12608 -10602 12628 -10538
rect 6329 -10618 12628 -10602
rect 6329 -10682 12544 -10618
rect 12608 -10682 12628 -10618
rect 6329 -10698 12628 -10682
rect 6329 -10762 12544 -10698
rect 12608 -10762 12628 -10698
rect 6329 -10778 12628 -10762
rect 6329 -10842 12544 -10778
rect 12608 -10842 12628 -10778
rect 6329 -10858 12628 -10842
rect 6329 -10922 12544 -10858
rect 12608 -10922 12628 -10858
rect 6329 -10938 12628 -10922
rect 6329 -11002 12544 -10938
rect 12608 -11002 12628 -10938
rect 6329 -11018 12628 -11002
rect 6329 -11082 12544 -11018
rect 12608 -11082 12628 -11018
rect 6329 -11098 12628 -11082
rect 6329 -11162 12544 -11098
rect 12608 -11162 12628 -11098
rect 6329 -11178 12628 -11162
rect 6329 -11242 12544 -11178
rect 12608 -11242 12628 -11178
rect 6329 -11258 12628 -11242
rect 6329 -11322 12544 -11258
rect 12608 -11322 12628 -11258
rect 6329 -11338 12628 -11322
rect 6329 -11402 12544 -11338
rect 12608 -11402 12628 -11338
rect 6329 -11418 12628 -11402
rect 6329 -11482 12544 -11418
rect 12608 -11482 12628 -11418
rect 6329 -11498 12628 -11482
rect 6329 -11562 12544 -11498
rect 12608 -11562 12628 -11498
rect 6329 -11578 12628 -11562
rect 6329 -11642 12544 -11578
rect 12608 -11642 12628 -11578
rect 6329 -11658 12628 -11642
rect 6329 -11722 12544 -11658
rect 12608 -11722 12628 -11658
rect 6329 -11738 12628 -11722
rect 6329 -11802 12544 -11738
rect 12608 -11802 12628 -11738
rect 6329 -11818 12628 -11802
rect 6329 -11882 12544 -11818
rect 12608 -11882 12628 -11818
rect 6329 -11898 12628 -11882
rect 6329 -11962 12544 -11898
rect 12608 -11962 12628 -11898
rect 6329 -11978 12628 -11962
rect 6329 -12042 12544 -11978
rect 12608 -12042 12628 -11978
rect 6329 -12058 12628 -12042
rect 6329 -12122 12544 -12058
rect 12608 -12122 12628 -12058
rect 6329 -12138 12628 -12122
rect 6329 -12202 12544 -12138
rect 12608 -12202 12628 -12138
rect 6329 -12218 12628 -12202
rect 6329 -12282 12544 -12218
rect 12608 -12282 12628 -12218
rect 6329 -12298 12628 -12282
rect 6329 -12362 12544 -12298
rect 12608 -12362 12628 -12298
rect 6329 -12378 12628 -12362
rect 6329 -12442 12544 -12378
rect 12608 -12442 12628 -12378
rect 6329 -12458 12628 -12442
rect 6329 -12522 12544 -12458
rect 12608 -12522 12628 -12458
rect 6329 -12550 12628 -12522
<< via3 >>
rect -6413 12458 -6349 12522
rect -6413 12378 -6349 12442
rect -6413 12298 -6349 12362
rect -6413 12218 -6349 12282
rect -6413 12138 -6349 12202
rect -6413 12058 -6349 12122
rect -6413 11978 -6349 12042
rect -6413 11898 -6349 11962
rect -6413 11818 -6349 11882
rect -6413 11738 -6349 11802
rect -6413 11658 -6349 11722
rect -6413 11578 -6349 11642
rect -6413 11498 -6349 11562
rect -6413 11418 -6349 11482
rect -6413 11338 -6349 11402
rect -6413 11258 -6349 11322
rect -6413 11178 -6349 11242
rect -6413 11098 -6349 11162
rect -6413 11018 -6349 11082
rect -6413 10938 -6349 11002
rect -6413 10858 -6349 10922
rect -6413 10778 -6349 10842
rect -6413 10698 -6349 10762
rect -6413 10618 -6349 10682
rect -6413 10538 -6349 10602
rect -6413 10458 -6349 10522
rect -6413 10378 -6349 10442
rect -6413 10298 -6349 10362
rect -6413 10218 -6349 10282
rect -6413 10138 -6349 10202
rect -6413 10058 -6349 10122
rect -6413 9978 -6349 10042
rect -6413 9898 -6349 9962
rect -6413 9818 -6349 9882
rect -6413 9738 -6349 9802
rect -6413 9658 -6349 9722
rect -6413 9578 -6349 9642
rect -6413 9498 -6349 9562
rect -6413 9418 -6349 9482
rect -6413 9338 -6349 9402
rect -6413 9258 -6349 9322
rect -6413 9178 -6349 9242
rect -6413 9098 -6349 9162
rect -6413 9018 -6349 9082
rect -6413 8938 -6349 9002
rect -6413 8858 -6349 8922
rect -6413 8778 -6349 8842
rect -6413 8698 -6349 8762
rect -6413 8618 -6349 8682
rect -6413 8538 -6349 8602
rect -6413 8458 -6349 8522
rect -6413 8378 -6349 8442
rect -6413 8298 -6349 8362
rect -6413 8218 -6349 8282
rect -6413 8138 -6349 8202
rect -6413 8058 -6349 8122
rect -6413 7978 -6349 8042
rect -6413 7898 -6349 7962
rect -6413 7818 -6349 7882
rect -6413 7738 -6349 7802
rect -6413 7658 -6349 7722
rect -6413 7578 -6349 7642
rect -6413 7498 -6349 7562
rect -6413 7418 -6349 7482
rect -6413 7338 -6349 7402
rect -6413 7258 -6349 7322
rect -6413 7178 -6349 7242
rect -6413 7098 -6349 7162
rect -6413 7018 -6349 7082
rect -6413 6938 -6349 7002
rect -6413 6858 -6349 6922
rect -6413 6778 -6349 6842
rect -6413 6698 -6349 6762
rect -6413 6618 -6349 6682
rect -6413 6538 -6349 6602
rect -6413 6458 -6349 6522
rect -6413 6378 -6349 6442
rect -94 12458 -30 12522
rect -94 12378 -30 12442
rect -94 12298 -30 12362
rect -94 12218 -30 12282
rect -94 12138 -30 12202
rect -94 12058 -30 12122
rect -94 11978 -30 12042
rect -94 11898 -30 11962
rect -94 11818 -30 11882
rect -94 11738 -30 11802
rect -94 11658 -30 11722
rect -94 11578 -30 11642
rect -94 11498 -30 11562
rect -94 11418 -30 11482
rect -94 11338 -30 11402
rect -94 11258 -30 11322
rect -94 11178 -30 11242
rect -94 11098 -30 11162
rect -94 11018 -30 11082
rect -94 10938 -30 11002
rect -94 10858 -30 10922
rect -94 10778 -30 10842
rect -94 10698 -30 10762
rect -94 10618 -30 10682
rect -94 10538 -30 10602
rect -94 10458 -30 10522
rect -94 10378 -30 10442
rect -94 10298 -30 10362
rect -94 10218 -30 10282
rect -94 10138 -30 10202
rect -94 10058 -30 10122
rect -94 9978 -30 10042
rect -94 9898 -30 9962
rect -94 9818 -30 9882
rect -94 9738 -30 9802
rect -94 9658 -30 9722
rect -94 9578 -30 9642
rect -94 9498 -30 9562
rect -94 9418 -30 9482
rect -94 9338 -30 9402
rect -94 9258 -30 9322
rect -94 9178 -30 9242
rect -94 9098 -30 9162
rect -94 9018 -30 9082
rect -94 8938 -30 9002
rect -94 8858 -30 8922
rect -94 8778 -30 8842
rect -94 8698 -30 8762
rect -94 8618 -30 8682
rect -94 8538 -30 8602
rect -94 8458 -30 8522
rect -94 8378 -30 8442
rect -94 8298 -30 8362
rect -94 8218 -30 8282
rect -94 8138 -30 8202
rect -94 8058 -30 8122
rect -94 7978 -30 8042
rect -94 7898 -30 7962
rect -94 7818 -30 7882
rect -94 7738 -30 7802
rect -94 7658 -30 7722
rect -94 7578 -30 7642
rect -94 7498 -30 7562
rect -94 7418 -30 7482
rect -94 7338 -30 7402
rect -94 7258 -30 7322
rect -94 7178 -30 7242
rect -94 7098 -30 7162
rect -94 7018 -30 7082
rect -94 6938 -30 7002
rect -94 6858 -30 6922
rect -94 6778 -30 6842
rect -94 6698 -30 6762
rect -94 6618 -30 6682
rect -94 6538 -30 6602
rect -94 6458 -30 6522
rect -94 6378 -30 6442
rect 6225 12458 6289 12522
rect 6225 12378 6289 12442
rect 6225 12298 6289 12362
rect 6225 12218 6289 12282
rect 6225 12138 6289 12202
rect 6225 12058 6289 12122
rect 6225 11978 6289 12042
rect 6225 11898 6289 11962
rect 6225 11818 6289 11882
rect 6225 11738 6289 11802
rect 6225 11658 6289 11722
rect 6225 11578 6289 11642
rect 6225 11498 6289 11562
rect 6225 11418 6289 11482
rect 6225 11338 6289 11402
rect 6225 11258 6289 11322
rect 6225 11178 6289 11242
rect 6225 11098 6289 11162
rect 6225 11018 6289 11082
rect 6225 10938 6289 11002
rect 6225 10858 6289 10922
rect 6225 10778 6289 10842
rect 6225 10698 6289 10762
rect 6225 10618 6289 10682
rect 6225 10538 6289 10602
rect 6225 10458 6289 10522
rect 6225 10378 6289 10442
rect 6225 10298 6289 10362
rect 6225 10218 6289 10282
rect 6225 10138 6289 10202
rect 6225 10058 6289 10122
rect 6225 9978 6289 10042
rect 6225 9898 6289 9962
rect 6225 9818 6289 9882
rect 6225 9738 6289 9802
rect 6225 9658 6289 9722
rect 6225 9578 6289 9642
rect 6225 9498 6289 9562
rect 6225 9418 6289 9482
rect 6225 9338 6289 9402
rect 6225 9258 6289 9322
rect 6225 9178 6289 9242
rect 6225 9098 6289 9162
rect 6225 9018 6289 9082
rect 6225 8938 6289 9002
rect 6225 8858 6289 8922
rect 6225 8778 6289 8842
rect 6225 8698 6289 8762
rect 6225 8618 6289 8682
rect 6225 8538 6289 8602
rect 6225 8458 6289 8522
rect 6225 8378 6289 8442
rect 6225 8298 6289 8362
rect 6225 8218 6289 8282
rect 6225 8138 6289 8202
rect 6225 8058 6289 8122
rect 6225 7978 6289 8042
rect 6225 7898 6289 7962
rect 6225 7818 6289 7882
rect 6225 7738 6289 7802
rect 6225 7658 6289 7722
rect 6225 7578 6289 7642
rect 6225 7498 6289 7562
rect 6225 7418 6289 7482
rect 6225 7338 6289 7402
rect 6225 7258 6289 7322
rect 6225 7178 6289 7242
rect 6225 7098 6289 7162
rect 6225 7018 6289 7082
rect 6225 6938 6289 7002
rect 6225 6858 6289 6922
rect 6225 6778 6289 6842
rect 6225 6698 6289 6762
rect 6225 6618 6289 6682
rect 6225 6538 6289 6602
rect 6225 6458 6289 6522
rect 6225 6378 6289 6442
rect 12544 12458 12608 12522
rect 12544 12378 12608 12442
rect 12544 12298 12608 12362
rect 12544 12218 12608 12282
rect 12544 12138 12608 12202
rect 12544 12058 12608 12122
rect 12544 11978 12608 12042
rect 12544 11898 12608 11962
rect 12544 11818 12608 11882
rect 12544 11738 12608 11802
rect 12544 11658 12608 11722
rect 12544 11578 12608 11642
rect 12544 11498 12608 11562
rect 12544 11418 12608 11482
rect 12544 11338 12608 11402
rect 12544 11258 12608 11322
rect 12544 11178 12608 11242
rect 12544 11098 12608 11162
rect 12544 11018 12608 11082
rect 12544 10938 12608 11002
rect 12544 10858 12608 10922
rect 12544 10778 12608 10842
rect 12544 10698 12608 10762
rect 12544 10618 12608 10682
rect 12544 10538 12608 10602
rect 12544 10458 12608 10522
rect 12544 10378 12608 10442
rect 12544 10298 12608 10362
rect 12544 10218 12608 10282
rect 12544 10138 12608 10202
rect 12544 10058 12608 10122
rect 12544 9978 12608 10042
rect 12544 9898 12608 9962
rect 12544 9818 12608 9882
rect 12544 9738 12608 9802
rect 12544 9658 12608 9722
rect 12544 9578 12608 9642
rect 12544 9498 12608 9562
rect 12544 9418 12608 9482
rect 12544 9338 12608 9402
rect 12544 9258 12608 9322
rect 12544 9178 12608 9242
rect 12544 9098 12608 9162
rect 12544 9018 12608 9082
rect 12544 8938 12608 9002
rect 12544 8858 12608 8922
rect 12544 8778 12608 8842
rect 12544 8698 12608 8762
rect 12544 8618 12608 8682
rect 12544 8538 12608 8602
rect 12544 8458 12608 8522
rect 12544 8378 12608 8442
rect 12544 8298 12608 8362
rect 12544 8218 12608 8282
rect 12544 8138 12608 8202
rect 12544 8058 12608 8122
rect 12544 7978 12608 8042
rect 12544 7898 12608 7962
rect 12544 7818 12608 7882
rect 12544 7738 12608 7802
rect 12544 7658 12608 7722
rect 12544 7578 12608 7642
rect 12544 7498 12608 7562
rect 12544 7418 12608 7482
rect 12544 7338 12608 7402
rect 12544 7258 12608 7322
rect 12544 7178 12608 7242
rect 12544 7098 12608 7162
rect 12544 7018 12608 7082
rect 12544 6938 12608 7002
rect 12544 6858 12608 6922
rect 12544 6778 12608 6842
rect 12544 6698 12608 6762
rect 12544 6618 12608 6682
rect 12544 6538 12608 6602
rect 12544 6458 12608 6522
rect 12544 6378 12608 6442
rect -6413 6158 -6349 6222
rect -6413 6078 -6349 6142
rect -6413 5998 -6349 6062
rect -6413 5918 -6349 5982
rect -6413 5838 -6349 5902
rect -6413 5758 -6349 5822
rect -6413 5678 -6349 5742
rect -6413 5598 -6349 5662
rect -6413 5518 -6349 5582
rect -6413 5438 -6349 5502
rect -6413 5358 -6349 5422
rect -6413 5278 -6349 5342
rect -6413 5198 -6349 5262
rect -6413 5118 -6349 5182
rect -6413 5038 -6349 5102
rect -6413 4958 -6349 5022
rect -6413 4878 -6349 4942
rect -6413 4798 -6349 4862
rect -6413 4718 -6349 4782
rect -6413 4638 -6349 4702
rect -6413 4558 -6349 4622
rect -6413 4478 -6349 4542
rect -6413 4398 -6349 4462
rect -6413 4318 -6349 4382
rect -6413 4238 -6349 4302
rect -6413 4158 -6349 4222
rect -6413 4078 -6349 4142
rect -6413 3998 -6349 4062
rect -6413 3918 -6349 3982
rect -6413 3838 -6349 3902
rect -6413 3758 -6349 3822
rect -6413 3678 -6349 3742
rect -6413 3598 -6349 3662
rect -6413 3518 -6349 3582
rect -6413 3438 -6349 3502
rect -6413 3358 -6349 3422
rect -6413 3278 -6349 3342
rect -6413 3198 -6349 3262
rect -6413 3118 -6349 3182
rect -6413 3038 -6349 3102
rect -6413 2958 -6349 3022
rect -6413 2878 -6349 2942
rect -6413 2798 -6349 2862
rect -6413 2718 -6349 2782
rect -6413 2638 -6349 2702
rect -6413 2558 -6349 2622
rect -6413 2478 -6349 2542
rect -6413 2398 -6349 2462
rect -6413 2318 -6349 2382
rect -6413 2238 -6349 2302
rect -6413 2158 -6349 2222
rect -6413 2078 -6349 2142
rect -6413 1998 -6349 2062
rect -6413 1918 -6349 1982
rect -6413 1838 -6349 1902
rect -6413 1758 -6349 1822
rect -6413 1678 -6349 1742
rect -6413 1598 -6349 1662
rect -6413 1518 -6349 1582
rect -6413 1438 -6349 1502
rect -6413 1358 -6349 1422
rect -6413 1278 -6349 1342
rect -6413 1198 -6349 1262
rect -6413 1118 -6349 1182
rect -6413 1038 -6349 1102
rect -6413 958 -6349 1022
rect -6413 878 -6349 942
rect -6413 798 -6349 862
rect -6413 718 -6349 782
rect -6413 638 -6349 702
rect -6413 558 -6349 622
rect -6413 478 -6349 542
rect -6413 398 -6349 462
rect -6413 318 -6349 382
rect -6413 238 -6349 302
rect -6413 158 -6349 222
rect -6413 78 -6349 142
rect -94 6158 -30 6222
rect -94 6078 -30 6142
rect -94 5998 -30 6062
rect -94 5918 -30 5982
rect -94 5838 -30 5902
rect -94 5758 -30 5822
rect -94 5678 -30 5742
rect -94 5598 -30 5662
rect -94 5518 -30 5582
rect -94 5438 -30 5502
rect -94 5358 -30 5422
rect -94 5278 -30 5342
rect -94 5198 -30 5262
rect -94 5118 -30 5182
rect -94 5038 -30 5102
rect -94 4958 -30 5022
rect -94 4878 -30 4942
rect -94 4798 -30 4862
rect -94 4718 -30 4782
rect -94 4638 -30 4702
rect -94 4558 -30 4622
rect -94 4478 -30 4542
rect -94 4398 -30 4462
rect -94 4318 -30 4382
rect -94 4238 -30 4302
rect -94 4158 -30 4222
rect -94 4078 -30 4142
rect -94 3998 -30 4062
rect -94 3918 -30 3982
rect -94 3838 -30 3902
rect -94 3758 -30 3822
rect -94 3678 -30 3742
rect -94 3598 -30 3662
rect -94 3518 -30 3582
rect -94 3438 -30 3502
rect -94 3358 -30 3422
rect -94 3278 -30 3342
rect -94 3198 -30 3262
rect -94 3118 -30 3182
rect -94 3038 -30 3102
rect -94 2958 -30 3022
rect -94 2878 -30 2942
rect -94 2798 -30 2862
rect -94 2718 -30 2782
rect -94 2638 -30 2702
rect -94 2558 -30 2622
rect -94 2478 -30 2542
rect -94 2398 -30 2462
rect -94 2318 -30 2382
rect -94 2238 -30 2302
rect -94 2158 -30 2222
rect -94 2078 -30 2142
rect -94 1998 -30 2062
rect -94 1918 -30 1982
rect -94 1838 -30 1902
rect -94 1758 -30 1822
rect -94 1678 -30 1742
rect -94 1598 -30 1662
rect -94 1518 -30 1582
rect -94 1438 -30 1502
rect -94 1358 -30 1422
rect -94 1278 -30 1342
rect -94 1198 -30 1262
rect -94 1118 -30 1182
rect -94 1038 -30 1102
rect -94 958 -30 1022
rect -94 878 -30 942
rect -94 798 -30 862
rect -94 718 -30 782
rect -94 638 -30 702
rect -94 558 -30 622
rect -94 478 -30 542
rect -94 398 -30 462
rect -94 318 -30 382
rect -94 238 -30 302
rect -94 158 -30 222
rect -94 78 -30 142
rect 6225 6158 6289 6222
rect 6225 6078 6289 6142
rect 6225 5998 6289 6062
rect 6225 5918 6289 5982
rect 6225 5838 6289 5902
rect 6225 5758 6289 5822
rect 6225 5678 6289 5742
rect 6225 5598 6289 5662
rect 6225 5518 6289 5582
rect 6225 5438 6289 5502
rect 6225 5358 6289 5422
rect 6225 5278 6289 5342
rect 6225 5198 6289 5262
rect 6225 5118 6289 5182
rect 6225 5038 6289 5102
rect 6225 4958 6289 5022
rect 6225 4878 6289 4942
rect 6225 4798 6289 4862
rect 6225 4718 6289 4782
rect 6225 4638 6289 4702
rect 6225 4558 6289 4622
rect 6225 4478 6289 4542
rect 6225 4398 6289 4462
rect 6225 4318 6289 4382
rect 6225 4238 6289 4302
rect 6225 4158 6289 4222
rect 6225 4078 6289 4142
rect 6225 3998 6289 4062
rect 6225 3918 6289 3982
rect 6225 3838 6289 3902
rect 6225 3758 6289 3822
rect 6225 3678 6289 3742
rect 6225 3598 6289 3662
rect 6225 3518 6289 3582
rect 6225 3438 6289 3502
rect 6225 3358 6289 3422
rect 6225 3278 6289 3342
rect 6225 3198 6289 3262
rect 6225 3118 6289 3182
rect 6225 3038 6289 3102
rect 6225 2958 6289 3022
rect 6225 2878 6289 2942
rect 6225 2798 6289 2862
rect 6225 2718 6289 2782
rect 6225 2638 6289 2702
rect 6225 2558 6289 2622
rect 6225 2478 6289 2542
rect 6225 2398 6289 2462
rect 6225 2318 6289 2382
rect 6225 2238 6289 2302
rect 6225 2158 6289 2222
rect 6225 2078 6289 2142
rect 6225 1998 6289 2062
rect 6225 1918 6289 1982
rect 6225 1838 6289 1902
rect 6225 1758 6289 1822
rect 6225 1678 6289 1742
rect 6225 1598 6289 1662
rect 6225 1518 6289 1582
rect 6225 1438 6289 1502
rect 6225 1358 6289 1422
rect 6225 1278 6289 1342
rect 6225 1198 6289 1262
rect 6225 1118 6289 1182
rect 6225 1038 6289 1102
rect 6225 958 6289 1022
rect 6225 878 6289 942
rect 6225 798 6289 862
rect 6225 718 6289 782
rect 6225 638 6289 702
rect 6225 558 6289 622
rect 6225 478 6289 542
rect 6225 398 6289 462
rect 6225 318 6289 382
rect 6225 238 6289 302
rect 6225 158 6289 222
rect 6225 78 6289 142
rect 12544 6158 12608 6222
rect 12544 6078 12608 6142
rect 12544 5998 12608 6062
rect 12544 5918 12608 5982
rect 12544 5838 12608 5902
rect 12544 5758 12608 5822
rect 12544 5678 12608 5742
rect 12544 5598 12608 5662
rect 12544 5518 12608 5582
rect 12544 5438 12608 5502
rect 12544 5358 12608 5422
rect 12544 5278 12608 5342
rect 12544 5198 12608 5262
rect 12544 5118 12608 5182
rect 12544 5038 12608 5102
rect 12544 4958 12608 5022
rect 12544 4878 12608 4942
rect 12544 4798 12608 4862
rect 12544 4718 12608 4782
rect 12544 4638 12608 4702
rect 12544 4558 12608 4622
rect 12544 4478 12608 4542
rect 12544 4398 12608 4462
rect 12544 4318 12608 4382
rect 12544 4238 12608 4302
rect 12544 4158 12608 4222
rect 12544 4078 12608 4142
rect 12544 3998 12608 4062
rect 12544 3918 12608 3982
rect 12544 3838 12608 3902
rect 12544 3758 12608 3822
rect 12544 3678 12608 3742
rect 12544 3598 12608 3662
rect 12544 3518 12608 3582
rect 12544 3438 12608 3502
rect 12544 3358 12608 3422
rect 12544 3278 12608 3342
rect 12544 3198 12608 3262
rect 12544 3118 12608 3182
rect 12544 3038 12608 3102
rect 12544 2958 12608 3022
rect 12544 2878 12608 2942
rect 12544 2798 12608 2862
rect 12544 2718 12608 2782
rect 12544 2638 12608 2702
rect 12544 2558 12608 2622
rect 12544 2478 12608 2542
rect 12544 2398 12608 2462
rect 12544 2318 12608 2382
rect 12544 2238 12608 2302
rect 12544 2158 12608 2222
rect 12544 2078 12608 2142
rect 12544 1998 12608 2062
rect 12544 1918 12608 1982
rect 12544 1838 12608 1902
rect 12544 1758 12608 1822
rect 12544 1678 12608 1742
rect 12544 1598 12608 1662
rect 12544 1518 12608 1582
rect 12544 1438 12608 1502
rect 12544 1358 12608 1422
rect 12544 1278 12608 1342
rect 12544 1198 12608 1262
rect 12544 1118 12608 1182
rect 12544 1038 12608 1102
rect 12544 958 12608 1022
rect 12544 878 12608 942
rect 12544 798 12608 862
rect 12544 718 12608 782
rect 12544 638 12608 702
rect 12544 558 12608 622
rect 12544 478 12608 542
rect 12544 398 12608 462
rect 12544 318 12608 382
rect 12544 238 12608 302
rect 12544 158 12608 222
rect 12544 78 12608 142
rect -6413 -142 -6349 -78
rect -6413 -222 -6349 -158
rect -6413 -302 -6349 -238
rect -6413 -382 -6349 -318
rect -6413 -462 -6349 -398
rect -6413 -542 -6349 -478
rect -6413 -622 -6349 -558
rect -6413 -702 -6349 -638
rect -6413 -782 -6349 -718
rect -6413 -862 -6349 -798
rect -6413 -942 -6349 -878
rect -6413 -1022 -6349 -958
rect -6413 -1102 -6349 -1038
rect -6413 -1182 -6349 -1118
rect -6413 -1262 -6349 -1198
rect -6413 -1342 -6349 -1278
rect -6413 -1422 -6349 -1358
rect -6413 -1502 -6349 -1438
rect -6413 -1582 -6349 -1518
rect -6413 -1662 -6349 -1598
rect -6413 -1742 -6349 -1678
rect -6413 -1822 -6349 -1758
rect -6413 -1902 -6349 -1838
rect -6413 -1982 -6349 -1918
rect -6413 -2062 -6349 -1998
rect -6413 -2142 -6349 -2078
rect -6413 -2222 -6349 -2158
rect -6413 -2302 -6349 -2238
rect -6413 -2382 -6349 -2318
rect -6413 -2462 -6349 -2398
rect -6413 -2542 -6349 -2478
rect -6413 -2622 -6349 -2558
rect -6413 -2702 -6349 -2638
rect -6413 -2782 -6349 -2718
rect -6413 -2862 -6349 -2798
rect -6413 -2942 -6349 -2878
rect -6413 -3022 -6349 -2958
rect -6413 -3102 -6349 -3038
rect -6413 -3182 -6349 -3118
rect -6413 -3262 -6349 -3198
rect -6413 -3342 -6349 -3278
rect -6413 -3422 -6349 -3358
rect -6413 -3502 -6349 -3438
rect -6413 -3582 -6349 -3518
rect -6413 -3662 -6349 -3598
rect -6413 -3742 -6349 -3678
rect -6413 -3822 -6349 -3758
rect -6413 -3902 -6349 -3838
rect -6413 -3982 -6349 -3918
rect -6413 -4062 -6349 -3998
rect -6413 -4142 -6349 -4078
rect -6413 -4222 -6349 -4158
rect -6413 -4302 -6349 -4238
rect -6413 -4382 -6349 -4318
rect -6413 -4462 -6349 -4398
rect -6413 -4542 -6349 -4478
rect -6413 -4622 -6349 -4558
rect -6413 -4702 -6349 -4638
rect -6413 -4782 -6349 -4718
rect -6413 -4862 -6349 -4798
rect -6413 -4942 -6349 -4878
rect -6413 -5022 -6349 -4958
rect -6413 -5102 -6349 -5038
rect -6413 -5182 -6349 -5118
rect -6413 -5262 -6349 -5198
rect -6413 -5342 -6349 -5278
rect -6413 -5422 -6349 -5358
rect -6413 -5502 -6349 -5438
rect -6413 -5582 -6349 -5518
rect -6413 -5662 -6349 -5598
rect -6413 -5742 -6349 -5678
rect -6413 -5822 -6349 -5758
rect -6413 -5902 -6349 -5838
rect -6413 -5982 -6349 -5918
rect -6413 -6062 -6349 -5998
rect -6413 -6142 -6349 -6078
rect -6413 -6222 -6349 -6158
rect -94 -142 -30 -78
rect -94 -222 -30 -158
rect -94 -302 -30 -238
rect -94 -382 -30 -318
rect -94 -462 -30 -398
rect -94 -542 -30 -478
rect -94 -622 -30 -558
rect -94 -702 -30 -638
rect -94 -782 -30 -718
rect -94 -862 -30 -798
rect -94 -942 -30 -878
rect -94 -1022 -30 -958
rect -94 -1102 -30 -1038
rect -94 -1182 -30 -1118
rect -94 -1262 -30 -1198
rect -94 -1342 -30 -1278
rect -94 -1422 -30 -1358
rect -94 -1502 -30 -1438
rect -94 -1582 -30 -1518
rect -94 -1662 -30 -1598
rect -94 -1742 -30 -1678
rect -94 -1822 -30 -1758
rect -94 -1902 -30 -1838
rect -94 -1982 -30 -1918
rect -94 -2062 -30 -1998
rect -94 -2142 -30 -2078
rect -94 -2222 -30 -2158
rect -94 -2302 -30 -2238
rect -94 -2382 -30 -2318
rect -94 -2462 -30 -2398
rect -94 -2542 -30 -2478
rect -94 -2622 -30 -2558
rect -94 -2702 -30 -2638
rect -94 -2782 -30 -2718
rect -94 -2862 -30 -2798
rect -94 -2942 -30 -2878
rect -94 -3022 -30 -2958
rect -94 -3102 -30 -3038
rect -94 -3182 -30 -3118
rect -94 -3262 -30 -3198
rect -94 -3342 -30 -3278
rect -94 -3422 -30 -3358
rect -94 -3502 -30 -3438
rect -94 -3582 -30 -3518
rect -94 -3662 -30 -3598
rect -94 -3742 -30 -3678
rect -94 -3822 -30 -3758
rect -94 -3902 -30 -3838
rect -94 -3982 -30 -3918
rect -94 -4062 -30 -3998
rect -94 -4142 -30 -4078
rect -94 -4222 -30 -4158
rect -94 -4302 -30 -4238
rect -94 -4382 -30 -4318
rect -94 -4462 -30 -4398
rect -94 -4542 -30 -4478
rect -94 -4622 -30 -4558
rect -94 -4702 -30 -4638
rect -94 -4782 -30 -4718
rect -94 -4862 -30 -4798
rect -94 -4942 -30 -4878
rect -94 -5022 -30 -4958
rect -94 -5102 -30 -5038
rect -94 -5182 -30 -5118
rect -94 -5262 -30 -5198
rect -94 -5342 -30 -5278
rect -94 -5422 -30 -5358
rect -94 -5502 -30 -5438
rect -94 -5582 -30 -5518
rect -94 -5662 -30 -5598
rect -94 -5742 -30 -5678
rect -94 -5822 -30 -5758
rect -94 -5902 -30 -5838
rect -94 -5982 -30 -5918
rect -94 -6062 -30 -5998
rect -94 -6142 -30 -6078
rect -94 -6222 -30 -6158
rect 6225 -142 6289 -78
rect 6225 -222 6289 -158
rect 6225 -302 6289 -238
rect 6225 -382 6289 -318
rect 6225 -462 6289 -398
rect 6225 -542 6289 -478
rect 6225 -622 6289 -558
rect 6225 -702 6289 -638
rect 6225 -782 6289 -718
rect 6225 -862 6289 -798
rect 6225 -942 6289 -878
rect 6225 -1022 6289 -958
rect 6225 -1102 6289 -1038
rect 6225 -1182 6289 -1118
rect 6225 -1262 6289 -1198
rect 6225 -1342 6289 -1278
rect 6225 -1422 6289 -1358
rect 6225 -1502 6289 -1438
rect 6225 -1582 6289 -1518
rect 6225 -1662 6289 -1598
rect 6225 -1742 6289 -1678
rect 6225 -1822 6289 -1758
rect 6225 -1902 6289 -1838
rect 6225 -1982 6289 -1918
rect 6225 -2062 6289 -1998
rect 6225 -2142 6289 -2078
rect 6225 -2222 6289 -2158
rect 6225 -2302 6289 -2238
rect 6225 -2382 6289 -2318
rect 6225 -2462 6289 -2398
rect 6225 -2542 6289 -2478
rect 6225 -2622 6289 -2558
rect 6225 -2702 6289 -2638
rect 6225 -2782 6289 -2718
rect 6225 -2862 6289 -2798
rect 6225 -2942 6289 -2878
rect 6225 -3022 6289 -2958
rect 6225 -3102 6289 -3038
rect 6225 -3182 6289 -3118
rect 6225 -3262 6289 -3198
rect 6225 -3342 6289 -3278
rect 6225 -3422 6289 -3358
rect 6225 -3502 6289 -3438
rect 6225 -3582 6289 -3518
rect 6225 -3662 6289 -3598
rect 6225 -3742 6289 -3678
rect 6225 -3822 6289 -3758
rect 6225 -3902 6289 -3838
rect 6225 -3982 6289 -3918
rect 6225 -4062 6289 -3998
rect 6225 -4142 6289 -4078
rect 6225 -4222 6289 -4158
rect 6225 -4302 6289 -4238
rect 6225 -4382 6289 -4318
rect 6225 -4462 6289 -4398
rect 6225 -4542 6289 -4478
rect 6225 -4622 6289 -4558
rect 6225 -4702 6289 -4638
rect 6225 -4782 6289 -4718
rect 6225 -4862 6289 -4798
rect 6225 -4942 6289 -4878
rect 6225 -5022 6289 -4958
rect 6225 -5102 6289 -5038
rect 6225 -5182 6289 -5118
rect 6225 -5262 6289 -5198
rect 6225 -5342 6289 -5278
rect 6225 -5422 6289 -5358
rect 6225 -5502 6289 -5438
rect 6225 -5582 6289 -5518
rect 6225 -5662 6289 -5598
rect 6225 -5742 6289 -5678
rect 6225 -5822 6289 -5758
rect 6225 -5902 6289 -5838
rect 6225 -5982 6289 -5918
rect 6225 -6062 6289 -5998
rect 6225 -6142 6289 -6078
rect 6225 -6222 6289 -6158
rect 12544 -142 12608 -78
rect 12544 -222 12608 -158
rect 12544 -302 12608 -238
rect 12544 -382 12608 -318
rect 12544 -462 12608 -398
rect 12544 -542 12608 -478
rect 12544 -622 12608 -558
rect 12544 -702 12608 -638
rect 12544 -782 12608 -718
rect 12544 -862 12608 -798
rect 12544 -942 12608 -878
rect 12544 -1022 12608 -958
rect 12544 -1102 12608 -1038
rect 12544 -1182 12608 -1118
rect 12544 -1262 12608 -1198
rect 12544 -1342 12608 -1278
rect 12544 -1422 12608 -1358
rect 12544 -1502 12608 -1438
rect 12544 -1582 12608 -1518
rect 12544 -1662 12608 -1598
rect 12544 -1742 12608 -1678
rect 12544 -1822 12608 -1758
rect 12544 -1902 12608 -1838
rect 12544 -1982 12608 -1918
rect 12544 -2062 12608 -1998
rect 12544 -2142 12608 -2078
rect 12544 -2222 12608 -2158
rect 12544 -2302 12608 -2238
rect 12544 -2382 12608 -2318
rect 12544 -2462 12608 -2398
rect 12544 -2542 12608 -2478
rect 12544 -2622 12608 -2558
rect 12544 -2702 12608 -2638
rect 12544 -2782 12608 -2718
rect 12544 -2862 12608 -2798
rect 12544 -2942 12608 -2878
rect 12544 -3022 12608 -2958
rect 12544 -3102 12608 -3038
rect 12544 -3182 12608 -3118
rect 12544 -3262 12608 -3198
rect 12544 -3342 12608 -3278
rect 12544 -3422 12608 -3358
rect 12544 -3502 12608 -3438
rect 12544 -3582 12608 -3518
rect 12544 -3662 12608 -3598
rect 12544 -3742 12608 -3678
rect 12544 -3822 12608 -3758
rect 12544 -3902 12608 -3838
rect 12544 -3982 12608 -3918
rect 12544 -4062 12608 -3998
rect 12544 -4142 12608 -4078
rect 12544 -4222 12608 -4158
rect 12544 -4302 12608 -4238
rect 12544 -4382 12608 -4318
rect 12544 -4462 12608 -4398
rect 12544 -4542 12608 -4478
rect 12544 -4622 12608 -4558
rect 12544 -4702 12608 -4638
rect 12544 -4782 12608 -4718
rect 12544 -4862 12608 -4798
rect 12544 -4942 12608 -4878
rect 12544 -5022 12608 -4958
rect 12544 -5102 12608 -5038
rect 12544 -5182 12608 -5118
rect 12544 -5262 12608 -5198
rect 12544 -5342 12608 -5278
rect 12544 -5422 12608 -5358
rect 12544 -5502 12608 -5438
rect 12544 -5582 12608 -5518
rect 12544 -5662 12608 -5598
rect 12544 -5742 12608 -5678
rect 12544 -5822 12608 -5758
rect 12544 -5902 12608 -5838
rect 12544 -5982 12608 -5918
rect 12544 -6062 12608 -5998
rect 12544 -6142 12608 -6078
rect 12544 -6222 12608 -6158
rect -6413 -6442 -6349 -6378
rect -6413 -6522 -6349 -6458
rect -6413 -6602 -6349 -6538
rect -6413 -6682 -6349 -6618
rect -6413 -6762 -6349 -6698
rect -6413 -6842 -6349 -6778
rect -6413 -6922 -6349 -6858
rect -6413 -7002 -6349 -6938
rect -6413 -7082 -6349 -7018
rect -6413 -7162 -6349 -7098
rect -6413 -7242 -6349 -7178
rect -6413 -7322 -6349 -7258
rect -6413 -7402 -6349 -7338
rect -6413 -7482 -6349 -7418
rect -6413 -7562 -6349 -7498
rect -6413 -7642 -6349 -7578
rect -6413 -7722 -6349 -7658
rect -6413 -7802 -6349 -7738
rect -6413 -7882 -6349 -7818
rect -6413 -7962 -6349 -7898
rect -6413 -8042 -6349 -7978
rect -6413 -8122 -6349 -8058
rect -6413 -8202 -6349 -8138
rect -6413 -8282 -6349 -8218
rect -6413 -8362 -6349 -8298
rect -6413 -8442 -6349 -8378
rect -6413 -8522 -6349 -8458
rect -6413 -8602 -6349 -8538
rect -6413 -8682 -6349 -8618
rect -6413 -8762 -6349 -8698
rect -6413 -8842 -6349 -8778
rect -6413 -8922 -6349 -8858
rect -6413 -9002 -6349 -8938
rect -6413 -9082 -6349 -9018
rect -6413 -9162 -6349 -9098
rect -6413 -9242 -6349 -9178
rect -6413 -9322 -6349 -9258
rect -6413 -9402 -6349 -9338
rect -6413 -9482 -6349 -9418
rect -6413 -9562 -6349 -9498
rect -6413 -9642 -6349 -9578
rect -6413 -9722 -6349 -9658
rect -6413 -9802 -6349 -9738
rect -6413 -9882 -6349 -9818
rect -6413 -9962 -6349 -9898
rect -6413 -10042 -6349 -9978
rect -6413 -10122 -6349 -10058
rect -6413 -10202 -6349 -10138
rect -6413 -10282 -6349 -10218
rect -6413 -10362 -6349 -10298
rect -6413 -10442 -6349 -10378
rect -6413 -10522 -6349 -10458
rect -6413 -10602 -6349 -10538
rect -6413 -10682 -6349 -10618
rect -6413 -10762 -6349 -10698
rect -6413 -10842 -6349 -10778
rect -6413 -10922 -6349 -10858
rect -6413 -11002 -6349 -10938
rect -6413 -11082 -6349 -11018
rect -6413 -11162 -6349 -11098
rect -6413 -11242 -6349 -11178
rect -6413 -11322 -6349 -11258
rect -6413 -11402 -6349 -11338
rect -6413 -11482 -6349 -11418
rect -6413 -11562 -6349 -11498
rect -6413 -11642 -6349 -11578
rect -6413 -11722 -6349 -11658
rect -6413 -11802 -6349 -11738
rect -6413 -11882 -6349 -11818
rect -6413 -11962 -6349 -11898
rect -6413 -12042 -6349 -11978
rect -6413 -12122 -6349 -12058
rect -6413 -12202 -6349 -12138
rect -6413 -12282 -6349 -12218
rect -6413 -12362 -6349 -12298
rect -6413 -12442 -6349 -12378
rect -6413 -12522 -6349 -12458
rect -94 -6442 -30 -6378
rect -94 -6522 -30 -6458
rect -94 -6602 -30 -6538
rect -94 -6682 -30 -6618
rect -94 -6762 -30 -6698
rect -94 -6842 -30 -6778
rect -94 -6922 -30 -6858
rect -94 -7002 -30 -6938
rect -94 -7082 -30 -7018
rect -94 -7162 -30 -7098
rect -94 -7242 -30 -7178
rect -94 -7322 -30 -7258
rect -94 -7402 -30 -7338
rect -94 -7482 -30 -7418
rect -94 -7562 -30 -7498
rect -94 -7642 -30 -7578
rect -94 -7722 -30 -7658
rect -94 -7802 -30 -7738
rect -94 -7882 -30 -7818
rect -94 -7962 -30 -7898
rect -94 -8042 -30 -7978
rect -94 -8122 -30 -8058
rect -94 -8202 -30 -8138
rect -94 -8282 -30 -8218
rect -94 -8362 -30 -8298
rect -94 -8442 -30 -8378
rect -94 -8522 -30 -8458
rect -94 -8602 -30 -8538
rect -94 -8682 -30 -8618
rect -94 -8762 -30 -8698
rect -94 -8842 -30 -8778
rect -94 -8922 -30 -8858
rect -94 -9002 -30 -8938
rect -94 -9082 -30 -9018
rect -94 -9162 -30 -9098
rect -94 -9242 -30 -9178
rect -94 -9322 -30 -9258
rect -94 -9402 -30 -9338
rect -94 -9482 -30 -9418
rect -94 -9562 -30 -9498
rect -94 -9642 -30 -9578
rect -94 -9722 -30 -9658
rect -94 -9802 -30 -9738
rect -94 -9882 -30 -9818
rect -94 -9962 -30 -9898
rect -94 -10042 -30 -9978
rect -94 -10122 -30 -10058
rect -94 -10202 -30 -10138
rect -94 -10282 -30 -10218
rect -94 -10362 -30 -10298
rect -94 -10442 -30 -10378
rect -94 -10522 -30 -10458
rect -94 -10602 -30 -10538
rect -94 -10682 -30 -10618
rect -94 -10762 -30 -10698
rect -94 -10842 -30 -10778
rect -94 -10922 -30 -10858
rect -94 -11002 -30 -10938
rect -94 -11082 -30 -11018
rect -94 -11162 -30 -11098
rect -94 -11242 -30 -11178
rect -94 -11322 -30 -11258
rect -94 -11402 -30 -11338
rect -94 -11482 -30 -11418
rect -94 -11562 -30 -11498
rect -94 -11642 -30 -11578
rect -94 -11722 -30 -11658
rect -94 -11802 -30 -11738
rect -94 -11882 -30 -11818
rect -94 -11962 -30 -11898
rect -94 -12042 -30 -11978
rect -94 -12122 -30 -12058
rect -94 -12202 -30 -12138
rect -94 -12282 -30 -12218
rect -94 -12362 -30 -12298
rect -94 -12442 -30 -12378
rect -94 -12522 -30 -12458
rect 6225 -6442 6289 -6378
rect 6225 -6522 6289 -6458
rect 6225 -6602 6289 -6538
rect 6225 -6682 6289 -6618
rect 6225 -6762 6289 -6698
rect 6225 -6842 6289 -6778
rect 6225 -6922 6289 -6858
rect 6225 -7002 6289 -6938
rect 6225 -7082 6289 -7018
rect 6225 -7162 6289 -7098
rect 6225 -7242 6289 -7178
rect 6225 -7322 6289 -7258
rect 6225 -7402 6289 -7338
rect 6225 -7482 6289 -7418
rect 6225 -7562 6289 -7498
rect 6225 -7642 6289 -7578
rect 6225 -7722 6289 -7658
rect 6225 -7802 6289 -7738
rect 6225 -7882 6289 -7818
rect 6225 -7962 6289 -7898
rect 6225 -8042 6289 -7978
rect 6225 -8122 6289 -8058
rect 6225 -8202 6289 -8138
rect 6225 -8282 6289 -8218
rect 6225 -8362 6289 -8298
rect 6225 -8442 6289 -8378
rect 6225 -8522 6289 -8458
rect 6225 -8602 6289 -8538
rect 6225 -8682 6289 -8618
rect 6225 -8762 6289 -8698
rect 6225 -8842 6289 -8778
rect 6225 -8922 6289 -8858
rect 6225 -9002 6289 -8938
rect 6225 -9082 6289 -9018
rect 6225 -9162 6289 -9098
rect 6225 -9242 6289 -9178
rect 6225 -9322 6289 -9258
rect 6225 -9402 6289 -9338
rect 6225 -9482 6289 -9418
rect 6225 -9562 6289 -9498
rect 6225 -9642 6289 -9578
rect 6225 -9722 6289 -9658
rect 6225 -9802 6289 -9738
rect 6225 -9882 6289 -9818
rect 6225 -9962 6289 -9898
rect 6225 -10042 6289 -9978
rect 6225 -10122 6289 -10058
rect 6225 -10202 6289 -10138
rect 6225 -10282 6289 -10218
rect 6225 -10362 6289 -10298
rect 6225 -10442 6289 -10378
rect 6225 -10522 6289 -10458
rect 6225 -10602 6289 -10538
rect 6225 -10682 6289 -10618
rect 6225 -10762 6289 -10698
rect 6225 -10842 6289 -10778
rect 6225 -10922 6289 -10858
rect 6225 -11002 6289 -10938
rect 6225 -11082 6289 -11018
rect 6225 -11162 6289 -11098
rect 6225 -11242 6289 -11178
rect 6225 -11322 6289 -11258
rect 6225 -11402 6289 -11338
rect 6225 -11482 6289 -11418
rect 6225 -11562 6289 -11498
rect 6225 -11642 6289 -11578
rect 6225 -11722 6289 -11658
rect 6225 -11802 6289 -11738
rect 6225 -11882 6289 -11818
rect 6225 -11962 6289 -11898
rect 6225 -12042 6289 -11978
rect 6225 -12122 6289 -12058
rect 6225 -12202 6289 -12138
rect 6225 -12282 6289 -12218
rect 6225 -12362 6289 -12298
rect 6225 -12442 6289 -12378
rect 6225 -12522 6289 -12458
rect 12544 -6442 12608 -6378
rect 12544 -6522 12608 -6458
rect 12544 -6602 12608 -6538
rect 12544 -6682 12608 -6618
rect 12544 -6762 12608 -6698
rect 12544 -6842 12608 -6778
rect 12544 -6922 12608 -6858
rect 12544 -7002 12608 -6938
rect 12544 -7082 12608 -7018
rect 12544 -7162 12608 -7098
rect 12544 -7242 12608 -7178
rect 12544 -7322 12608 -7258
rect 12544 -7402 12608 -7338
rect 12544 -7482 12608 -7418
rect 12544 -7562 12608 -7498
rect 12544 -7642 12608 -7578
rect 12544 -7722 12608 -7658
rect 12544 -7802 12608 -7738
rect 12544 -7882 12608 -7818
rect 12544 -7962 12608 -7898
rect 12544 -8042 12608 -7978
rect 12544 -8122 12608 -8058
rect 12544 -8202 12608 -8138
rect 12544 -8282 12608 -8218
rect 12544 -8362 12608 -8298
rect 12544 -8442 12608 -8378
rect 12544 -8522 12608 -8458
rect 12544 -8602 12608 -8538
rect 12544 -8682 12608 -8618
rect 12544 -8762 12608 -8698
rect 12544 -8842 12608 -8778
rect 12544 -8922 12608 -8858
rect 12544 -9002 12608 -8938
rect 12544 -9082 12608 -9018
rect 12544 -9162 12608 -9098
rect 12544 -9242 12608 -9178
rect 12544 -9322 12608 -9258
rect 12544 -9402 12608 -9338
rect 12544 -9482 12608 -9418
rect 12544 -9562 12608 -9498
rect 12544 -9642 12608 -9578
rect 12544 -9722 12608 -9658
rect 12544 -9802 12608 -9738
rect 12544 -9882 12608 -9818
rect 12544 -9962 12608 -9898
rect 12544 -10042 12608 -9978
rect 12544 -10122 12608 -10058
rect 12544 -10202 12608 -10138
rect 12544 -10282 12608 -10218
rect 12544 -10362 12608 -10298
rect 12544 -10442 12608 -10378
rect 12544 -10522 12608 -10458
rect 12544 -10602 12608 -10538
rect 12544 -10682 12608 -10618
rect 12544 -10762 12608 -10698
rect 12544 -10842 12608 -10778
rect 12544 -10922 12608 -10858
rect 12544 -11002 12608 -10938
rect 12544 -11082 12608 -11018
rect 12544 -11162 12608 -11098
rect 12544 -11242 12608 -11178
rect 12544 -11322 12608 -11258
rect 12544 -11402 12608 -11338
rect 12544 -11482 12608 -11418
rect 12544 -11562 12608 -11498
rect 12544 -11642 12608 -11578
rect 12544 -11722 12608 -11658
rect 12544 -11802 12608 -11738
rect 12544 -11882 12608 -11818
rect 12544 -11962 12608 -11898
rect 12544 -12042 12608 -11978
rect 12544 -12122 12608 -12058
rect 12544 -12202 12608 -12138
rect 12544 -12282 12608 -12218
rect 12544 -12362 12608 -12298
rect 12544 -12442 12608 -12378
rect 12544 -12522 12608 -12458
<< mimcap >>
rect -12528 12402 -6528 12450
rect -12528 6498 -12480 12402
rect -6576 6498 -6528 12402
rect -12528 6450 -6528 6498
rect -6209 12402 -209 12450
rect -6209 6498 -6161 12402
rect -257 6498 -209 12402
rect -6209 6450 -209 6498
rect 110 12402 6110 12450
rect 110 6498 158 12402
rect 6062 6498 6110 12402
rect 110 6450 6110 6498
rect 6429 12402 12429 12450
rect 6429 6498 6477 12402
rect 12381 6498 12429 12402
rect 6429 6450 12429 6498
rect -12528 6102 -6528 6150
rect -12528 198 -12480 6102
rect -6576 198 -6528 6102
rect -12528 150 -6528 198
rect -6209 6102 -209 6150
rect -6209 198 -6161 6102
rect -257 198 -209 6102
rect -6209 150 -209 198
rect 110 6102 6110 6150
rect 110 198 158 6102
rect 6062 198 6110 6102
rect 110 150 6110 198
rect 6429 6102 12429 6150
rect 6429 198 6477 6102
rect 12381 198 12429 6102
rect 6429 150 12429 198
rect -12528 -198 -6528 -150
rect -12528 -6102 -12480 -198
rect -6576 -6102 -6528 -198
rect -12528 -6150 -6528 -6102
rect -6209 -198 -209 -150
rect -6209 -6102 -6161 -198
rect -257 -6102 -209 -198
rect -6209 -6150 -209 -6102
rect 110 -198 6110 -150
rect 110 -6102 158 -198
rect 6062 -6102 6110 -198
rect 110 -6150 6110 -6102
rect 6429 -198 12429 -150
rect 6429 -6102 6477 -198
rect 12381 -6102 12429 -198
rect 6429 -6150 12429 -6102
rect -12528 -6498 -6528 -6450
rect -12528 -12402 -12480 -6498
rect -6576 -12402 -6528 -6498
rect -12528 -12450 -6528 -12402
rect -6209 -6498 -209 -6450
rect -6209 -12402 -6161 -6498
rect -257 -12402 -209 -6498
rect -6209 -12450 -209 -12402
rect 110 -6498 6110 -6450
rect 110 -12402 158 -6498
rect 6062 -12402 6110 -6498
rect 110 -12450 6110 -12402
rect 6429 -6498 12429 -6450
rect 6429 -12402 6477 -6498
rect 12381 -12402 12429 -6498
rect 6429 -12450 12429 -12402
<< mimcapcontact >>
rect -12480 6498 -6576 12402
rect -6161 6498 -257 12402
rect 158 6498 6062 12402
rect 6477 6498 12381 12402
rect -12480 198 -6576 6102
rect -6161 198 -257 6102
rect 158 198 6062 6102
rect 6477 198 12381 6102
rect -12480 -6102 -6576 -198
rect -6161 -6102 -257 -198
rect 158 -6102 6062 -198
rect 6477 -6102 12381 -198
rect -12480 -12402 -6576 -6498
rect -6161 -12402 -257 -6498
rect 158 -12402 6062 -6498
rect 6477 -12402 12381 -6498
<< metal4 >>
rect -9580 12411 -9476 12600
rect -6460 12538 -6356 12600
rect -6460 12522 -6333 12538
rect -6460 12458 -6413 12522
rect -6349 12458 -6333 12522
rect -6460 12442 -6333 12458
rect -12489 12402 -6567 12411
rect -12489 6498 -12480 12402
rect -6576 6498 -6567 12402
rect -12489 6489 -6567 6498
rect -6460 12378 -6413 12442
rect -6349 12378 -6333 12442
rect -3261 12411 -3157 12600
rect -141 12538 -37 12600
rect -141 12522 -14 12538
rect -141 12458 -94 12522
rect -30 12458 -14 12522
rect -141 12442 -14 12458
rect -6460 12362 -6333 12378
rect -6460 12298 -6413 12362
rect -6349 12298 -6333 12362
rect -6460 12282 -6333 12298
rect -6460 12218 -6413 12282
rect -6349 12218 -6333 12282
rect -6460 12202 -6333 12218
rect -6460 12138 -6413 12202
rect -6349 12138 -6333 12202
rect -6460 12122 -6333 12138
rect -6460 12058 -6413 12122
rect -6349 12058 -6333 12122
rect -6460 12042 -6333 12058
rect -6460 11978 -6413 12042
rect -6349 11978 -6333 12042
rect -6460 11962 -6333 11978
rect -6460 11898 -6413 11962
rect -6349 11898 -6333 11962
rect -6460 11882 -6333 11898
rect -6460 11818 -6413 11882
rect -6349 11818 -6333 11882
rect -6460 11802 -6333 11818
rect -6460 11738 -6413 11802
rect -6349 11738 -6333 11802
rect -6460 11722 -6333 11738
rect -6460 11658 -6413 11722
rect -6349 11658 -6333 11722
rect -6460 11642 -6333 11658
rect -6460 11578 -6413 11642
rect -6349 11578 -6333 11642
rect -6460 11562 -6333 11578
rect -6460 11498 -6413 11562
rect -6349 11498 -6333 11562
rect -6460 11482 -6333 11498
rect -6460 11418 -6413 11482
rect -6349 11418 -6333 11482
rect -6460 11402 -6333 11418
rect -6460 11338 -6413 11402
rect -6349 11338 -6333 11402
rect -6460 11322 -6333 11338
rect -6460 11258 -6413 11322
rect -6349 11258 -6333 11322
rect -6460 11242 -6333 11258
rect -6460 11178 -6413 11242
rect -6349 11178 -6333 11242
rect -6460 11162 -6333 11178
rect -6460 11098 -6413 11162
rect -6349 11098 -6333 11162
rect -6460 11082 -6333 11098
rect -6460 11018 -6413 11082
rect -6349 11018 -6333 11082
rect -6460 11002 -6333 11018
rect -6460 10938 -6413 11002
rect -6349 10938 -6333 11002
rect -6460 10922 -6333 10938
rect -6460 10858 -6413 10922
rect -6349 10858 -6333 10922
rect -6460 10842 -6333 10858
rect -6460 10778 -6413 10842
rect -6349 10778 -6333 10842
rect -6460 10762 -6333 10778
rect -6460 10698 -6413 10762
rect -6349 10698 -6333 10762
rect -6460 10682 -6333 10698
rect -6460 10618 -6413 10682
rect -6349 10618 -6333 10682
rect -6460 10602 -6333 10618
rect -6460 10538 -6413 10602
rect -6349 10538 -6333 10602
rect -6460 10522 -6333 10538
rect -6460 10458 -6413 10522
rect -6349 10458 -6333 10522
rect -6460 10442 -6333 10458
rect -6460 10378 -6413 10442
rect -6349 10378 -6333 10442
rect -6460 10362 -6333 10378
rect -6460 10298 -6413 10362
rect -6349 10298 -6333 10362
rect -6460 10282 -6333 10298
rect -6460 10218 -6413 10282
rect -6349 10218 -6333 10282
rect -6460 10202 -6333 10218
rect -6460 10138 -6413 10202
rect -6349 10138 -6333 10202
rect -6460 10122 -6333 10138
rect -6460 10058 -6413 10122
rect -6349 10058 -6333 10122
rect -6460 10042 -6333 10058
rect -6460 9978 -6413 10042
rect -6349 9978 -6333 10042
rect -6460 9962 -6333 9978
rect -6460 9898 -6413 9962
rect -6349 9898 -6333 9962
rect -6460 9882 -6333 9898
rect -6460 9818 -6413 9882
rect -6349 9818 -6333 9882
rect -6460 9802 -6333 9818
rect -6460 9738 -6413 9802
rect -6349 9738 -6333 9802
rect -6460 9722 -6333 9738
rect -6460 9658 -6413 9722
rect -6349 9658 -6333 9722
rect -6460 9642 -6333 9658
rect -6460 9578 -6413 9642
rect -6349 9578 -6333 9642
rect -6460 9562 -6333 9578
rect -6460 9498 -6413 9562
rect -6349 9498 -6333 9562
rect -6460 9482 -6333 9498
rect -6460 9418 -6413 9482
rect -6349 9418 -6333 9482
rect -6460 9402 -6333 9418
rect -6460 9338 -6413 9402
rect -6349 9338 -6333 9402
rect -6460 9322 -6333 9338
rect -6460 9258 -6413 9322
rect -6349 9258 -6333 9322
rect -6460 9242 -6333 9258
rect -6460 9178 -6413 9242
rect -6349 9178 -6333 9242
rect -6460 9162 -6333 9178
rect -6460 9098 -6413 9162
rect -6349 9098 -6333 9162
rect -6460 9082 -6333 9098
rect -6460 9018 -6413 9082
rect -6349 9018 -6333 9082
rect -6460 9002 -6333 9018
rect -6460 8938 -6413 9002
rect -6349 8938 -6333 9002
rect -6460 8922 -6333 8938
rect -6460 8858 -6413 8922
rect -6349 8858 -6333 8922
rect -6460 8842 -6333 8858
rect -6460 8778 -6413 8842
rect -6349 8778 -6333 8842
rect -6460 8762 -6333 8778
rect -6460 8698 -6413 8762
rect -6349 8698 -6333 8762
rect -6460 8682 -6333 8698
rect -6460 8618 -6413 8682
rect -6349 8618 -6333 8682
rect -6460 8602 -6333 8618
rect -6460 8538 -6413 8602
rect -6349 8538 -6333 8602
rect -6460 8522 -6333 8538
rect -6460 8458 -6413 8522
rect -6349 8458 -6333 8522
rect -6460 8442 -6333 8458
rect -6460 8378 -6413 8442
rect -6349 8378 -6333 8442
rect -6460 8362 -6333 8378
rect -6460 8298 -6413 8362
rect -6349 8298 -6333 8362
rect -6460 8282 -6333 8298
rect -6460 8218 -6413 8282
rect -6349 8218 -6333 8282
rect -6460 8202 -6333 8218
rect -6460 8138 -6413 8202
rect -6349 8138 -6333 8202
rect -6460 8122 -6333 8138
rect -6460 8058 -6413 8122
rect -6349 8058 -6333 8122
rect -6460 8042 -6333 8058
rect -6460 7978 -6413 8042
rect -6349 7978 -6333 8042
rect -6460 7962 -6333 7978
rect -6460 7898 -6413 7962
rect -6349 7898 -6333 7962
rect -6460 7882 -6333 7898
rect -6460 7818 -6413 7882
rect -6349 7818 -6333 7882
rect -6460 7802 -6333 7818
rect -6460 7738 -6413 7802
rect -6349 7738 -6333 7802
rect -6460 7722 -6333 7738
rect -6460 7658 -6413 7722
rect -6349 7658 -6333 7722
rect -6460 7642 -6333 7658
rect -6460 7578 -6413 7642
rect -6349 7578 -6333 7642
rect -6460 7562 -6333 7578
rect -6460 7498 -6413 7562
rect -6349 7498 -6333 7562
rect -6460 7482 -6333 7498
rect -6460 7418 -6413 7482
rect -6349 7418 -6333 7482
rect -6460 7402 -6333 7418
rect -6460 7338 -6413 7402
rect -6349 7338 -6333 7402
rect -6460 7322 -6333 7338
rect -6460 7258 -6413 7322
rect -6349 7258 -6333 7322
rect -6460 7242 -6333 7258
rect -6460 7178 -6413 7242
rect -6349 7178 -6333 7242
rect -6460 7162 -6333 7178
rect -6460 7098 -6413 7162
rect -6349 7098 -6333 7162
rect -6460 7082 -6333 7098
rect -6460 7018 -6413 7082
rect -6349 7018 -6333 7082
rect -6460 7002 -6333 7018
rect -6460 6938 -6413 7002
rect -6349 6938 -6333 7002
rect -6460 6922 -6333 6938
rect -6460 6858 -6413 6922
rect -6349 6858 -6333 6922
rect -6460 6842 -6333 6858
rect -6460 6778 -6413 6842
rect -6349 6778 -6333 6842
rect -6460 6762 -6333 6778
rect -6460 6698 -6413 6762
rect -6349 6698 -6333 6762
rect -6460 6682 -6333 6698
rect -6460 6618 -6413 6682
rect -6349 6618 -6333 6682
rect -6460 6602 -6333 6618
rect -6460 6538 -6413 6602
rect -6349 6538 -6333 6602
rect -6460 6522 -6333 6538
rect -9580 6111 -9476 6489
rect -6460 6458 -6413 6522
rect -6349 6458 -6333 6522
rect -6170 12402 -248 12411
rect -6170 6498 -6161 12402
rect -257 6498 -248 12402
rect -6170 6489 -248 6498
rect -141 12378 -94 12442
rect -30 12378 -14 12442
rect 3058 12411 3162 12600
rect 6178 12538 6282 12600
rect 6178 12522 6305 12538
rect 6178 12458 6225 12522
rect 6289 12458 6305 12522
rect 6178 12442 6305 12458
rect -141 12362 -14 12378
rect -141 12298 -94 12362
rect -30 12298 -14 12362
rect -141 12282 -14 12298
rect -141 12218 -94 12282
rect -30 12218 -14 12282
rect -141 12202 -14 12218
rect -141 12138 -94 12202
rect -30 12138 -14 12202
rect -141 12122 -14 12138
rect -141 12058 -94 12122
rect -30 12058 -14 12122
rect -141 12042 -14 12058
rect -141 11978 -94 12042
rect -30 11978 -14 12042
rect -141 11962 -14 11978
rect -141 11898 -94 11962
rect -30 11898 -14 11962
rect -141 11882 -14 11898
rect -141 11818 -94 11882
rect -30 11818 -14 11882
rect -141 11802 -14 11818
rect -141 11738 -94 11802
rect -30 11738 -14 11802
rect -141 11722 -14 11738
rect -141 11658 -94 11722
rect -30 11658 -14 11722
rect -141 11642 -14 11658
rect -141 11578 -94 11642
rect -30 11578 -14 11642
rect -141 11562 -14 11578
rect -141 11498 -94 11562
rect -30 11498 -14 11562
rect -141 11482 -14 11498
rect -141 11418 -94 11482
rect -30 11418 -14 11482
rect -141 11402 -14 11418
rect -141 11338 -94 11402
rect -30 11338 -14 11402
rect -141 11322 -14 11338
rect -141 11258 -94 11322
rect -30 11258 -14 11322
rect -141 11242 -14 11258
rect -141 11178 -94 11242
rect -30 11178 -14 11242
rect -141 11162 -14 11178
rect -141 11098 -94 11162
rect -30 11098 -14 11162
rect -141 11082 -14 11098
rect -141 11018 -94 11082
rect -30 11018 -14 11082
rect -141 11002 -14 11018
rect -141 10938 -94 11002
rect -30 10938 -14 11002
rect -141 10922 -14 10938
rect -141 10858 -94 10922
rect -30 10858 -14 10922
rect -141 10842 -14 10858
rect -141 10778 -94 10842
rect -30 10778 -14 10842
rect -141 10762 -14 10778
rect -141 10698 -94 10762
rect -30 10698 -14 10762
rect -141 10682 -14 10698
rect -141 10618 -94 10682
rect -30 10618 -14 10682
rect -141 10602 -14 10618
rect -141 10538 -94 10602
rect -30 10538 -14 10602
rect -141 10522 -14 10538
rect -141 10458 -94 10522
rect -30 10458 -14 10522
rect -141 10442 -14 10458
rect -141 10378 -94 10442
rect -30 10378 -14 10442
rect -141 10362 -14 10378
rect -141 10298 -94 10362
rect -30 10298 -14 10362
rect -141 10282 -14 10298
rect -141 10218 -94 10282
rect -30 10218 -14 10282
rect -141 10202 -14 10218
rect -141 10138 -94 10202
rect -30 10138 -14 10202
rect -141 10122 -14 10138
rect -141 10058 -94 10122
rect -30 10058 -14 10122
rect -141 10042 -14 10058
rect -141 9978 -94 10042
rect -30 9978 -14 10042
rect -141 9962 -14 9978
rect -141 9898 -94 9962
rect -30 9898 -14 9962
rect -141 9882 -14 9898
rect -141 9818 -94 9882
rect -30 9818 -14 9882
rect -141 9802 -14 9818
rect -141 9738 -94 9802
rect -30 9738 -14 9802
rect -141 9722 -14 9738
rect -141 9658 -94 9722
rect -30 9658 -14 9722
rect -141 9642 -14 9658
rect -141 9578 -94 9642
rect -30 9578 -14 9642
rect -141 9562 -14 9578
rect -141 9498 -94 9562
rect -30 9498 -14 9562
rect -141 9482 -14 9498
rect -141 9418 -94 9482
rect -30 9418 -14 9482
rect -141 9402 -14 9418
rect -141 9338 -94 9402
rect -30 9338 -14 9402
rect -141 9322 -14 9338
rect -141 9258 -94 9322
rect -30 9258 -14 9322
rect -141 9242 -14 9258
rect -141 9178 -94 9242
rect -30 9178 -14 9242
rect -141 9162 -14 9178
rect -141 9098 -94 9162
rect -30 9098 -14 9162
rect -141 9082 -14 9098
rect -141 9018 -94 9082
rect -30 9018 -14 9082
rect -141 9002 -14 9018
rect -141 8938 -94 9002
rect -30 8938 -14 9002
rect -141 8922 -14 8938
rect -141 8858 -94 8922
rect -30 8858 -14 8922
rect -141 8842 -14 8858
rect -141 8778 -94 8842
rect -30 8778 -14 8842
rect -141 8762 -14 8778
rect -141 8698 -94 8762
rect -30 8698 -14 8762
rect -141 8682 -14 8698
rect -141 8618 -94 8682
rect -30 8618 -14 8682
rect -141 8602 -14 8618
rect -141 8538 -94 8602
rect -30 8538 -14 8602
rect -141 8522 -14 8538
rect -141 8458 -94 8522
rect -30 8458 -14 8522
rect -141 8442 -14 8458
rect -141 8378 -94 8442
rect -30 8378 -14 8442
rect -141 8362 -14 8378
rect -141 8298 -94 8362
rect -30 8298 -14 8362
rect -141 8282 -14 8298
rect -141 8218 -94 8282
rect -30 8218 -14 8282
rect -141 8202 -14 8218
rect -141 8138 -94 8202
rect -30 8138 -14 8202
rect -141 8122 -14 8138
rect -141 8058 -94 8122
rect -30 8058 -14 8122
rect -141 8042 -14 8058
rect -141 7978 -94 8042
rect -30 7978 -14 8042
rect -141 7962 -14 7978
rect -141 7898 -94 7962
rect -30 7898 -14 7962
rect -141 7882 -14 7898
rect -141 7818 -94 7882
rect -30 7818 -14 7882
rect -141 7802 -14 7818
rect -141 7738 -94 7802
rect -30 7738 -14 7802
rect -141 7722 -14 7738
rect -141 7658 -94 7722
rect -30 7658 -14 7722
rect -141 7642 -14 7658
rect -141 7578 -94 7642
rect -30 7578 -14 7642
rect -141 7562 -14 7578
rect -141 7498 -94 7562
rect -30 7498 -14 7562
rect -141 7482 -14 7498
rect -141 7418 -94 7482
rect -30 7418 -14 7482
rect -141 7402 -14 7418
rect -141 7338 -94 7402
rect -30 7338 -14 7402
rect -141 7322 -14 7338
rect -141 7258 -94 7322
rect -30 7258 -14 7322
rect -141 7242 -14 7258
rect -141 7178 -94 7242
rect -30 7178 -14 7242
rect -141 7162 -14 7178
rect -141 7098 -94 7162
rect -30 7098 -14 7162
rect -141 7082 -14 7098
rect -141 7018 -94 7082
rect -30 7018 -14 7082
rect -141 7002 -14 7018
rect -141 6938 -94 7002
rect -30 6938 -14 7002
rect -141 6922 -14 6938
rect -141 6858 -94 6922
rect -30 6858 -14 6922
rect -141 6842 -14 6858
rect -141 6778 -94 6842
rect -30 6778 -14 6842
rect -141 6762 -14 6778
rect -141 6698 -94 6762
rect -30 6698 -14 6762
rect -141 6682 -14 6698
rect -141 6618 -94 6682
rect -30 6618 -14 6682
rect -141 6602 -14 6618
rect -141 6538 -94 6602
rect -30 6538 -14 6602
rect -141 6522 -14 6538
rect -6460 6442 -6333 6458
rect -6460 6378 -6413 6442
rect -6349 6378 -6333 6442
rect -6460 6362 -6333 6378
rect -6460 6238 -6356 6362
rect -6460 6222 -6333 6238
rect -6460 6158 -6413 6222
rect -6349 6158 -6333 6222
rect -6460 6142 -6333 6158
rect -12489 6102 -6567 6111
rect -12489 198 -12480 6102
rect -6576 198 -6567 6102
rect -12489 189 -6567 198
rect -6460 6078 -6413 6142
rect -6349 6078 -6333 6142
rect -3261 6111 -3157 6489
rect -141 6458 -94 6522
rect -30 6458 -14 6522
rect 149 12402 6071 12411
rect 149 6498 158 12402
rect 6062 6498 6071 12402
rect 149 6489 6071 6498
rect 6178 12378 6225 12442
rect 6289 12378 6305 12442
rect 9377 12411 9481 12600
rect 12497 12538 12601 12600
rect 12497 12522 12624 12538
rect 12497 12458 12544 12522
rect 12608 12458 12624 12522
rect 12497 12442 12624 12458
rect 6178 12362 6305 12378
rect 6178 12298 6225 12362
rect 6289 12298 6305 12362
rect 6178 12282 6305 12298
rect 6178 12218 6225 12282
rect 6289 12218 6305 12282
rect 6178 12202 6305 12218
rect 6178 12138 6225 12202
rect 6289 12138 6305 12202
rect 6178 12122 6305 12138
rect 6178 12058 6225 12122
rect 6289 12058 6305 12122
rect 6178 12042 6305 12058
rect 6178 11978 6225 12042
rect 6289 11978 6305 12042
rect 6178 11962 6305 11978
rect 6178 11898 6225 11962
rect 6289 11898 6305 11962
rect 6178 11882 6305 11898
rect 6178 11818 6225 11882
rect 6289 11818 6305 11882
rect 6178 11802 6305 11818
rect 6178 11738 6225 11802
rect 6289 11738 6305 11802
rect 6178 11722 6305 11738
rect 6178 11658 6225 11722
rect 6289 11658 6305 11722
rect 6178 11642 6305 11658
rect 6178 11578 6225 11642
rect 6289 11578 6305 11642
rect 6178 11562 6305 11578
rect 6178 11498 6225 11562
rect 6289 11498 6305 11562
rect 6178 11482 6305 11498
rect 6178 11418 6225 11482
rect 6289 11418 6305 11482
rect 6178 11402 6305 11418
rect 6178 11338 6225 11402
rect 6289 11338 6305 11402
rect 6178 11322 6305 11338
rect 6178 11258 6225 11322
rect 6289 11258 6305 11322
rect 6178 11242 6305 11258
rect 6178 11178 6225 11242
rect 6289 11178 6305 11242
rect 6178 11162 6305 11178
rect 6178 11098 6225 11162
rect 6289 11098 6305 11162
rect 6178 11082 6305 11098
rect 6178 11018 6225 11082
rect 6289 11018 6305 11082
rect 6178 11002 6305 11018
rect 6178 10938 6225 11002
rect 6289 10938 6305 11002
rect 6178 10922 6305 10938
rect 6178 10858 6225 10922
rect 6289 10858 6305 10922
rect 6178 10842 6305 10858
rect 6178 10778 6225 10842
rect 6289 10778 6305 10842
rect 6178 10762 6305 10778
rect 6178 10698 6225 10762
rect 6289 10698 6305 10762
rect 6178 10682 6305 10698
rect 6178 10618 6225 10682
rect 6289 10618 6305 10682
rect 6178 10602 6305 10618
rect 6178 10538 6225 10602
rect 6289 10538 6305 10602
rect 6178 10522 6305 10538
rect 6178 10458 6225 10522
rect 6289 10458 6305 10522
rect 6178 10442 6305 10458
rect 6178 10378 6225 10442
rect 6289 10378 6305 10442
rect 6178 10362 6305 10378
rect 6178 10298 6225 10362
rect 6289 10298 6305 10362
rect 6178 10282 6305 10298
rect 6178 10218 6225 10282
rect 6289 10218 6305 10282
rect 6178 10202 6305 10218
rect 6178 10138 6225 10202
rect 6289 10138 6305 10202
rect 6178 10122 6305 10138
rect 6178 10058 6225 10122
rect 6289 10058 6305 10122
rect 6178 10042 6305 10058
rect 6178 9978 6225 10042
rect 6289 9978 6305 10042
rect 6178 9962 6305 9978
rect 6178 9898 6225 9962
rect 6289 9898 6305 9962
rect 6178 9882 6305 9898
rect 6178 9818 6225 9882
rect 6289 9818 6305 9882
rect 6178 9802 6305 9818
rect 6178 9738 6225 9802
rect 6289 9738 6305 9802
rect 6178 9722 6305 9738
rect 6178 9658 6225 9722
rect 6289 9658 6305 9722
rect 6178 9642 6305 9658
rect 6178 9578 6225 9642
rect 6289 9578 6305 9642
rect 6178 9562 6305 9578
rect 6178 9498 6225 9562
rect 6289 9498 6305 9562
rect 6178 9482 6305 9498
rect 6178 9418 6225 9482
rect 6289 9418 6305 9482
rect 6178 9402 6305 9418
rect 6178 9338 6225 9402
rect 6289 9338 6305 9402
rect 6178 9322 6305 9338
rect 6178 9258 6225 9322
rect 6289 9258 6305 9322
rect 6178 9242 6305 9258
rect 6178 9178 6225 9242
rect 6289 9178 6305 9242
rect 6178 9162 6305 9178
rect 6178 9098 6225 9162
rect 6289 9098 6305 9162
rect 6178 9082 6305 9098
rect 6178 9018 6225 9082
rect 6289 9018 6305 9082
rect 6178 9002 6305 9018
rect 6178 8938 6225 9002
rect 6289 8938 6305 9002
rect 6178 8922 6305 8938
rect 6178 8858 6225 8922
rect 6289 8858 6305 8922
rect 6178 8842 6305 8858
rect 6178 8778 6225 8842
rect 6289 8778 6305 8842
rect 6178 8762 6305 8778
rect 6178 8698 6225 8762
rect 6289 8698 6305 8762
rect 6178 8682 6305 8698
rect 6178 8618 6225 8682
rect 6289 8618 6305 8682
rect 6178 8602 6305 8618
rect 6178 8538 6225 8602
rect 6289 8538 6305 8602
rect 6178 8522 6305 8538
rect 6178 8458 6225 8522
rect 6289 8458 6305 8522
rect 6178 8442 6305 8458
rect 6178 8378 6225 8442
rect 6289 8378 6305 8442
rect 6178 8362 6305 8378
rect 6178 8298 6225 8362
rect 6289 8298 6305 8362
rect 6178 8282 6305 8298
rect 6178 8218 6225 8282
rect 6289 8218 6305 8282
rect 6178 8202 6305 8218
rect 6178 8138 6225 8202
rect 6289 8138 6305 8202
rect 6178 8122 6305 8138
rect 6178 8058 6225 8122
rect 6289 8058 6305 8122
rect 6178 8042 6305 8058
rect 6178 7978 6225 8042
rect 6289 7978 6305 8042
rect 6178 7962 6305 7978
rect 6178 7898 6225 7962
rect 6289 7898 6305 7962
rect 6178 7882 6305 7898
rect 6178 7818 6225 7882
rect 6289 7818 6305 7882
rect 6178 7802 6305 7818
rect 6178 7738 6225 7802
rect 6289 7738 6305 7802
rect 6178 7722 6305 7738
rect 6178 7658 6225 7722
rect 6289 7658 6305 7722
rect 6178 7642 6305 7658
rect 6178 7578 6225 7642
rect 6289 7578 6305 7642
rect 6178 7562 6305 7578
rect 6178 7498 6225 7562
rect 6289 7498 6305 7562
rect 6178 7482 6305 7498
rect 6178 7418 6225 7482
rect 6289 7418 6305 7482
rect 6178 7402 6305 7418
rect 6178 7338 6225 7402
rect 6289 7338 6305 7402
rect 6178 7322 6305 7338
rect 6178 7258 6225 7322
rect 6289 7258 6305 7322
rect 6178 7242 6305 7258
rect 6178 7178 6225 7242
rect 6289 7178 6305 7242
rect 6178 7162 6305 7178
rect 6178 7098 6225 7162
rect 6289 7098 6305 7162
rect 6178 7082 6305 7098
rect 6178 7018 6225 7082
rect 6289 7018 6305 7082
rect 6178 7002 6305 7018
rect 6178 6938 6225 7002
rect 6289 6938 6305 7002
rect 6178 6922 6305 6938
rect 6178 6858 6225 6922
rect 6289 6858 6305 6922
rect 6178 6842 6305 6858
rect 6178 6778 6225 6842
rect 6289 6778 6305 6842
rect 6178 6762 6305 6778
rect 6178 6698 6225 6762
rect 6289 6698 6305 6762
rect 6178 6682 6305 6698
rect 6178 6618 6225 6682
rect 6289 6618 6305 6682
rect 6178 6602 6305 6618
rect 6178 6538 6225 6602
rect 6289 6538 6305 6602
rect 6178 6522 6305 6538
rect -141 6442 -14 6458
rect -141 6378 -94 6442
rect -30 6378 -14 6442
rect -141 6362 -14 6378
rect -141 6238 -37 6362
rect -141 6222 -14 6238
rect -141 6158 -94 6222
rect -30 6158 -14 6222
rect -141 6142 -14 6158
rect -6460 6062 -6333 6078
rect -6460 5998 -6413 6062
rect -6349 5998 -6333 6062
rect -6460 5982 -6333 5998
rect -6460 5918 -6413 5982
rect -6349 5918 -6333 5982
rect -6460 5902 -6333 5918
rect -6460 5838 -6413 5902
rect -6349 5838 -6333 5902
rect -6460 5822 -6333 5838
rect -6460 5758 -6413 5822
rect -6349 5758 -6333 5822
rect -6460 5742 -6333 5758
rect -6460 5678 -6413 5742
rect -6349 5678 -6333 5742
rect -6460 5662 -6333 5678
rect -6460 5598 -6413 5662
rect -6349 5598 -6333 5662
rect -6460 5582 -6333 5598
rect -6460 5518 -6413 5582
rect -6349 5518 -6333 5582
rect -6460 5502 -6333 5518
rect -6460 5438 -6413 5502
rect -6349 5438 -6333 5502
rect -6460 5422 -6333 5438
rect -6460 5358 -6413 5422
rect -6349 5358 -6333 5422
rect -6460 5342 -6333 5358
rect -6460 5278 -6413 5342
rect -6349 5278 -6333 5342
rect -6460 5262 -6333 5278
rect -6460 5198 -6413 5262
rect -6349 5198 -6333 5262
rect -6460 5182 -6333 5198
rect -6460 5118 -6413 5182
rect -6349 5118 -6333 5182
rect -6460 5102 -6333 5118
rect -6460 5038 -6413 5102
rect -6349 5038 -6333 5102
rect -6460 5022 -6333 5038
rect -6460 4958 -6413 5022
rect -6349 4958 -6333 5022
rect -6460 4942 -6333 4958
rect -6460 4878 -6413 4942
rect -6349 4878 -6333 4942
rect -6460 4862 -6333 4878
rect -6460 4798 -6413 4862
rect -6349 4798 -6333 4862
rect -6460 4782 -6333 4798
rect -6460 4718 -6413 4782
rect -6349 4718 -6333 4782
rect -6460 4702 -6333 4718
rect -6460 4638 -6413 4702
rect -6349 4638 -6333 4702
rect -6460 4622 -6333 4638
rect -6460 4558 -6413 4622
rect -6349 4558 -6333 4622
rect -6460 4542 -6333 4558
rect -6460 4478 -6413 4542
rect -6349 4478 -6333 4542
rect -6460 4462 -6333 4478
rect -6460 4398 -6413 4462
rect -6349 4398 -6333 4462
rect -6460 4382 -6333 4398
rect -6460 4318 -6413 4382
rect -6349 4318 -6333 4382
rect -6460 4302 -6333 4318
rect -6460 4238 -6413 4302
rect -6349 4238 -6333 4302
rect -6460 4222 -6333 4238
rect -6460 4158 -6413 4222
rect -6349 4158 -6333 4222
rect -6460 4142 -6333 4158
rect -6460 4078 -6413 4142
rect -6349 4078 -6333 4142
rect -6460 4062 -6333 4078
rect -6460 3998 -6413 4062
rect -6349 3998 -6333 4062
rect -6460 3982 -6333 3998
rect -6460 3918 -6413 3982
rect -6349 3918 -6333 3982
rect -6460 3902 -6333 3918
rect -6460 3838 -6413 3902
rect -6349 3838 -6333 3902
rect -6460 3822 -6333 3838
rect -6460 3758 -6413 3822
rect -6349 3758 -6333 3822
rect -6460 3742 -6333 3758
rect -6460 3678 -6413 3742
rect -6349 3678 -6333 3742
rect -6460 3662 -6333 3678
rect -6460 3598 -6413 3662
rect -6349 3598 -6333 3662
rect -6460 3582 -6333 3598
rect -6460 3518 -6413 3582
rect -6349 3518 -6333 3582
rect -6460 3502 -6333 3518
rect -6460 3438 -6413 3502
rect -6349 3438 -6333 3502
rect -6460 3422 -6333 3438
rect -6460 3358 -6413 3422
rect -6349 3358 -6333 3422
rect -6460 3342 -6333 3358
rect -6460 3278 -6413 3342
rect -6349 3278 -6333 3342
rect -6460 3262 -6333 3278
rect -6460 3198 -6413 3262
rect -6349 3198 -6333 3262
rect -6460 3182 -6333 3198
rect -6460 3118 -6413 3182
rect -6349 3118 -6333 3182
rect -6460 3102 -6333 3118
rect -6460 3038 -6413 3102
rect -6349 3038 -6333 3102
rect -6460 3022 -6333 3038
rect -6460 2958 -6413 3022
rect -6349 2958 -6333 3022
rect -6460 2942 -6333 2958
rect -6460 2878 -6413 2942
rect -6349 2878 -6333 2942
rect -6460 2862 -6333 2878
rect -6460 2798 -6413 2862
rect -6349 2798 -6333 2862
rect -6460 2782 -6333 2798
rect -6460 2718 -6413 2782
rect -6349 2718 -6333 2782
rect -6460 2702 -6333 2718
rect -6460 2638 -6413 2702
rect -6349 2638 -6333 2702
rect -6460 2622 -6333 2638
rect -6460 2558 -6413 2622
rect -6349 2558 -6333 2622
rect -6460 2542 -6333 2558
rect -6460 2478 -6413 2542
rect -6349 2478 -6333 2542
rect -6460 2462 -6333 2478
rect -6460 2398 -6413 2462
rect -6349 2398 -6333 2462
rect -6460 2382 -6333 2398
rect -6460 2318 -6413 2382
rect -6349 2318 -6333 2382
rect -6460 2302 -6333 2318
rect -6460 2238 -6413 2302
rect -6349 2238 -6333 2302
rect -6460 2222 -6333 2238
rect -6460 2158 -6413 2222
rect -6349 2158 -6333 2222
rect -6460 2142 -6333 2158
rect -6460 2078 -6413 2142
rect -6349 2078 -6333 2142
rect -6460 2062 -6333 2078
rect -6460 1998 -6413 2062
rect -6349 1998 -6333 2062
rect -6460 1982 -6333 1998
rect -6460 1918 -6413 1982
rect -6349 1918 -6333 1982
rect -6460 1902 -6333 1918
rect -6460 1838 -6413 1902
rect -6349 1838 -6333 1902
rect -6460 1822 -6333 1838
rect -6460 1758 -6413 1822
rect -6349 1758 -6333 1822
rect -6460 1742 -6333 1758
rect -6460 1678 -6413 1742
rect -6349 1678 -6333 1742
rect -6460 1662 -6333 1678
rect -6460 1598 -6413 1662
rect -6349 1598 -6333 1662
rect -6460 1582 -6333 1598
rect -6460 1518 -6413 1582
rect -6349 1518 -6333 1582
rect -6460 1502 -6333 1518
rect -6460 1438 -6413 1502
rect -6349 1438 -6333 1502
rect -6460 1422 -6333 1438
rect -6460 1358 -6413 1422
rect -6349 1358 -6333 1422
rect -6460 1342 -6333 1358
rect -6460 1278 -6413 1342
rect -6349 1278 -6333 1342
rect -6460 1262 -6333 1278
rect -6460 1198 -6413 1262
rect -6349 1198 -6333 1262
rect -6460 1182 -6333 1198
rect -6460 1118 -6413 1182
rect -6349 1118 -6333 1182
rect -6460 1102 -6333 1118
rect -6460 1038 -6413 1102
rect -6349 1038 -6333 1102
rect -6460 1022 -6333 1038
rect -6460 958 -6413 1022
rect -6349 958 -6333 1022
rect -6460 942 -6333 958
rect -6460 878 -6413 942
rect -6349 878 -6333 942
rect -6460 862 -6333 878
rect -6460 798 -6413 862
rect -6349 798 -6333 862
rect -6460 782 -6333 798
rect -6460 718 -6413 782
rect -6349 718 -6333 782
rect -6460 702 -6333 718
rect -6460 638 -6413 702
rect -6349 638 -6333 702
rect -6460 622 -6333 638
rect -6460 558 -6413 622
rect -6349 558 -6333 622
rect -6460 542 -6333 558
rect -6460 478 -6413 542
rect -6349 478 -6333 542
rect -6460 462 -6333 478
rect -6460 398 -6413 462
rect -6349 398 -6333 462
rect -6460 382 -6333 398
rect -6460 318 -6413 382
rect -6349 318 -6333 382
rect -6460 302 -6333 318
rect -6460 238 -6413 302
rect -6349 238 -6333 302
rect -6460 222 -6333 238
rect -9580 -189 -9476 189
rect -6460 158 -6413 222
rect -6349 158 -6333 222
rect -6170 6102 -248 6111
rect -6170 198 -6161 6102
rect -257 198 -248 6102
rect -6170 189 -248 198
rect -141 6078 -94 6142
rect -30 6078 -14 6142
rect 3058 6111 3162 6489
rect 6178 6458 6225 6522
rect 6289 6458 6305 6522
rect 6468 12402 12390 12411
rect 6468 6498 6477 12402
rect 12381 6498 12390 12402
rect 6468 6489 12390 6498
rect 12497 12378 12544 12442
rect 12608 12378 12624 12442
rect 12497 12362 12624 12378
rect 12497 12298 12544 12362
rect 12608 12298 12624 12362
rect 12497 12282 12624 12298
rect 12497 12218 12544 12282
rect 12608 12218 12624 12282
rect 12497 12202 12624 12218
rect 12497 12138 12544 12202
rect 12608 12138 12624 12202
rect 12497 12122 12624 12138
rect 12497 12058 12544 12122
rect 12608 12058 12624 12122
rect 12497 12042 12624 12058
rect 12497 11978 12544 12042
rect 12608 11978 12624 12042
rect 12497 11962 12624 11978
rect 12497 11898 12544 11962
rect 12608 11898 12624 11962
rect 12497 11882 12624 11898
rect 12497 11818 12544 11882
rect 12608 11818 12624 11882
rect 12497 11802 12624 11818
rect 12497 11738 12544 11802
rect 12608 11738 12624 11802
rect 12497 11722 12624 11738
rect 12497 11658 12544 11722
rect 12608 11658 12624 11722
rect 12497 11642 12624 11658
rect 12497 11578 12544 11642
rect 12608 11578 12624 11642
rect 12497 11562 12624 11578
rect 12497 11498 12544 11562
rect 12608 11498 12624 11562
rect 12497 11482 12624 11498
rect 12497 11418 12544 11482
rect 12608 11418 12624 11482
rect 12497 11402 12624 11418
rect 12497 11338 12544 11402
rect 12608 11338 12624 11402
rect 12497 11322 12624 11338
rect 12497 11258 12544 11322
rect 12608 11258 12624 11322
rect 12497 11242 12624 11258
rect 12497 11178 12544 11242
rect 12608 11178 12624 11242
rect 12497 11162 12624 11178
rect 12497 11098 12544 11162
rect 12608 11098 12624 11162
rect 12497 11082 12624 11098
rect 12497 11018 12544 11082
rect 12608 11018 12624 11082
rect 12497 11002 12624 11018
rect 12497 10938 12544 11002
rect 12608 10938 12624 11002
rect 12497 10922 12624 10938
rect 12497 10858 12544 10922
rect 12608 10858 12624 10922
rect 12497 10842 12624 10858
rect 12497 10778 12544 10842
rect 12608 10778 12624 10842
rect 12497 10762 12624 10778
rect 12497 10698 12544 10762
rect 12608 10698 12624 10762
rect 12497 10682 12624 10698
rect 12497 10618 12544 10682
rect 12608 10618 12624 10682
rect 12497 10602 12624 10618
rect 12497 10538 12544 10602
rect 12608 10538 12624 10602
rect 12497 10522 12624 10538
rect 12497 10458 12544 10522
rect 12608 10458 12624 10522
rect 12497 10442 12624 10458
rect 12497 10378 12544 10442
rect 12608 10378 12624 10442
rect 12497 10362 12624 10378
rect 12497 10298 12544 10362
rect 12608 10298 12624 10362
rect 12497 10282 12624 10298
rect 12497 10218 12544 10282
rect 12608 10218 12624 10282
rect 12497 10202 12624 10218
rect 12497 10138 12544 10202
rect 12608 10138 12624 10202
rect 12497 10122 12624 10138
rect 12497 10058 12544 10122
rect 12608 10058 12624 10122
rect 12497 10042 12624 10058
rect 12497 9978 12544 10042
rect 12608 9978 12624 10042
rect 12497 9962 12624 9978
rect 12497 9898 12544 9962
rect 12608 9898 12624 9962
rect 12497 9882 12624 9898
rect 12497 9818 12544 9882
rect 12608 9818 12624 9882
rect 12497 9802 12624 9818
rect 12497 9738 12544 9802
rect 12608 9738 12624 9802
rect 12497 9722 12624 9738
rect 12497 9658 12544 9722
rect 12608 9658 12624 9722
rect 12497 9642 12624 9658
rect 12497 9578 12544 9642
rect 12608 9578 12624 9642
rect 12497 9562 12624 9578
rect 12497 9498 12544 9562
rect 12608 9498 12624 9562
rect 12497 9482 12624 9498
rect 12497 9418 12544 9482
rect 12608 9418 12624 9482
rect 12497 9402 12624 9418
rect 12497 9338 12544 9402
rect 12608 9338 12624 9402
rect 12497 9322 12624 9338
rect 12497 9258 12544 9322
rect 12608 9258 12624 9322
rect 12497 9242 12624 9258
rect 12497 9178 12544 9242
rect 12608 9178 12624 9242
rect 12497 9162 12624 9178
rect 12497 9098 12544 9162
rect 12608 9098 12624 9162
rect 12497 9082 12624 9098
rect 12497 9018 12544 9082
rect 12608 9018 12624 9082
rect 12497 9002 12624 9018
rect 12497 8938 12544 9002
rect 12608 8938 12624 9002
rect 12497 8922 12624 8938
rect 12497 8858 12544 8922
rect 12608 8858 12624 8922
rect 12497 8842 12624 8858
rect 12497 8778 12544 8842
rect 12608 8778 12624 8842
rect 12497 8762 12624 8778
rect 12497 8698 12544 8762
rect 12608 8698 12624 8762
rect 12497 8682 12624 8698
rect 12497 8618 12544 8682
rect 12608 8618 12624 8682
rect 12497 8602 12624 8618
rect 12497 8538 12544 8602
rect 12608 8538 12624 8602
rect 12497 8522 12624 8538
rect 12497 8458 12544 8522
rect 12608 8458 12624 8522
rect 12497 8442 12624 8458
rect 12497 8378 12544 8442
rect 12608 8378 12624 8442
rect 12497 8362 12624 8378
rect 12497 8298 12544 8362
rect 12608 8298 12624 8362
rect 12497 8282 12624 8298
rect 12497 8218 12544 8282
rect 12608 8218 12624 8282
rect 12497 8202 12624 8218
rect 12497 8138 12544 8202
rect 12608 8138 12624 8202
rect 12497 8122 12624 8138
rect 12497 8058 12544 8122
rect 12608 8058 12624 8122
rect 12497 8042 12624 8058
rect 12497 7978 12544 8042
rect 12608 7978 12624 8042
rect 12497 7962 12624 7978
rect 12497 7898 12544 7962
rect 12608 7898 12624 7962
rect 12497 7882 12624 7898
rect 12497 7818 12544 7882
rect 12608 7818 12624 7882
rect 12497 7802 12624 7818
rect 12497 7738 12544 7802
rect 12608 7738 12624 7802
rect 12497 7722 12624 7738
rect 12497 7658 12544 7722
rect 12608 7658 12624 7722
rect 12497 7642 12624 7658
rect 12497 7578 12544 7642
rect 12608 7578 12624 7642
rect 12497 7562 12624 7578
rect 12497 7498 12544 7562
rect 12608 7498 12624 7562
rect 12497 7482 12624 7498
rect 12497 7418 12544 7482
rect 12608 7418 12624 7482
rect 12497 7402 12624 7418
rect 12497 7338 12544 7402
rect 12608 7338 12624 7402
rect 12497 7322 12624 7338
rect 12497 7258 12544 7322
rect 12608 7258 12624 7322
rect 12497 7242 12624 7258
rect 12497 7178 12544 7242
rect 12608 7178 12624 7242
rect 12497 7162 12624 7178
rect 12497 7098 12544 7162
rect 12608 7098 12624 7162
rect 12497 7082 12624 7098
rect 12497 7018 12544 7082
rect 12608 7018 12624 7082
rect 12497 7002 12624 7018
rect 12497 6938 12544 7002
rect 12608 6938 12624 7002
rect 12497 6922 12624 6938
rect 12497 6858 12544 6922
rect 12608 6858 12624 6922
rect 12497 6842 12624 6858
rect 12497 6778 12544 6842
rect 12608 6778 12624 6842
rect 12497 6762 12624 6778
rect 12497 6698 12544 6762
rect 12608 6698 12624 6762
rect 12497 6682 12624 6698
rect 12497 6618 12544 6682
rect 12608 6618 12624 6682
rect 12497 6602 12624 6618
rect 12497 6538 12544 6602
rect 12608 6538 12624 6602
rect 12497 6522 12624 6538
rect 6178 6442 6305 6458
rect 6178 6378 6225 6442
rect 6289 6378 6305 6442
rect 6178 6362 6305 6378
rect 6178 6238 6282 6362
rect 6178 6222 6305 6238
rect 6178 6158 6225 6222
rect 6289 6158 6305 6222
rect 6178 6142 6305 6158
rect -141 6062 -14 6078
rect -141 5998 -94 6062
rect -30 5998 -14 6062
rect -141 5982 -14 5998
rect -141 5918 -94 5982
rect -30 5918 -14 5982
rect -141 5902 -14 5918
rect -141 5838 -94 5902
rect -30 5838 -14 5902
rect -141 5822 -14 5838
rect -141 5758 -94 5822
rect -30 5758 -14 5822
rect -141 5742 -14 5758
rect -141 5678 -94 5742
rect -30 5678 -14 5742
rect -141 5662 -14 5678
rect -141 5598 -94 5662
rect -30 5598 -14 5662
rect -141 5582 -14 5598
rect -141 5518 -94 5582
rect -30 5518 -14 5582
rect -141 5502 -14 5518
rect -141 5438 -94 5502
rect -30 5438 -14 5502
rect -141 5422 -14 5438
rect -141 5358 -94 5422
rect -30 5358 -14 5422
rect -141 5342 -14 5358
rect -141 5278 -94 5342
rect -30 5278 -14 5342
rect -141 5262 -14 5278
rect -141 5198 -94 5262
rect -30 5198 -14 5262
rect -141 5182 -14 5198
rect -141 5118 -94 5182
rect -30 5118 -14 5182
rect -141 5102 -14 5118
rect -141 5038 -94 5102
rect -30 5038 -14 5102
rect -141 5022 -14 5038
rect -141 4958 -94 5022
rect -30 4958 -14 5022
rect -141 4942 -14 4958
rect -141 4878 -94 4942
rect -30 4878 -14 4942
rect -141 4862 -14 4878
rect -141 4798 -94 4862
rect -30 4798 -14 4862
rect -141 4782 -14 4798
rect -141 4718 -94 4782
rect -30 4718 -14 4782
rect -141 4702 -14 4718
rect -141 4638 -94 4702
rect -30 4638 -14 4702
rect -141 4622 -14 4638
rect -141 4558 -94 4622
rect -30 4558 -14 4622
rect -141 4542 -14 4558
rect -141 4478 -94 4542
rect -30 4478 -14 4542
rect -141 4462 -14 4478
rect -141 4398 -94 4462
rect -30 4398 -14 4462
rect -141 4382 -14 4398
rect -141 4318 -94 4382
rect -30 4318 -14 4382
rect -141 4302 -14 4318
rect -141 4238 -94 4302
rect -30 4238 -14 4302
rect -141 4222 -14 4238
rect -141 4158 -94 4222
rect -30 4158 -14 4222
rect -141 4142 -14 4158
rect -141 4078 -94 4142
rect -30 4078 -14 4142
rect -141 4062 -14 4078
rect -141 3998 -94 4062
rect -30 3998 -14 4062
rect -141 3982 -14 3998
rect -141 3918 -94 3982
rect -30 3918 -14 3982
rect -141 3902 -14 3918
rect -141 3838 -94 3902
rect -30 3838 -14 3902
rect -141 3822 -14 3838
rect -141 3758 -94 3822
rect -30 3758 -14 3822
rect -141 3742 -14 3758
rect -141 3678 -94 3742
rect -30 3678 -14 3742
rect -141 3662 -14 3678
rect -141 3598 -94 3662
rect -30 3598 -14 3662
rect -141 3582 -14 3598
rect -141 3518 -94 3582
rect -30 3518 -14 3582
rect -141 3502 -14 3518
rect -141 3438 -94 3502
rect -30 3438 -14 3502
rect -141 3422 -14 3438
rect -141 3358 -94 3422
rect -30 3358 -14 3422
rect -141 3342 -14 3358
rect -141 3278 -94 3342
rect -30 3278 -14 3342
rect -141 3262 -14 3278
rect -141 3198 -94 3262
rect -30 3198 -14 3262
rect -141 3182 -14 3198
rect -141 3118 -94 3182
rect -30 3118 -14 3182
rect -141 3102 -14 3118
rect -141 3038 -94 3102
rect -30 3038 -14 3102
rect -141 3022 -14 3038
rect -141 2958 -94 3022
rect -30 2958 -14 3022
rect -141 2942 -14 2958
rect -141 2878 -94 2942
rect -30 2878 -14 2942
rect -141 2862 -14 2878
rect -141 2798 -94 2862
rect -30 2798 -14 2862
rect -141 2782 -14 2798
rect -141 2718 -94 2782
rect -30 2718 -14 2782
rect -141 2702 -14 2718
rect -141 2638 -94 2702
rect -30 2638 -14 2702
rect -141 2622 -14 2638
rect -141 2558 -94 2622
rect -30 2558 -14 2622
rect -141 2542 -14 2558
rect -141 2478 -94 2542
rect -30 2478 -14 2542
rect -141 2462 -14 2478
rect -141 2398 -94 2462
rect -30 2398 -14 2462
rect -141 2382 -14 2398
rect -141 2318 -94 2382
rect -30 2318 -14 2382
rect -141 2302 -14 2318
rect -141 2238 -94 2302
rect -30 2238 -14 2302
rect -141 2222 -14 2238
rect -141 2158 -94 2222
rect -30 2158 -14 2222
rect -141 2142 -14 2158
rect -141 2078 -94 2142
rect -30 2078 -14 2142
rect -141 2062 -14 2078
rect -141 1998 -94 2062
rect -30 1998 -14 2062
rect -141 1982 -14 1998
rect -141 1918 -94 1982
rect -30 1918 -14 1982
rect -141 1902 -14 1918
rect -141 1838 -94 1902
rect -30 1838 -14 1902
rect -141 1822 -14 1838
rect -141 1758 -94 1822
rect -30 1758 -14 1822
rect -141 1742 -14 1758
rect -141 1678 -94 1742
rect -30 1678 -14 1742
rect -141 1662 -14 1678
rect -141 1598 -94 1662
rect -30 1598 -14 1662
rect -141 1582 -14 1598
rect -141 1518 -94 1582
rect -30 1518 -14 1582
rect -141 1502 -14 1518
rect -141 1438 -94 1502
rect -30 1438 -14 1502
rect -141 1422 -14 1438
rect -141 1358 -94 1422
rect -30 1358 -14 1422
rect -141 1342 -14 1358
rect -141 1278 -94 1342
rect -30 1278 -14 1342
rect -141 1262 -14 1278
rect -141 1198 -94 1262
rect -30 1198 -14 1262
rect -141 1182 -14 1198
rect -141 1118 -94 1182
rect -30 1118 -14 1182
rect -141 1102 -14 1118
rect -141 1038 -94 1102
rect -30 1038 -14 1102
rect -141 1022 -14 1038
rect -141 958 -94 1022
rect -30 958 -14 1022
rect -141 942 -14 958
rect -141 878 -94 942
rect -30 878 -14 942
rect -141 862 -14 878
rect -141 798 -94 862
rect -30 798 -14 862
rect -141 782 -14 798
rect -141 718 -94 782
rect -30 718 -14 782
rect -141 702 -14 718
rect -141 638 -94 702
rect -30 638 -14 702
rect -141 622 -14 638
rect -141 558 -94 622
rect -30 558 -14 622
rect -141 542 -14 558
rect -141 478 -94 542
rect -30 478 -14 542
rect -141 462 -14 478
rect -141 398 -94 462
rect -30 398 -14 462
rect -141 382 -14 398
rect -141 318 -94 382
rect -30 318 -14 382
rect -141 302 -14 318
rect -141 238 -94 302
rect -30 238 -14 302
rect -141 222 -14 238
rect -6460 142 -6333 158
rect -6460 78 -6413 142
rect -6349 78 -6333 142
rect -6460 62 -6333 78
rect -6460 -62 -6356 62
rect -6460 -78 -6333 -62
rect -6460 -142 -6413 -78
rect -6349 -142 -6333 -78
rect -6460 -158 -6333 -142
rect -12489 -198 -6567 -189
rect -12489 -6102 -12480 -198
rect -6576 -6102 -6567 -198
rect -12489 -6111 -6567 -6102
rect -6460 -222 -6413 -158
rect -6349 -222 -6333 -158
rect -3261 -189 -3157 189
rect -141 158 -94 222
rect -30 158 -14 222
rect 149 6102 6071 6111
rect 149 198 158 6102
rect 6062 198 6071 6102
rect 149 189 6071 198
rect 6178 6078 6225 6142
rect 6289 6078 6305 6142
rect 9377 6111 9481 6489
rect 12497 6458 12544 6522
rect 12608 6458 12624 6522
rect 12497 6442 12624 6458
rect 12497 6378 12544 6442
rect 12608 6378 12624 6442
rect 12497 6362 12624 6378
rect 12497 6238 12601 6362
rect 12497 6222 12624 6238
rect 12497 6158 12544 6222
rect 12608 6158 12624 6222
rect 12497 6142 12624 6158
rect 6178 6062 6305 6078
rect 6178 5998 6225 6062
rect 6289 5998 6305 6062
rect 6178 5982 6305 5998
rect 6178 5918 6225 5982
rect 6289 5918 6305 5982
rect 6178 5902 6305 5918
rect 6178 5838 6225 5902
rect 6289 5838 6305 5902
rect 6178 5822 6305 5838
rect 6178 5758 6225 5822
rect 6289 5758 6305 5822
rect 6178 5742 6305 5758
rect 6178 5678 6225 5742
rect 6289 5678 6305 5742
rect 6178 5662 6305 5678
rect 6178 5598 6225 5662
rect 6289 5598 6305 5662
rect 6178 5582 6305 5598
rect 6178 5518 6225 5582
rect 6289 5518 6305 5582
rect 6178 5502 6305 5518
rect 6178 5438 6225 5502
rect 6289 5438 6305 5502
rect 6178 5422 6305 5438
rect 6178 5358 6225 5422
rect 6289 5358 6305 5422
rect 6178 5342 6305 5358
rect 6178 5278 6225 5342
rect 6289 5278 6305 5342
rect 6178 5262 6305 5278
rect 6178 5198 6225 5262
rect 6289 5198 6305 5262
rect 6178 5182 6305 5198
rect 6178 5118 6225 5182
rect 6289 5118 6305 5182
rect 6178 5102 6305 5118
rect 6178 5038 6225 5102
rect 6289 5038 6305 5102
rect 6178 5022 6305 5038
rect 6178 4958 6225 5022
rect 6289 4958 6305 5022
rect 6178 4942 6305 4958
rect 6178 4878 6225 4942
rect 6289 4878 6305 4942
rect 6178 4862 6305 4878
rect 6178 4798 6225 4862
rect 6289 4798 6305 4862
rect 6178 4782 6305 4798
rect 6178 4718 6225 4782
rect 6289 4718 6305 4782
rect 6178 4702 6305 4718
rect 6178 4638 6225 4702
rect 6289 4638 6305 4702
rect 6178 4622 6305 4638
rect 6178 4558 6225 4622
rect 6289 4558 6305 4622
rect 6178 4542 6305 4558
rect 6178 4478 6225 4542
rect 6289 4478 6305 4542
rect 6178 4462 6305 4478
rect 6178 4398 6225 4462
rect 6289 4398 6305 4462
rect 6178 4382 6305 4398
rect 6178 4318 6225 4382
rect 6289 4318 6305 4382
rect 6178 4302 6305 4318
rect 6178 4238 6225 4302
rect 6289 4238 6305 4302
rect 6178 4222 6305 4238
rect 6178 4158 6225 4222
rect 6289 4158 6305 4222
rect 6178 4142 6305 4158
rect 6178 4078 6225 4142
rect 6289 4078 6305 4142
rect 6178 4062 6305 4078
rect 6178 3998 6225 4062
rect 6289 3998 6305 4062
rect 6178 3982 6305 3998
rect 6178 3918 6225 3982
rect 6289 3918 6305 3982
rect 6178 3902 6305 3918
rect 6178 3838 6225 3902
rect 6289 3838 6305 3902
rect 6178 3822 6305 3838
rect 6178 3758 6225 3822
rect 6289 3758 6305 3822
rect 6178 3742 6305 3758
rect 6178 3678 6225 3742
rect 6289 3678 6305 3742
rect 6178 3662 6305 3678
rect 6178 3598 6225 3662
rect 6289 3598 6305 3662
rect 6178 3582 6305 3598
rect 6178 3518 6225 3582
rect 6289 3518 6305 3582
rect 6178 3502 6305 3518
rect 6178 3438 6225 3502
rect 6289 3438 6305 3502
rect 6178 3422 6305 3438
rect 6178 3358 6225 3422
rect 6289 3358 6305 3422
rect 6178 3342 6305 3358
rect 6178 3278 6225 3342
rect 6289 3278 6305 3342
rect 6178 3262 6305 3278
rect 6178 3198 6225 3262
rect 6289 3198 6305 3262
rect 6178 3182 6305 3198
rect 6178 3118 6225 3182
rect 6289 3118 6305 3182
rect 6178 3102 6305 3118
rect 6178 3038 6225 3102
rect 6289 3038 6305 3102
rect 6178 3022 6305 3038
rect 6178 2958 6225 3022
rect 6289 2958 6305 3022
rect 6178 2942 6305 2958
rect 6178 2878 6225 2942
rect 6289 2878 6305 2942
rect 6178 2862 6305 2878
rect 6178 2798 6225 2862
rect 6289 2798 6305 2862
rect 6178 2782 6305 2798
rect 6178 2718 6225 2782
rect 6289 2718 6305 2782
rect 6178 2702 6305 2718
rect 6178 2638 6225 2702
rect 6289 2638 6305 2702
rect 6178 2622 6305 2638
rect 6178 2558 6225 2622
rect 6289 2558 6305 2622
rect 6178 2542 6305 2558
rect 6178 2478 6225 2542
rect 6289 2478 6305 2542
rect 6178 2462 6305 2478
rect 6178 2398 6225 2462
rect 6289 2398 6305 2462
rect 6178 2382 6305 2398
rect 6178 2318 6225 2382
rect 6289 2318 6305 2382
rect 6178 2302 6305 2318
rect 6178 2238 6225 2302
rect 6289 2238 6305 2302
rect 6178 2222 6305 2238
rect 6178 2158 6225 2222
rect 6289 2158 6305 2222
rect 6178 2142 6305 2158
rect 6178 2078 6225 2142
rect 6289 2078 6305 2142
rect 6178 2062 6305 2078
rect 6178 1998 6225 2062
rect 6289 1998 6305 2062
rect 6178 1982 6305 1998
rect 6178 1918 6225 1982
rect 6289 1918 6305 1982
rect 6178 1902 6305 1918
rect 6178 1838 6225 1902
rect 6289 1838 6305 1902
rect 6178 1822 6305 1838
rect 6178 1758 6225 1822
rect 6289 1758 6305 1822
rect 6178 1742 6305 1758
rect 6178 1678 6225 1742
rect 6289 1678 6305 1742
rect 6178 1662 6305 1678
rect 6178 1598 6225 1662
rect 6289 1598 6305 1662
rect 6178 1582 6305 1598
rect 6178 1518 6225 1582
rect 6289 1518 6305 1582
rect 6178 1502 6305 1518
rect 6178 1438 6225 1502
rect 6289 1438 6305 1502
rect 6178 1422 6305 1438
rect 6178 1358 6225 1422
rect 6289 1358 6305 1422
rect 6178 1342 6305 1358
rect 6178 1278 6225 1342
rect 6289 1278 6305 1342
rect 6178 1262 6305 1278
rect 6178 1198 6225 1262
rect 6289 1198 6305 1262
rect 6178 1182 6305 1198
rect 6178 1118 6225 1182
rect 6289 1118 6305 1182
rect 6178 1102 6305 1118
rect 6178 1038 6225 1102
rect 6289 1038 6305 1102
rect 6178 1022 6305 1038
rect 6178 958 6225 1022
rect 6289 958 6305 1022
rect 6178 942 6305 958
rect 6178 878 6225 942
rect 6289 878 6305 942
rect 6178 862 6305 878
rect 6178 798 6225 862
rect 6289 798 6305 862
rect 6178 782 6305 798
rect 6178 718 6225 782
rect 6289 718 6305 782
rect 6178 702 6305 718
rect 6178 638 6225 702
rect 6289 638 6305 702
rect 6178 622 6305 638
rect 6178 558 6225 622
rect 6289 558 6305 622
rect 6178 542 6305 558
rect 6178 478 6225 542
rect 6289 478 6305 542
rect 6178 462 6305 478
rect 6178 398 6225 462
rect 6289 398 6305 462
rect 6178 382 6305 398
rect 6178 318 6225 382
rect 6289 318 6305 382
rect 6178 302 6305 318
rect 6178 238 6225 302
rect 6289 238 6305 302
rect 6178 222 6305 238
rect -141 142 -14 158
rect -141 78 -94 142
rect -30 78 -14 142
rect -141 62 -14 78
rect -141 -62 -37 62
rect -141 -78 -14 -62
rect -141 -142 -94 -78
rect -30 -142 -14 -78
rect -141 -158 -14 -142
rect -6460 -238 -6333 -222
rect -6460 -302 -6413 -238
rect -6349 -302 -6333 -238
rect -6460 -318 -6333 -302
rect -6460 -382 -6413 -318
rect -6349 -382 -6333 -318
rect -6460 -398 -6333 -382
rect -6460 -462 -6413 -398
rect -6349 -462 -6333 -398
rect -6460 -478 -6333 -462
rect -6460 -542 -6413 -478
rect -6349 -542 -6333 -478
rect -6460 -558 -6333 -542
rect -6460 -622 -6413 -558
rect -6349 -622 -6333 -558
rect -6460 -638 -6333 -622
rect -6460 -702 -6413 -638
rect -6349 -702 -6333 -638
rect -6460 -718 -6333 -702
rect -6460 -782 -6413 -718
rect -6349 -782 -6333 -718
rect -6460 -798 -6333 -782
rect -6460 -862 -6413 -798
rect -6349 -862 -6333 -798
rect -6460 -878 -6333 -862
rect -6460 -942 -6413 -878
rect -6349 -942 -6333 -878
rect -6460 -958 -6333 -942
rect -6460 -1022 -6413 -958
rect -6349 -1022 -6333 -958
rect -6460 -1038 -6333 -1022
rect -6460 -1102 -6413 -1038
rect -6349 -1102 -6333 -1038
rect -6460 -1118 -6333 -1102
rect -6460 -1182 -6413 -1118
rect -6349 -1182 -6333 -1118
rect -6460 -1198 -6333 -1182
rect -6460 -1262 -6413 -1198
rect -6349 -1262 -6333 -1198
rect -6460 -1278 -6333 -1262
rect -6460 -1342 -6413 -1278
rect -6349 -1342 -6333 -1278
rect -6460 -1358 -6333 -1342
rect -6460 -1422 -6413 -1358
rect -6349 -1422 -6333 -1358
rect -6460 -1438 -6333 -1422
rect -6460 -1502 -6413 -1438
rect -6349 -1502 -6333 -1438
rect -6460 -1518 -6333 -1502
rect -6460 -1582 -6413 -1518
rect -6349 -1582 -6333 -1518
rect -6460 -1598 -6333 -1582
rect -6460 -1662 -6413 -1598
rect -6349 -1662 -6333 -1598
rect -6460 -1678 -6333 -1662
rect -6460 -1742 -6413 -1678
rect -6349 -1742 -6333 -1678
rect -6460 -1758 -6333 -1742
rect -6460 -1822 -6413 -1758
rect -6349 -1822 -6333 -1758
rect -6460 -1838 -6333 -1822
rect -6460 -1902 -6413 -1838
rect -6349 -1902 -6333 -1838
rect -6460 -1918 -6333 -1902
rect -6460 -1982 -6413 -1918
rect -6349 -1982 -6333 -1918
rect -6460 -1998 -6333 -1982
rect -6460 -2062 -6413 -1998
rect -6349 -2062 -6333 -1998
rect -6460 -2078 -6333 -2062
rect -6460 -2142 -6413 -2078
rect -6349 -2142 -6333 -2078
rect -6460 -2158 -6333 -2142
rect -6460 -2222 -6413 -2158
rect -6349 -2222 -6333 -2158
rect -6460 -2238 -6333 -2222
rect -6460 -2302 -6413 -2238
rect -6349 -2302 -6333 -2238
rect -6460 -2318 -6333 -2302
rect -6460 -2382 -6413 -2318
rect -6349 -2382 -6333 -2318
rect -6460 -2398 -6333 -2382
rect -6460 -2462 -6413 -2398
rect -6349 -2462 -6333 -2398
rect -6460 -2478 -6333 -2462
rect -6460 -2542 -6413 -2478
rect -6349 -2542 -6333 -2478
rect -6460 -2558 -6333 -2542
rect -6460 -2622 -6413 -2558
rect -6349 -2622 -6333 -2558
rect -6460 -2638 -6333 -2622
rect -6460 -2702 -6413 -2638
rect -6349 -2702 -6333 -2638
rect -6460 -2718 -6333 -2702
rect -6460 -2782 -6413 -2718
rect -6349 -2782 -6333 -2718
rect -6460 -2798 -6333 -2782
rect -6460 -2862 -6413 -2798
rect -6349 -2862 -6333 -2798
rect -6460 -2878 -6333 -2862
rect -6460 -2942 -6413 -2878
rect -6349 -2942 -6333 -2878
rect -6460 -2958 -6333 -2942
rect -6460 -3022 -6413 -2958
rect -6349 -3022 -6333 -2958
rect -6460 -3038 -6333 -3022
rect -6460 -3102 -6413 -3038
rect -6349 -3102 -6333 -3038
rect -6460 -3118 -6333 -3102
rect -6460 -3182 -6413 -3118
rect -6349 -3182 -6333 -3118
rect -6460 -3198 -6333 -3182
rect -6460 -3262 -6413 -3198
rect -6349 -3262 -6333 -3198
rect -6460 -3278 -6333 -3262
rect -6460 -3342 -6413 -3278
rect -6349 -3342 -6333 -3278
rect -6460 -3358 -6333 -3342
rect -6460 -3422 -6413 -3358
rect -6349 -3422 -6333 -3358
rect -6460 -3438 -6333 -3422
rect -6460 -3502 -6413 -3438
rect -6349 -3502 -6333 -3438
rect -6460 -3518 -6333 -3502
rect -6460 -3582 -6413 -3518
rect -6349 -3582 -6333 -3518
rect -6460 -3598 -6333 -3582
rect -6460 -3662 -6413 -3598
rect -6349 -3662 -6333 -3598
rect -6460 -3678 -6333 -3662
rect -6460 -3742 -6413 -3678
rect -6349 -3742 -6333 -3678
rect -6460 -3758 -6333 -3742
rect -6460 -3822 -6413 -3758
rect -6349 -3822 -6333 -3758
rect -6460 -3838 -6333 -3822
rect -6460 -3902 -6413 -3838
rect -6349 -3902 -6333 -3838
rect -6460 -3918 -6333 -3902
rect -6460 -3982 -6413 -3918
rect -6349 -3982 -6333 -3918
rect -6460 -3998 -6333 -3982
rect -6460 -4062 -6413 -3998
rect -6349 -4062 -6333 -3998
rect -6460 -4078 -6333 -4062
rect -6460 -4142 -6413 -4078
rect -6349 -4142 -6333 -4078
rect -6460 -4158 -6333 -4142
rect -6460 -4222 -6413 -4158
rect -6349 -4222 -6333 -4158
rect -6460 -4238 -6333 -4222
rect -6460 -4302 -6413 -4238
rect -6349 -4302 -6333 -4238
rect -6460 -4318 -6333 -4302
rect -6460 -4382 -6413 -4318
rect -6349 -4382 -6333 -4318
rect -6460 -4398 -6333 -4382
rect -6460 -4462 -6413 -4398
rect -6349 -4462 -6333 -4398
rect -6460 -4478 -6333 -4462
rect -6460 -4542 -6413 -4478
rect -6349 -4542 -6333 -4478
rect -6460 -4558 -6333 -4542
rect -6460 -4622 -6413 -4558
rect -6349 -4622 -6333 -4558
rect -6460 -4638 -6333 -4622
rect -6460 -4702 -6413 -4638
rect -6349 -4702 -6333 -4638
rect -6460 -4718 -6333 -4702
rect -6460 -4782 -6413 -4718
rect -6349 -4782 -6333 -4718
rect -6460 -4798 -6333 -4782
rect -6460 -4862 -6413 -4798
rect -6349 -4862 -6333 -4798
rect -6460 -4878 -6333 -4862
rect -6460 -4942 -6413 -4878
rect -6349 -4942 -6333 -4878
rect -6460 -4958 -6333 -4942
rect -6460 -5022 -6413 -4958
rect -6349 -5022 -6333 -4958
rect -6460 -5038 -6333 -5022
rect -6460 -5102 -6413 -5038
rect -6349 -5102 -6333 -5038
rect -6460 -5118 -6333 -5102
rect -6460 -5182 -6413 -5118
rect -6349 -5182 -6333 -5118
rect -6460 -5198 -6333 -5182
rect -6460 -5262 -6413 -5198
rect -6349 -5262 -6333 -5198
rect -6460 -5278 -6333 -5262
rect -6460 -5342 -6413 -5278
rect -6349 -5342 -6333 -5278
rect -6460 -5358 -6333 -5342
rect -6460 -5422 -6413 -5358
rect -6349 -5422 -6333 -5358
rect -6460 -5438 -6333 -5422
rect -6460 -5502 -6413 -5438
rect -6349 -5502 -6333 -5438
rect -6460 -5518 -6333 -5502
rect -6460 -5582 -6413 -5518
rect -6349 -5582 -6333 -5518
rect -6460 -5598 -6333 -5582
rect -6460 -5662 -6413 -5598
rect -6349 -5662 -6333 -5598
rect -6460 -5678 -6333 -5662
rect -6460 -5742 -6413 -5678
rect -6349 -5742 -6333 -5678
rect -6460 -5758 -6333 -5742
rect -6460 -5822 -6413 -5758
rect -6349 -5822 -6333 -5758
rect -6460 -5838 -6333 -5822
rect -6460 -5902 -6413 -5838
rect -6349 -5902 -6333 -5838
rect -6460 -5918 -6333 -5902
rect -6460 -5982 -6413 -5918
rect -6349 -5982 -6333 -5918
rect -6460 -5998 -6333 -5982
rect -6460 -6062 -6413 -5998
rect -6349 -6062 -6333 -5998
rect -6460 -6078 -6333 -6062
rect -9580 -6489 -9476 -6111
rect -6460 -6142 -6413 -6078
rect -6349 -6142 -6333 -6078
rect -6170 -198 -248 -189
rect -6170 -6102 -6161 -198
rect -257 -6102 -248 -198
rect -6170 -6111 -248 -6102
rect -141 -222 -94 -158
rect -30 -222 -14 -158
rect 3058 -189 3162 189
rect 6178 158 6225 222
rect 6289 158 6305 222
rect 6468 6102 12390 6111
rect 6468 198 6477 6102
rect 12381 198 12390 6102
rect 6468 189 12390 198
rect 12497 6078 12544 6142
rect 12608 6078 12624 6142
rect 12497 6062 12624 6078
rect 12497 5998 12544 6062
rect 12608 5998 12624 6062
rect 12497 5982 12624 5998
rect 12497 5918 12544 5982
rect 12608 5918 12624 5982
rect 12497 5902 12624 5918
rect 12497 5838 12544 5902
rect 12608 5838 12624 5902
rect 12497 5822 12624 5838
rect 12497 5758 12544 5822
rect 12608 5758 12624 5822
rect 12497 5742 12624 5758
rect 12497 5678 12544 5742
rect 12608 5678 12624 5742
rect 12497 5662 12624 5678
rect 12497 5598 12544 5662
rect 12608 5598 12624 5662
rect 12497 5582 12624 5598
rect 12497 5518 12544 5582
rect 12608 5518 12624 5582
rect 12497 5502 12624 5518
rect 12497 5438 12544 5502
rect 12608 5438 12624 5502
rect 12497 5422 12624 5438
rect 12497 5358 12544 5422
rect 12608 5358 12624 5422
rect 12497 5342 12624 5358
rect 12497 5278 12544 5342
rect 12608 5278 12624 5342
rect 12497 5262 12624 5278
rect 12497 5198 12544 5262
rect 12608 5198 12624 5262
rect 12497 5182 12624 5198
rect 12497 5118 12544 5182
rect 12608 5118 12624 5182
rect 12497 5102 12624 5118
rect 12497 5038 12544 5102
rect 12608 5038 12624 5102
rect 12497 5022 12624 5038
rect 12497 4958 12544 5022
rect 12608 4958 12624 5022
rect 12497 4942 12624 4958
rect 12497 4878 12544 4942
rect 12608 4878 12624 4942
rect 12497 4862 12624 4878
rect 12497 4798 12544 4862
rect 12608 4798 12624 4862
rect 12497 4782 12624 4798
rect 12497 4718 12544 4782
rect 12608 4718 12624 4782
rect 12497 4702 12624 4718
rect 12497 4638 12544 4702
rect 12608 4638 12624 4702
rect 12497 4622 12624 4638
rect 12497 4558 12544 4622
rect 12608 4558 12624 4622
rect 12497 4542 12624 4558
rect 12497 4478 12544 4542
rect 12608 4478 12624 4542
rect 12497 4462 12624 4478
rect 12497 4398 12544 4462
rect 12608 4398 12624 4462
rect 12497 4382 12624 4398
rect 12497 4318 12544 4382
rect 12608 4318 12624 4382
rect 12497 4302 12624 4318
rect 12497 4238 12544 4302
rect 12608 4238 12624 4302
rect 12497 4222 12624 4238
rect 12497 4158 12544 4222
rect 12608 4158 12624 4222
rect 12497 4142 12624 4158
rect 12497 4078 12544 4142
rect 12608 4078 12624 4142
rect 12497 4062 12624 4078
rect 12497 3998 12544 4062
rect 12608 3998 12624 4062
rect 12497 3982 12624 3998
rect 12497 3918 12544 3982
rect 12608 3918 12624 3982
rect 12497 3902 12624 3918
rect 12497 3838 12544 3902
rect 12608 3838 12624 3902
rect 12497 3822 12624 3838
rect 12497 3758 12544 3822
rect 12608 3758 12624 3822
rect 12497 3742 12624 3758
rect 12497 3678 12544 3742
rect 12608 3678 12624 3742
rect 12497 3662 12624 3678
rect 12497 3598 12544 3662
rect 12608 3598 12624 3662
rect 12497 3582 12624 3598
rect 12497 3518 12544 3582
rect 12608 3518 12624 3582
rect 12497 3502 12624 3518
rect 12497 3438 12544 3502
rect 12608 3438 12624 3502
rect 12497 3422 12624 3438
rect 12497 3358 12544 3422
rect 12608 3358 12624 3422
rect 12497 3342 12624 3358
rect 12497 3278 12544 3342
rect 12608 3278 12624 3342
rect 12497 3262 12624 3278
rect 12497 3198 12544 3262
rect 12608 3198 12624 3262
rect 12497 3182 12624 3198
rect 12497 3118 12544 3182
rect 12608 3118 12624 3182
rect 12497 3102 12624 3118
rect 12497 3038 12544 3102
rect 12608 3038 12624 3102
rect 12497 3022 12624 3038
rect 12497 2958 12544 3022
rect 12608 2958 12624 3022
rect 12497 2942 12624 2958
rect 12497 2878 12544 2942
rect 12608 2878 12624 2942
rect 12497 2862 12624 2878
rect 12497 2798 12544 2862
rect 12608 2798 12624 2862
rect 12497 2782 12624 2798
rect 12497 2718 12544 2782
rect 12608 2718 12624 2782
rect 12497 2702 12624 2718
rect 12497 2638 12544 2702
rect 12608 2638 12624 2702
rect 12497 2622 12624 2638
rect 12497 2558 12544 2622
rect 12608 2558 12624 2622
rect 12497 2542 12624 2558
rect 12497 2478 12544 2542
rect 12608 2478 12624 2542
rect 12497 2462 12624 2478
rect 12497 2398 12544 2462
rect 12608 2398 12624 2462
rect 12497 2382 12624 2398
rect 12497 2318 12544 2382
rect 12608 2318 12624 2382
rect 12497 2302 12624 2318
rect 12497 2238 12544 2302
rect 12608 2238 12624 2302
rect 12497 2222 12624 2238
rect 12497 2158 12544 2222
rect 12608 2158 12624 2222
rect 12497 2142 12624 2158
rect 12497 2078 12544 2142
rect 12608 2078 12624 2142
rect 12497 2062 12624 2078
rect 12497 1998 12544 2062
rect 12608 1998 12624 2062
rect 12497 1982 12624 1998
rect 12497 1918 12544 1982
rect 12608 1918 12624 1982
rect 12497 1902 12624 1918
rect 12497 1838 12544 1902
rect 12608 1838 12624 1902
rect 12497 1822 12624 1838
rect 12497 1758 12544 1822
rect 12608 1758 12624 1822
rect 12497 1742 12624 1758
rect 12497 1678 12544 1742
rect 12608 1678 12624 1742
rect 12497 1662 12624 1678
rect 12497 1598 12544 1662
rect 12608 1598 12624 1662
rect 12497 1582 12624 1598
rect 12497 1518 12544 1582
rect 12608 1518 12624 1582
rect 12497 1502 12624 1518
rect 12497 1438 12544 1502
rect 12608 1438 12624 1502
rect 12497 1422 12624 1438
rect 12497 1358 12544 1422
rect 12608 1358 12624 1422
rect 12497 1342 12624 1358
rect 12497 1278 12544 1342
rect 12608 1278 12624 1342
rect 12497 1262 12624 1278
rect 12497 1198 12544 1262
rect 12608 1198 12624 1262
rect 12497 1182 12624 1198
rect 12497 1118 12544 1182
rect 12608 1118 12624 1182
rect 12497 1102 12624 1118
rect 12497 1038 12544 1102
rect 12608 1038 12624 1102
rect 12497 1022 12624 1038
rect 12497 958 12544 1022
rect 12608 958 12624 1022
rect 12497 942 12624 958
rect 12497 878 12544 942
rect 12608 878 12624 942
rect 12497 862 12624 878
rect 12497 798 12544 862
rect 12608 798 12624 862
rect 12497 782 12624 798
rect 12497 718 12544 782
rect 12608 718 12624 782
rect 12497 702 12624 718
rect 12497 638 12544 702
rect 12608 638 12624 702
rect 12497 622 12624 638
rect 12497 558 12544 622
rect 12608 558 12624 622
rect 12497 542 12624 558
rect 12497 478 12544 542
rect 12608 478 12624 542
rect 12497 462 12624 478
rect 12497 398 12544 462
rect 12608 398 12624 462
rect 12497 382 12624 398
rect 12497 318 12544 382
rect 12608 318 12624 382
rect 12497 302 12624 318
rect 12497 238 12544 302
rect 12608 238 12624 302
rect 12497 222 12624 238
rect 6178 142 6305 158
rect 6178 78 6225 142
rect 6289 78 6305 142
rect 6178 62 6305 78
rect 6178 -62 6282 62
rect 6178 -78 6305 -62
rect 6178 -142 6225 -78
rect 6289 -142 6305 -78
rect 6178 -158 6305 -142
rect -141 -238 -14 -222
rect -141 -302 -94 -238
rect -30 -302 -14 -238
rect -141 -318 -14 -302
rect -141 -382 -94 -318
rect -30 -382 -14 -318
rect -141 -398 -14 -382
rect -141 -462 -94 -398
rect -30 -462 -14 -398
rect -141 -478 -14 -462
rect -141 -542 -94 -478
rect -30 -542 -14 -478
rect -141 -558 -14 -542
rect -141 -622 -94 -558
rect -30 -622 -14 -558
rect -141 -638 -14 -622
rect -141 -702 -94 -638
rect -30 -702 -14 -638
rect -141 -718 -14 -702
rect -141 -782 -94 -718
rect -30 -782 -14 -718
rect -141 -798 -14 -782
rect -141 -862 -94 -798
rect -30 -862 -14 -798
rect -141 -878 -14 -862
rect -141 -942 -94 -878
rect -30 -942 -14 -878
rect -141 -958 -14 -942
rect -141 -1022 -94 -958
rect -30 -1022 -14 -958
rect -141 -1038 -14 -1022
rect -141 -1102 -94 -1038
rect -30 -1102 -14 -1038
rect -141 -1118 -14 -1102
rect -141 -1182 -94 -1118
rect -30 -1182 -14 -1118
rect -141 -1198 -14 -1182
rect -141 -1262 -94 -1198
rect -30 -1262 -14 -1198
rect -141 -1278 -14 -1262
rect -141 -1342 -94 -1278
rect -30 -1342 -14 -1278
rect -141 -1358 -14 -1342
rect -141 -1422 -94 -1358
rect -30 -1422 -14 -1358
rect -141 -1438 -14 -1422
rect -141 -1502 -94 -1438
rect -30 -1502 -14 -1438
rect -141 -1518 -14 -1502
rect -141 -1582 -94 -1518
rect -30 -1582 -14 -1518
rect -141 -1598 -14 -1582
rect -141 -1662 -94 -1598
rect -30 -1662 -14 -1598
rect -141 -1678 -14 -1662
rect -141 -1742 -94 -1678
rect -30 -1742 -14 -1678
rect -141 -1758 -14 -1742
rect -141 -1822 -94 -1758
rect -30 -1822 -14 -1758
rect -141 -1838 -14 -1822
rect -141 -1902 -94 -1838
rect -30 -1902 -14 -1838
rect -141 -1918 -14 -1902
rect -141 -1982 -94 -1918
rect -30 -1982 -14 -1918
rect -141 -1998 -14 -1982
rect -141 -2062 -94 -1998
rect -30 -2062 -14 -1998
rect -141 -2078 -14 -2062
rect -141 -2142 -94 -2078
rect -30 -2142 -14 -2078
rect -141 -2158 -14 -2142
rect -141 -2222 -94 -2158
rect -30 -2222 -14 -2158
rect -141 -2238 -14 -2222
rect -141 -2302 -94 -2238
rect -30 -2302 -14 -2238
rect -141 -2318 -14 -2302
rect -141 -2382 -94 -2318
rect -30 -2382 -14 -2318
rect -141 -2398 -14 -2382
rect -141 -2462 -94 -2398
rect -30 -2462 -14 -2398
rect -141 -2478 -14 -2462
rect -141 -2542 -94 -2478
rect -30 -2542 -14 -2478
rect -141 -2558 -14 -2542
rect -141 -2622 -94 -2558
rect -30 -2622 -14 -2558
rect -141 -2638 -14 -2622
rect -141 -2702 -94 -2638
rect -30 -2702 -14 -2638
rect -141 -2718 -14 -2702
rect -141 -2782 -94 -2718
rect -30 -2782 -14 -2718
rect -141 -2798 -14 -2782
rect -141 -2862 -94 -2798
rect -30 -2862 -14 -2798
rect -141 -2878 -14 -2862
rect -141 -2942 -94 -2878
rect -30 -2942 -14 -2878
rect -141 -2958 -14 -2942
rect -141 -3022 -94 -2958
rect -30 -3022 -14 -2958
rect -141 -3038 -14 -3022
rect -141 -3102 -94 -3038
rect -30 -3102 -14 -3038
rect -141 -3118 -14 -3102
rect -141 -3182 -94 -3118
rect -30 -3182 -14 -3118
rect -141 -3198 -14 -3182
rect -141 -3262 -94 -3198
rect -30 -3262 -14 -3198
rect -141 -3278 -14 -3262
rect -141 -3342 -94 -3278
rect -30 -3342 -14 -3278
rect -141 -3358 -14 -3342
rect -141 -3422 -94 -3358
rect -30 -3422 -14 -3358
rect -141 -3438 -14 -3422
rect -141 -3502 -94 -3438
rect -30 -3502 -14 -3438
rect -141 -3518 -14 -3502
rect -141 -3582 -94 -3518
rect -30 -3582 -14 -3518
rect -141 -3598 -14 -3582
rect -141 -3662 -94 -3598
rect -30 -3662 -14 -3598
rect -141 -3678 -14 -3662
rect -141 -3742 -94 -3678
rect -30 -3742 -14 -3678
rect -141 -3758 -14 -3742
rect -141 -3822 -94 -3758
rect -30 -3822 -14 -3758
rect -141 -3838 -14 -3822
rect -141 -3902 -94 -3838
rect -30 -3902 -14 -3838
rect -141 -3918 -14 -3902
rect -141 -3982 -94 -3918
rect -30 -3982 -14 -3918
rect -141 -3998 -14 -3982
rect -141 -4062 -94 -3998
rect -30 -4062 -14 -3998
rect -141 -4078 -14 -4062
rect -141 -4142 -94 -4078
rect -30 -4142 -14 -4078
rect -141 -4158 -14 -4142
rect -141 -4222 -94 -4158
rect -30 -4222 -14 -4158
rect -141 -4238 -14 -4222
rect -141 -4302 -94 -4238
rect -30 -4302 -14 -4238
rect -141 -4318 -14 -4302
rect -141 -4382 -94 -4318
rect -30 -4382 -14 -4318
rect -141 -4398 -14 -4382
rect -141 -4462 -94 -4398
rect -30 -4462 -14 -4398
rect -141 -4478 -14 -4462
rect -141 -4542 -94 -4478
rect -30 -4542 -14 -4478
rect -141 -4558 -14 -4542
rect -141 -4622 -94 -4558
rect -30 -4622 -14 -4558
rect -141 -4638 -14 -4622
rect -141 -4702 -94 -4638
rect -30 -4702 -14 -4638
rect -141 -4718 -14 -4702
rect -141 -4782 -94 -4718
rect -30 -4782 -14 -4718
rect -141 -4798 -14 -4782
rect -141 -4862 -94 -4798
rect -30 -4862 -14 -4798
rect -141 -4878 -14 -4862
rect -141 -4942 -94 -4878
rect -30 -4942 -14 -4878
rect -141 -4958 -14 -4942
rect -141 -5022 -94 -4958
rect -30 -5022 -14 -4958
rect -141 -5038 -14 -5022
rect -141 -5102 -94 -5038
rect -30 -5102 -14 -5038
rect -141 -5118 -14 -5102
rect -141 -5182 -94 -5118
rect -30 -5182 -14 -5118
rect -141 -5198 -14 -5182
rect -141 -5262 -94 -5198
rect -30 -5262 -14 -5198
rect -141 -5278 -14 -5262
rect -141 -5342 -94 -5278
rect -30 -5342 -14 -5278
rect -141 -5358 -14 -5342
rect -141 -5422 -94 -5358
rect -30 -5422 -14 -5358
rect -141 -5438 -14 -5422
rect -141 -5502 -94 -5438
rect -30 -5502 -14 -5438
rect -141 -5518 -14 -5502
rect -141 -5582 -94 -5518
rect -30 -5582 -14 -5518
rect -141 -5598 -14 -5582
rect -141 -5662 -94 -5598
rect -30 -5662 -14 -5598
rect -141 -5678 -14 -5662
rect -141 -5742 -94 -5678
rect -30 -5742 -14 -5678
rect -141 -5758 -14 -5742
rect -141 -5822 -94 -5758
rect -30 -5822 -14 -5758
rect -141 -5838 -14 -5822
rect -141 -5902 -94 -5838
rect -30 -5902 -14 -5838
rect -141 -5918 -14 -5902
rect -141 -5982 -94 -5918
rect -30 -5982 -14 -5918
rect -141 -5998 -14 -5982
rect -141 -6062 -94 -5998
rect -30 -6062 -14 -5998
rect -141 -6078 -14 -6062
rect -6460 -6158 -6333 -6142
rect -6460 -6222 -6413 -6158
rect -6349 -6222 -6333 -6158
rect -6460 -6238 -6333 -6222
rect -6460 -6362 -6356 -6238
rect -6460 -6378 -6333 -6362
rect -6460 -6442 -6413 -6378
rect -6349 -6442 -6333 -6378
rect -6460 -6458 -6333 -6442
rect -12489 -6498 -6567 -6489
rect -12489 -12402 -12480 -6498
rect -6576 -12402 -6567 -6498
rect -12489 -12411 -6567 -12402
rect -6460 -6522 -6413 -6458
rect -6349 -6522 -6333 -6458
rect -3261 -6489 -3157 -6111
rect -141 -6142 -94 -6078
rect -30 -6142 -14 -6078
rect 149 -198 6071 -189
rect 149 -6102 158 -198
rect 6062 -6102 6071 -198
rect 149 -6111 6071 -6102
rect 6178 -222 6225 -158
rect 6289 -222 6305 -158
rect 9377 -189 9481 189
rect 12497 158 12544 222
rect 12608 158 12624 222
rect 12497 142 12624 158
rect 12497 78 12544 142
rect 12608 78 12624 142
rect 12497 62 12624 78
rect 12497 -62 12601 62
rect 12497 -78 12624 -62
rect 12497 -142 12544 -78
rect 12608 -142 12624 -78
rect 12497 -158 12624 -142
rect 6178 -238 6305 -222
rect 6178 -302 6225 -238
rect 6289 -302 6305 -238
rect 6178 -318 6305 -302
rect 6178 -382 6225 -318
rect 6289 -382 6305 -318
rect 6178 -398 6305 -382
rect 6178 -462 6225 -398
rect 6289 -462 6305 -398
rect 6178 -478 6305 -462
rect 6178 -542 6225 -478
rect 6289 -542 6305 -478
rect 6178 -558 6305 -542
rect 6178 -622 6225 -558
rect 6289 -622 6305 -558
rect 6178 -638 6305 -622
rect 6178 -702 6225 -638
rect 6289 -702 6305 -638
rect 6178 -718 6305 -702
rect 6178 -782 6225 -718
rect 6289 -782 6305 -718
rect 6178 -798 6305 -782
rect 6178 -862 6225 -798
rect 6289 -862 6305 -798
rect 6178 -878 6305 -862
rect 6178 -942 6225 -878
rect 6289 -942 6305 -878
rect 6178 -958 6305 -942
rect 6178 -1022 6225 -958
rect 6289 -1022 6305 -958
rect 6178 -1038 6305 -1022
rect 6178 -1102 6225 -1038
rect 6289 -1102 6305 -1038
rect 6178 -1118 6305 -1102
rect 6178 -1182 6225 -1118
rect 6289 -1182 6305 -1118
rect 6178 -1198 6305 -1182
rect 6178 -1262 6225 -1198
rect 6289 -1262 6305 -1198
rect 6178 -1278 6305 -1262
rect 6178 -1342 6225 -1278
rect 6289 -1342 6305 -1278
rect 6178 -1358 6305 -1342
rect 6178 -1422 6225 -1358
rect 6289 -1422 6305 -1358
rect 6178 -1438 6305 -1422
rect 6178 -1502 6225 -1438
rect 6289 -1502 6305 -1438
rect 6178 -1518 6305 -1502
rect 6178 -1582 6225 -1518
rect 6289 -1582 6305 -1518
rect 6178 -1598 6305 -1582
rect 6178 -1662 6225 -1598
rect 6289 -1662 6305 -1598
rect 6178 -1678 6305 -1662
rect 6178 -1742 6225 -1678
rect 6289 -1742 6305 -1678
rect 6178 -1758 6305 -1742
rect 6178 -1822 6225 -1758
rect 6289 -1822 6305 -1758
rect 6178 -1838 6305 -1822
rect 6178 -1902 6225 -1838
rect 6289 -1902 6305 -1838
rect 6178 -1918 6305 -1902
rect 6178 -1982 6225 -1918
rect 6289 -1982 6305 -1918
rect 6178 -1998 6305 -1982
rect 6178 -2062 6225 -1998
rect 6289 -2062 6305 -1998
rect 6178 -2078 6305 -2062
rect 6178 -2142 6225 -2078
rect 6289 -2142 6305 -2078
rect 6178 -2158 6305 -2142
rect 6178 -2222 6225 -2158
rect 6289 -2222 6305 -2158
rect 6178 -2238 6305 -2222
rect 6178 -2302 6225 -2238
rect 6289 -2302 6305 -2238
rect 6178 -2318 6305 -2302
rect 6178 -2382 6225 -2318
rect 6289 -2382 6305 -2318
rect 6178 -2398 6305 -2382
rect 6178 -2462 6225 -2398
rect 6289 -2462 6305 -2398
rect 6178 -2478 6305 -2462
rect 6178 -2542 6225 -2478
rect 6289 -2542 6305 -2478
rect 6178 -2558 6305 -2542
rect 6178 -2622 6225 -2558
rect 6289 -2622 6305 -2558
rect 6178 -2638 6305 -2622
rect 6178 -2702 6225 -2638
rect 6289 -2702 6305 -2638
rect 6178 -2718 6305 -2702
rect 6178 -2782 6225 -2718
rect 6289 -2782 6305 -2718
rect 6178 -2798 6305 -2782
rect 6178 -2862 6225 -2798
rect 6289 -2862 6305 -2798
rect 6178 -2878 6305 -2862
rect 6178 -2942 6225 -2878
rect 6289 -2942 6305 -2878
rect 6178 -2958 6305 -2942
rect 6178 -3022 6225 -2958
rect 6289 -3022 6305 -2958
rect 6178 -3038 6305 -3022
rect 6178 -3102 6225 -3038
rect 6289 -3102 6305 -3038
rect 6178 -3118 6305 -3102
rect 6178 -3182 6225 -3118
rect 6289 -3182 6305 -3118
rect 6178 -3198 6305 -3182
rect 6178 -3262 6225 -3198
rect 6289 -3262 6305 -3198
rect 6178 -3278 6305 -3262
rect 6178 -3342 6225 -3278
rect 6289 -3342 6305 -3278
rect 6178 -3358 6305 -3342
rect 6178 -3422 6225 -3358
rect 6289 -3422 6305 -3358
rect 6178 -3438 6305 -3422
rect 6178 -3502 6225 -3438
rect 6289 -3502 6305 -3438
rect 6178 -3518 6305 -3502
rect 6178 -3582 6225 -3518
rect 6289 -3582 6305 -3518
rect 6178 -3598 6305 -3582
rect 6178 -3662 6225 -3598
rect 6289 -3662 6305 -3598
rect 6178 -3678 6305 -3662
rect 6178 -3742 6225 -3678
rect 6289 -3742 6305 -3678
rect 6178 -3758 6305 -3742
rect 6178 -3822 6225 -3758
rect 6289 -3822 6305 -3758
rect 6178 -3838 6305 -3822
rect 6178 -3902 6225 -3838
rect 6289 -3902 6305 -3838
rect 6178 -3918 6305 -3902
rect 6178 -3982 6225 -3918
rect 6289 -3982 6305 -3918
rect 6178 -3998 6305 -3982
rect 6178 -4062 6225 -3998
rect 6289 -4062 6305 -3998
rect 6178 -4078 6305 -4062
rect 6178 -4142 6225 -4078
rect 6289 -4142 6305 -4078
rect 6178 -4158 6305 -4142
rect 6178 -4222 6225 -4158
rect 6289 -4222 6305 -4158
rect 6178 -4238 6305 -4222
rect 6178 -4302 6225 -4238
rect 6289 -4302 6305 -4238
rect 6178 -4318 6305 -4302
rect 6178 -4382 6225 -4318
rect 6289 -4382 6305 -4318
rect 6178 -4398 6305 -4382
rect 6178 -4462 6225 -4398
rect 6289 -4462 6305 -4398
rect 6178 -4478 6305 -4462
rect 6178 -4542 6225 -4478
rect 6289 -4542 6305 -4478
rect 6178 -4558 6305 -4542
rect 6178 -4622 6225 -4558
rect 6289 -4622 6305 -4558
rect 6178 -4638 6305 -4622
rect 6178 -4702 6225 -4638
rect 6289 -4702 6305 -4638
rect 6178 -4718 6305 -4702
rect 6178 -4782 6225 -4718
rect 6289 -4782 6305 -4718
rect 6178 -4798 6305 -4782
rect 6178 -4862 6225 -4798
rect 6289 -4862 6305 -4798
rect 6178 -4878 6305 -4862
rect 6178 -4942 6225 -4878
rect 6289 -4942 6305 -4878
rect 6178 -4958 6305 -4942
rect 6178 -5022 6225 -4958
rect 6289 -5022 6305 -4958
rect 6178 -5038 6305 -5022
rect 6178 -5102 6225 -5038
rect 6289 -5102 6305 -5038
rect 6178 -5118 6305 -5102
rect 6178 -5182 6225 -5118
rect 6289 -5182 6305 -5118
rect 6178 -5198 6305 -5182
rect 6178 -5262 6225 -5198
rect 6289 -5262 6305 -5198
rect 6178 -5278 6305 -5262
rect 6178 -5342 6225 -5278
rect 6289 -5342 6305 -5278
rect 6178 -5358 6305 -5342
rect 6178 -5422 6225 -5358
rect 6289 -5422 6305 -5358
rect 6178 -5438 6305 -5422
rect 6178 -5502 6225 -5438
rect 6289 -5502 6305 -5438
rect 6178 -5518 6305 -5502
rect 6178 -5582 6225 -5518
rect 6289 -5582 6305 -5518
rect 6178 -5598 6305 -5582
rect 6178 -5662 6225 -5598
rect 6289 -5662 6305 -5598
rect 6178 -5678 6305 -5662
rect 6178 -5742 6225 -5678
rect 6289 -5742 6305 -5678
rect 6178 -5758 6305 -5742
rect 6178 -5822 6225 -5758
rect 6289 -5822 6305 -5758
rect 6178 -5838 6305 -5822
rect 6178 -5902 6225 -5838
rect 6289 -5902 6305 -5838
rect 6178 -5918 6305 -5902
rect 6178 -5982 6225 -5918
rect 6289 -5982 6305 -5918
rect 6178 -5998 6305 -5982
rect 6178 -6062 6225 -5998
rect 6289 -6062 6305 -5998
rect 6178 -6078 6305 -6062
rect -141 -6158 -14 -6142
rect -141 -6222 -94 -6158
rect -30 -6222 -14 -6158
rect -141 -6238 -14 -6222
rect -141 -6362 -37 -6238
rect -141 -6378 -14 -6362
rect -141 -6442 -94 -6378
rect -30 -6442 -14 -6378
rect -141 -6458 -14 -6442
rect -6460 -6538 -6333 -6522
rect -6460 -6602 -6413 -6538
rect -6349 -6602 -6333 -6538
rect -6460 -6618 -6333 -6602
rect -6460 -6682 -6413 -6618
rect -6349 -6682 -6333 -6618
rect -6460 -6698 -6333 -6682
rect -6460 -6762 -6413 -6698
rect -6349 -6762 -6333 -6698
rect -6460 -6778 -6333 -6762
rect -6460 -6842 -6413 -6778
rect -6349 -6842 -6333 -6778
rect -6460 -6858 -6333 -6842
rect -6460 -6922 -6413 -6858
rect -6349 -6922 -6333 -6858
rect -6460 -6938 -6333 -6922
rect -6460 -7002 -6413 -6938
rect -6349 -7002 -6333 -6938
rect -6460 -7018 -6333 -7002
rect -6460 -7082 -6413 -7018
rect -6349 -7082 -6333 -7018
rect -6460 -7098 -6333 -7082
rect -6460 -7162 -6413 -7098
rect -6349 -7162 -6333 -7098
rect -6460 -7178 -6333 -7162
rect -6460 -7242 -6413 -7178
rect -6349 -7242 -6333 -7178
rect -6460 -7258 -6333 -7242
rect -6460 -7322 -6413 -7258
rect -6349 -7322 -6333 -7258
rect -6460 -7338 -6333 -7322
rect -6460 -7402 -6413 -7338
rect -6349 -7402 -6333 -7338
rect -6460 -7418 -6333 -7402
rect -6460 -7482 -6413 -7418
rect -6349 -7482 -6333 -7418
rect -6460 -7498 -6333 -7482
rect -6460 -7562 -6413 -7498
rect -6349 -7562 -6333 -7498
rect -6460 -7578 -6333 -7562
rect -6460 -7642 -6413 -7578
rect -6349 -7642 -6333 -7578
rect -6460 -7658 -6333 -7642
rect -6460 -7722 -6413 -7658
rect -6349 -7722 -6333 -7658
rect -6460 -7738 -6333 -7722
rect -6460 -7802 -6413 -7738
rect -6349 -7802 -6333 -7738
rect -6460 -7818 -6333 -7802
rect -6460 -7882 -6413 -7818
rect -6349 -7882 -6333 -7818
rect -6460 -7898 -6333 -7882
rect -6460 -7962 -6413 -7898
rect -6349 -7962 -6333 -7898
rect -6460 -7978 -6333 -7962
rect -6460 -8042 -6413 -7978
rect -6349 -8042 -6333 -7978
rect -6460 -8058 -6333 -8042
rect -6460 -8122 -6413 -8058
rect -6349 -8122 -6333 -8058
rect -6460 -8138 -6333 -8122
rect -6460 -8202 -6413 -8138
rect -6349 -8202 -6333 -8138
rect -6460 -8218 -6333 -8202
rect -6460 -8282 -6413 -8218
rect -6349 -8282 -6333 -8218
rect -6460 -8298 -6333 -8282
rect -6460 -8362 -6413 -8298
rect -6349 -8362 -6333 -8298
rect -6460 -8378 -6333 -8362
rect -6460 -8442 -6413 -8378
rect -6349 -8442 -6333 -8378
rect -6460 -8458 -6333 -8442
rect -6460 -8522 -6413 -8458
rect -6349 -8522 -6333 -8458
rect -6460 -8538 -6333 -8522
rect -6460 -8602 -6413 -8538
rect -6349 -8602 -6333 -8538
rect -6460 -8618 -6333 -8602
rect -6460 -8682 -6413 -8618
rect -6349 -8682 -6333 -8618
rect -6460 -8698 -6333 -8682
rect -6460 -8762 -6413 -8698
rect -6349 -8762 -6333 -8698
rect -6460 -8778 -6333 -8762
rect -6460 -8842 -6413 -8778
rect -6349 -8842 -6333 -8778
rect -6460 -8858 -6333 -8842
rect -6460 -8922 -6413 -8858
rect -6349 -8922 -6333 -8858
rect -6460 -8938 -6333 -8922
rect -6460 -9002 -6413 -8938
rect -6349 -9002 -6333 -8938
rect -6460 -9018 -6333 -9002
rect -6460 -9082 -6413 -9018
rect -6349 -9082 -6333 -9018
rect -6460 -9098 -6333 -9082
rect -6460 -9162 -6413 -9098
rect -6349 -9162 -6333 -9098
rect -6460 -9178 -6333 -9162
rect -6460 -9242 -6413 -9178
rect -6349 -9242 -6333 -9178
rect -6460 -9258 -6333 -9242
rect -6460 -9322 -6413 -9258
rect -6349 -9322 -6333 -9258
rect -6460 -9338 -6333 -9322
rect -6460 -9402 -6413 -9338
rect -6349 -9402 -6333 -9338
rect -6460 -9418 -6333 -9402
rect -6460 -9482 -6413 -9418
rect -6349 -9482 -6333 -9418
rect -6460 -9498 -6333 -9482
rect -6460 -9562 -6413 -9498
rect -6349 -9562 -6333 -9498
rect -6460 -9578 -6333 -9562
rect -6460 -9642 -6413 -9578
rect -6349 -9642 -6333 -9578
rect -6460 -9658 -6333 -9642
rect -6460 -9722 -6413 -9658
rect -6349 -9722 -6333 -9658
rect -6460 -9738 -6333 -9722
rect -6460 -9802 -6413 -9738
rect -6349 -9802 -6333 -9738
rect -6460 -9818 -6333 -9802
rect -6460 -9882 -6413 -9818
rect -6349 -9882 -6333 -9818
rect -6460 -9898 -6333 -9882
rect -6460 -9962 -6413 -9898
rect -6349 -9962 -6333 -9898
rect -6460 -9978 -6333 -9962
rect -6460 -10042 -6413 -9978
rect -6349 -10042 -6333 -9978
rect -6460 -10058 -6333 -10042
rect -6460 -10122 -6413 -10058
rect -6349 -10122 -6333 -10058
rect -6460 -10138 -6333 -10122
rect -6460 -10202 -6413 -10138
rect -6349 -10202 -6333 -10138
rect -6460 -10218 -6333 -10202
rect -6460 -10282 -6413 -10218
rect -6349 -10282 -6333 -10218
rect -6460 -10298 -6333 -10282
rect -6460 -10362 -6413 -10298
rect -6349 -10362 -6333 -10298
rect -6460 -10378 -6333 -10362
rect -6460 -10442 -6413 -10378
rect -6349 -10442 -6333 -10378
rect -6460 -10458 -6333 -10442
rect -6460 -10522 -6413 -10458
rect -6349 -10522 -6333 -10458
rect -6460 -10538 -6333 -10522
rect -6460 -10602 -6413 -10538
rect -6349 -10602 -6333 -10538
rect -6460 -10618 -6333 -10602
rect -6460 -10682 -6413 -10618
rect -6349 -10682 -6333 -10618
rect -6460 -10698 -6333 -10682
rect -6460 -10762 -6413 -10698
rect -6349 -10762 -6333 -10698
rect -6460 -10778 -6333 -10762
rect -6460 -10842 -6413 -10778
rect -6349 -10842 -6333 -10778
rect -6460 -10858 -6333 -10842
rect -6460 -10922 -6413 -10858
rect -6349 -10922 -6333 -10858
rect -6460 -10938 -6333 -10922
rect -6460 -11002 -6413 -10938
rect -6349 -11002 -6333 -10938
rect -6460 -11018 -6333 -11002
rect -6460 -11082 -6413 -11018
rect -6349 -11082 -6333 -11018
rect -6460 -11098 -6333 -11082
rect -6460 -11162 -6413 -11098
rect -6349 -11162 -6333 -11098
rect -6460 -11178 -6333 -11162
rect -6460 -11242 -6413 -11178
rect -6349 -11242 -6333 -11178
rect -6460 -11258 -6333 -11242
rect -6460 -11322 -6413 -11258
rect -6349 -11322 -6333 -11258
rect -6460 -11338 -6333 -11322
rect -6460 -11402 -6413 -11338
rect -6349 -11402 -6333 -11338
rect -6460 -11418 -6333 -11402
rect -6460 -11482 -6413 -11418
rect -6349 -11482 -6333 -11418
rect -6460 -11498 -6333 -11482
rect -6460 -11562 -6413 -11498
rect -6349 -11562 -6333 -11498
rect -6460 -11578 -6333 -11562
rect -6460 -11642 -6413 -11578
rect -6349 -11642 -6333 -11578
rect -6460 -11658 -6333 -11642
rect -6460 -11722 -6413 -11658
rect -6349 -11722 -6333 -11658
rect -6460 -11738 -6333 -11722
rect -6460 -11802 -6413 -11738
rect -6349 -11802 -6333 -11738
rect -6460 -11818 -6333 -11802
rect -6460 -11882 -6413 -11818
rect -6349 -11882 -6333 -11818
rect -6460 -11898 -6333 -11882
rect -6460 -11962 -6413 -11898
rect -6349 -11962 -6333 -11898
rect -6460 -11978 -6333 -11962
rect -6460 -12042 -6413 -11978
rect -6349 -12042 -6333 -11978
rect -6460 -12058 -6333 -12042
rect -6460 -12122 -6413 -12058
rect -6349 -12122 -6333 -12058
rect -6460 -12138 -6333 -12122
rect -6460 -12202 -6413 -12138
rect -6349 -12202 -6333 -12138
rect -6460 -12218 -6333 -12202
rect -6460 -12282 -6413 -12218
rect -6349 -12282 -6333 -12218
rect -6460 -12298 -6333 -12282
rect -6460 -12362 -6413 -12298
rect -6349 -12362 -6333 -12298
rect -6460 -12378 -6333 -12362
rect -9580 -12600 -9476 -12411
rect -6460 -12442 -6413 -12378
rect -6349 -12442 -6333 -12378
rect -6170 -6498 -248 -6489
rect -6170 -12402 -6161 -6498
rect -257 -12402 -248 -6498
rect -6170 -12411 -248 -12402
rect -141 -6522 -94 -6458
rect -30 -6522 -14 -6458
rect 3058 -6489 3162 -6111
rect 6178 -6142 6225 -6078
rect 6289 -6142 6305 -6078
rect 6468 -198 12390 -189
rect 6468 -6102 6477 -198
rect 12381 -6102 12390 -198
rect 6468 -6111 12390 -6102
rect 12497 -222 12544 -158
rect 12608 -222 12624 -158
rect 12497 -238 12624 -222
rect 12497 -302 12544 -238
rect 12608 -302 12624 -238
rect 12497 -318 12624 -302
rect 12497 -382 12544 -318
rect 12608 -382 12624 -318
rect 12497 -398 12624 -382
rect 12497 -462 12544 -398
rect 12608 -462 12624 -398
rect 12497 -478 12624 -462
rect 12497 -542 12544 -478
rect 12608 -542 12624 -478
rect 12497 -558 12624 -542
rect 12497 -622 12544 -558
rect 12608 -622 12624 -558
rect 12497 -638 12624 -622
rect 12497 -702 12544 -638
rect 12608 -702 12624 -638
rect 12497 -718 12624 -702
rect 12497 -782 12544 -718
rect 12608 -782 12624 -718
rect 12497 -798 12624 -782
rect 12497 -862 12544 -798
rect 12608 -862 12624 -798
rect 12497 -878 12624 -862
rect 12497 -942 12544 -878
rect 12608 -942 12624 -878
rect 12497 -958 12624 -942
rect 12497 -1022 12544 -958
rect 12608 -1022 12624 -958
rect 12497 -1038 12624 -1022
rect 12497 -1102 12544 -1038
rect 12608 -1102 12624 -1038
rect 12497 -1118 12624 -1102
rect 12497 -1182 12544 -1118
rect 12608 -1182 12624 -1118
rect 12497 -1198 12624 -1182
rect 12497 -1262 12544 -1198
rect 12608 -1262 12624 -1198
rect 12497 -1278 12624 -1262
rect 12497 -1342 12544 -1278
rect 12608 -1342 12624 -1278
rect 12497 -1358 12624 -1342
rect 12497 -1422 12544 -1358
rect 12608 -1422 12624 -1358
rect 12497 -1438 12624 -1422
rect 12497 -1502 12544 -1438
rect 12608 -1502 12624 -1438
rect 12497 -1518 12624 -1502
rect 12497 -1582 12544 -1518
rect 12608 -1582 12624 -1518
rect 12497 -1598 12624 -1582
rect 12497 -1662 12544 -1598
rect 12608 -1662 12624 -1598
rect 12497 -1678 12624 -1662
rect 12497 -1742 12544 -1678
rect 12608 -1742 12624 -1678
rect 12497 -1758 12624 -1742
rect 12497 -1822 12544 -1758
rect 12608 -1822 12624 -1758
rect 12497 -1838 12624 -1822
rect 12497 -1902 12544 -1838
rect 12608 -1902 12624 -1838
rect 12497 -1918 12624 -1902
rect 12497 -1982 12544 -1918
rect 12608 -1982 12624 -1918
rect 12497 -1998 12624 -1982
rect 12497 -2062 12544 -1998
rect 12608 -2062 12624 -1998
rect 12497 -2078 12624 -2062
rect 12497 -2142 12544 -2078
rect 12608 -2142 12624 -2078
rect 12497 -2158 12624 -2142
rect 12497 -2222 12544 -2158
rect 12608 -2222 12624 -2158
rect 12497 -2238 12624 -2222
rect 12497 -2302 12544 -2238
rect 12608 -2302 12624 -2238
rect 12497 -2318 12624 -2302
rect 12497 -2382 12544 -2318
rect 12608 -2382 12624 -2318
rect 12497 -2398 12624 -2382
rect 12497 -2462 12544 -2398
rect 12608 -2462 12624 -2398
rect 12497 -2478 12624 -2462
rect 12497 -2542 12544 -2478
rect 12608 -2542 12624 -2478
rect 12497 -2558 12624 -2542
rect 12497 -2622 12544 -2558
rect 12608 -2622 12624 -2558
rect 12497 -2638 12624 -2622
rect 12497 -2702 12544 -2638
rect 12608 -2702 12624 -2638
rect 12497 -2718 12624 -2702
rect 12497 -2782 12544 -2718
rect 12608 -2782 12624 -2718
rect 12497 -2798 12624 -2782
rect 12497 -2862 12544 -2798
rect 12608 -2862 12624 -2798
rect 12497 -2878 12624 -2862
rect 12497 -2942 12544 -2878
rect 12608 -2942 12624 -2878
rect 12497 -2958 12624 -2942
rect 12497 -3022 12544 -2958
rect 12608 -3022 12624 -2958
rect 12497 -3038 12624 -3022
rect 12497 -3102 12544 -3038
rect 12608 -3102 12624 -3038
rect 12497 -3118 12624 -3102
rect 12497 -3182 12544 -3118
rect 12608 -3182 12624 -3118
rect 12497 -3198 12624 -3182
rect 12497 -3262 12544 -3198
rect 12608 -3262 12624 -3198
rect 12497 -3278 12624 -3262
rect 12497 -3342 12544 -3278
rect 12608 -3342 12624 -3278
rect 12497 -3358 12624 -3342
rect 12497 -3422 12544 -3358
rect 12608 -3422 12624 -3358
rect 12497 -3438 12624 -3422
rect 12497 -3502 12544 -3438
rect 12608 -3502 12624 -3438
rect 12497 -3518 12624 -3502
rect 12497 -3582 12544 -3518
rect 12608 -3582 12624 -3518
rect 12497 -3598 12624 -3582
rect 12497 -3662 12544 -3598
rect 12608 -3662 12624 -3598
rect 12497 -3678 12624 -3662
rect 12497 -3742 12544 -3678
rect 12608 -3742 12624 -3678
rect 12497 -3758 12624 -3742
rect 12497 -3822 12544 -3758
rect 12608 -3822 12624 -3758
rect 12497 -3838 12624 -3822
rect 12497 -3902 12544 -3838
rect 12608 -3902 12624 -3838
rect 12497 -3918 12624 -3902
rect 12497 -3982 12544 -3918
rect 12608 -3982 12624 -3918
rect 12497 -3998 12624 -3982
rect 12497 -4062 12544 -3998
rect 12608 -4062 12624 -3998
rect 12497 -4078 12624 -4062
rect 12497 -4142 12544 -4078
rect 12608 -4142 12624 -4078
rect 12497 -4158 12624 -4142
rect 12497 -4222 12544 -4158
rect 12608 -4222 12624 -4158
rect 12497 -4238 12624 -4222
rect 12497 -4302 12544 -4238
rect 12608 -4302 12624 -4238
rect 12497 -4318 12624 -4302
rect 12497 -4382 12544 -4318
rect 12608 -4382 12624 -4318
rect 12497 -4398 12624 -4382
rect 12497 -4462 12544 -4398
rect 12608 -4462 12624 -4398
rect 12497 -4478 12624 -4462
rect 12497 -4542 12544 -4478
rect 12608 -4542 12624 -4478
rect 12497 -4558 12624 -4542
rect 12497 -4622 12544 -4558
rect 12608 -4622 12624 -4558
rect 12497 -4638 12624 -4622
rect 12497 -4702 12544 -4638
rect 12608 -4702 12624 -4638
rect 12497 -4718 12624 -4702
rect 12497 -4782 12544 -4718
rect 12608 -4782 12624 -4718
rect 12497 -4798 12624 -4782
rect 12497 -4862 12544 -4798
rect 12608 -4862 12624 -4798
rect 12497 -4878 12624 -4862
rect 12497 -4942 12544 -4878
rect 12608 -4942 12624 -4878
rect 12497 -4958 12624 -4942
rect 12497 -5022 12544 -4958
rect 12608 -5022 12624 -4958
rect 12497 -5038 12624 -5022
rect 12497 -5102 12544 -5038
rect 12608 -5102 12624 -5038
rect 12497 -5118 12624 -5102
rect 12497 -5182 12544 -5118
rect 12608 -5182 12624 -5118
rect 12497 -5198 12624 -5182
rect 12497 -5262 12544 -5198
rect 12608 -5262 12624 -5198
rect 12497 -5278 12624 -5262
rect 12497 -5342 12544 -5278
rect 12608 -5342 12624 -5278
rect 12497 -5358 12624 -5342
rect 12497 -5422 12544 -5358
rect 12608 -5422 12624 -5358
rect 12497 -5438 12624 -5422
rect 12497 -5502 12544 -5438
rect 12608 -5502 12624 -5438
rect 12497 -5518 12624 -5502
rect 12497 -5582 12544 -5518
rect 12608 -5582 12624 -5518
rect 12497 -5598 12624 -5582
rect 12497 -5662 12544 -5598
rect 12608 -5662 12624 -5598
rect 12497 -5678 12624 -5662
rect 12497 -5742 12544 -5678
rect 12608 -5742 12624 -5678
rect 12497 -5758 12624 -5742
rect 12497 -5822 12544 -5758
rect 12608 -5822 12624 -5758
rect 12497 -5838 12624 -5822
rect 12497 -5902 12544 -5838
rect 12608 -5902 12624 -5838
rect 12497 -5918 12624 -5902
rect 12497 -5982 12544 -5918
rect 12608 -5982 12624 -5918
rect 12497 -5998 12624 -5982
rect 12497 -6062 12544 -5998
rect 12608 -6062 12624 -5998
rect 12497 -6078 12624 -6062
rect 6178 -6158 6305 -6142
rect 6178 -6222 6225 -6158
rect 6289 -6222 6305 -6158
rect 6178 -6238 6305 -6222
rect 6178 -6362 6282 -6238
rect 6178 -6378 6305 -6362
rect 6178 -6442 6225 -6378
rect 6289 -6442 6305 -6378
rect 6178 -6458 6305 -6442
rect -141 -6538 -14 -6522
rect -141 -6602 -94 -6538
rect -30 -6602 -14 -6538
rect -141 -6618 -14 -6602
rect -141 -6682 -94 -6618
rect -30 -6682 -14 -6618
rect -141 -6698 -14 -6682
rect -141 -6762 -94 -6698
rect -30 -6762 -14 -6698
rect -141 -6778 -14 -6762
rect -141 -6842 -94 -6778
rect -30 -6842 -14 -6778
rect -141 -6858 -14 -6842
rect -141 -6922 -94 -6858
rect -30 -6922 -14 -6858
rect -141 -6938 -14 -6922
rect -141 -7002 -94 -6938
rect -30 -7002 -14 -6938
rect -141 -7018 -14 -7002
rect -141 -7082 -94 -7018
rect -30 -7082 -14 -7018
rect -141 -7098 -14 -7082
rect -141 -7162 -94 -7098
rect -30 -7162 -14 -7098
rect -141 -7178 -14 -7162
rect -141 -7242 -94 -7178
rect -30 -7242 -14 -7178
rect -141 -7258 -14 -7242
rect -141 -7322 -94 -7258
rect -30 -7322 -14 -7258
rect -141 -7338 -14 -7322
rect -141 -7402 -94 -7338
rect -30 -7402 -14 -7338
rect -141 -7418 -14 -7402
rect -141 -7482 -94 -7418
rect -30 -7482 -14 -7418
rect -141 -7498 -14 -7482
rect -141 -7562 -94 -7498
rect -30 -7562 -14 -7498
rect -141 -7578 -14 -7562
rect -141 -7642 -94 -7578
rect -30 -7642 -14 -7578
rect -141 -7658 -14 -7642
rect -141 -7722 -94 -7658
rect -30 -7722 -14 -7658
rect -141 -7738 -14 -7722
rect -141 -7802 -94 -7738
rect -30 -7802 -14 -7738
rect -141 -7818 -14 -7802
rect -141 -7882 -94 -7818
rect -30 -7882 -14 -7818
rect -141 -7898 -14 -7882
rect -141 -7962 -94 -7898
rect -30 -7962 -14 -7898
rect -141 -7978 -14 -7962
rect -141 -8042 -94 -7978
rect -30 -8042 -14 -7978
rect -141 -8058 -14 -8042
rect -141 -8122 -94 -8058
rect -30 -8122 -14 -8058
rect -141 -8138 -14 -8122
rect -141 -8202 -94 -8138
rect -30 -8202 -14 -8138
rect -141 -8218 -14 -8202
rect -141 -8282 -94 -8218
rect -30 -8282 -14 -8218
rect -141 -8298 -14 -8282
rect -141 -8362 -94 -8298
rect -30 -8362 -14 -8298
rect -141 -8378 -14 -8362
rect -141 -8442 -94 -8378
rect -30 -8442 -14 -8378
rect -141 -8458 -14 -8442
rect -141 -8522 -94 -8458
rect -30 -8522 -14 -8458
rect -141 -8538 -14 -8522
rect -141 -8602 -94 -8538
rect -30 -8602 -14 -8538
rect -141 -8618 -14 -8602
rect -141 -8682 -94 -8618
rect -30 -8682 -14 -8618
rect -141 -8698 -14 -8682
rect -141 -8762 -94 -8698
rect -30 -8762 -14 -8698
rect -141 -8778 -14 -8762
rect -141 -8842 -94 -8778
rect -30 -8842 -14 -8778
rect -141 -8858 -14 -8842
rect -141 -8922 -94 -8858
rect -30 -8922 -14 -8858
rect -141 -8938 -14 -8922
rect -141 -9002 -94 -8938
rect -30 -9002 -14 -8938
rect -141 -9018 -14 -9002
rect -141 -9082 -94 -9018
rect -30 -9082 -14 -9018
rect -141 -9098 -14 -9082
rect -141 -9162 -94 -9098
rect -30 -9162 -14 -9098
rect -141 -9178 -14 -9162
rect -141 -9242 -94 -9178
rect -30 -9242 -14 -9178
rect -141 -9258 -14 -9242
rect -141 -9322 -94 -9258
rect -30 -9322 -14 -9258
rect -141 -9338 -14 -9322
rect -141 -9402 -94 -9338
rect -30 -9402 -14 -9338
rect -141 -9418 -14 -9402
rect -141 -9482 -94 -9418
rect -30 -9482 -14 -9418
rect -141 -9498 -14 -9482
rect -141 -9562 -94 -9498
rect -30 -9562 -14 -9498
rect -141 -9578 -14 -9562
rect -141 -9642 -94 -9578
rect -30 -9642 -14 -9578
rect -141 -9658 -14 -9642
rect -141 -9722 -94 -9658
rect -30 -9722 -14 -9658
rect -141 -9738 -14 -9722
rect -141 -9802 -94 -9738
rect -30 -9802 -14 -9738
rect -141 -9818 -14 -9802
rect -141 -9882 -94 -9818
rect -30 -9882 -14 -9818
rect -141 -9898 -14 -9882
rect -141 -9962 -94 -9898
rect -30 -9962 -14 -9898
rect -141 -9978 -14 -9962
rect -141 -10042 -94 -9978
rect -30 -10042 -14 -9978
rect -141 -10058 -14 -10042
rect -141 -10122 -94 -10058
rect -30 -10122 -14 -10058
rect -141 -10138 -14 -10122
rect -141 -10202 -94 -10138
rect -30 -10202 -14 -10138
rect -141 -10218 -14 -10202
rect -141 -10282 -94 -10218
rect -30 -10282 -14 -10218
rect -141 -10298 -14 -10282
rect -141 -10362 -94 -10298
rect -30 -10362 -14 -10298
rect -141 -10378 -14 -10362
rect -141 -10442 -94 -10378
rect -30 -10442 -14 -10378
rect -141 -10458 -14 -10442
rect -141 -10522 -94 -10458
rect -30 -10522 -14 -10458
rect -141 -10538 -14 -10522
rect -141 -10602 -94 -10538
rect -30 -10602 -14 -10538
rect -141 -10618 -14 -10602
rect -141 -10682 -94 -10618
rect -30 -10682 -14 -10618
rect -141 -10698 -14 -10682
rect -141 -10762 -94 -10698
rect -30 -10762 -14 -10698
rect -141 -10778 -14 -10762
rect -141 -10842 -94 -10778
rect -30 -10842 -14 -10778
rect -141 -10858 -14 -10842
rect -141 -10922 -94 -10858
rect -30 -10922 -14 -10858
rect -141 -10938 -14 -10922
rect -141 -11002 -94 -10938
rect -30 -11002 -14 -10938
rect -141 -11018 -14 -11002
rect -141 -11082 -94 -11018
rect -30 -11082 -14 -11018
rect -141 -11098 -14 -11082
rect -141 -11162 -94 -11098
rect -30 -11162 -14 -11098
rect -141 -11178 -14 -11162
rect -141 -11242 -94 -11178
rect -30 -11242 -14 -11178
rect -141 -11258 -14 -11242
rect -141 -11322 -94 -11258
rect -30 -11322 -14 -11258
rect -141 -11338 -14 -11322
rect -141 -11402 -94 -11338
rect -30 -11402 -14 -11338
rect -141 -11418 -14 -11402
rect -141 -11482 -94 -11418
rect -30 -11482 -14 -11418
rect -141 -11498 -14 -11482
rect -141 -11562 -94 -11498
rect -30 -11562 -14 -11498
rect -141 -11578 -14 -11562
rect -141 -11642 -94 -11578
rect -30 -11642 -14 -11578
rect -141 -11658 -14 -11642
rect -141 -11722 -94 -11658
rect -30 -11722 -14 -11658
rect -141 -11738 -14 -11722
rect -141 -11802 -94 -11738
rect -30 -11802 -14 -11738
rect -141 -11818 -14 -11802
rect -141 -11882 -94 -11818
rect -30 -11882 -14 -11818
rect -141 -11898 -14 -11882
rect -141 -11962 -94 -11898
rect -30 -11962 -14 -11898
rect -141 -11978 -14 -11962
rect -141 -12042 -94 -11978
rect -30 -12042 -14 -11978
rect -141 -12058 -14 -12042
rect -141 -12122 -94 -12058
rect -30 -12122 -14 -12058
rect -141 -12138 -14 -12122
rect -141 -12202 -94 -12138
rect -30 -12202 -14 -12138
rect -141 -12218 -14 -12202
rect -141 -12282 -94 -12218
rect -30 -12282 -14 -12218
rect -141 -12298 -14 -12282
rect -141 -12362 -94 -12298
rect -30 -12362 -14 -12298
rect -141 -12378 -14 -12362
rect -6460 -12458 -6333 -12442
rect -6460 -12522 -6413 -12458
rect -6349 -12522 -6333 -12458
rect -6460 -12538 -6333 -12522
rect -6460 -12600 -6356 -12538
rect -3261 -12600 -3157 -12411
rect -141 -12442 -94 -12378
rect -30 -12442 -14 -12378
rect 149 -6498 6071 -6489
rect 149 -12402 158 -6498
rect 6062 -12402 6071 -6498
rect 149 -12411 6071 -12402
rect 6178 -6522 6225 -6458
rect 6289 -6522 6305 -6458
rect 9377 -6489 9481 -6111
rect 12497 -6142 12544 -6078
rect 12608 -6142 12624 -6078
rect 12497 -6158 12624 -6142
rect 12497 -6222 12544 -6158
rect 12608 -6222 12624 -6158
rect 12497 -6238 12624 -6222
rect 12497 -6362 12601 -6238
rect 12497 -6378 12624 -6362
rect 12497 -6442 12544 -6378
rect 12608 -6442 12624 -6378
rect 12497 -6458 12624 -6442
rect 6178 -6538 6305 -6522
rect 6178 -6602 6225 -6538
rect 6289 -6602 6305 -6538
rect 6178 -6618 6305 -6602
rect 6178 -6682 6225 -6618
rect 6289 -6682 6305 -6618
rect 6178 -6698 6305 -6682
rect 6178 -6762 6225 -6698
rect 6289 -6762 6305 -6698
rect 6178 -6778 6305 -6762
rect 6178 -6842 6225 -6778
rect 6289 -6842 6305 -6778
rect 6178 -6858 6305 -6842
rect 6178 -6922 6225 -6858
rect 6289 -6922 6305 -6858
rect 6178 -6938 6305 -6922
rect 6178 -7002 6225 -6938
rect 6289 -7002 6305 -6938
rect 6178 -7018 6305 -7002
rect 6178 -7082 6225 -7018
rect 6289 -7082 6305 -7018
rect 6178 -7098 6305 -7082
rect 6178 -7162 6225 -7098
rect 6289 -7162 6305 -7098
rect 6178 -7178 6305 -7162
rect 6178 -7242 6225 -7178
rect 6289 -7242 6305 -7178
rect 6178 -7258 6305 -7242
rect 6178 -7322 6225 -7258
rect 6289 -7322 6305 -7258
rect 6178 -7338 6305 -7322
rect 6178 -7402 6225 -7338
rect 6289 -7402 6305 -7338
rect 6178 -7418 6305 -7402
rect 6178 -7482 6225 -7418
rect 6289 -7482 6305 -7418
rect 6178 -7498 6305 -7482
rect 6178 -7562 6225 -7498
rect 6289 -7562 6305 -7498
rect 6178 -7578 6305 -7562
rect 6178 -7642 6225 -7578
rect 6289 -7642 6305 -7578
rect 6178 -7658 6305 -7642
rect 6178 -7722 6225 -7658
rect 6289 -7722 6305 -7658
rect 6178 -7738 6305 -7722
rect 6178 -7802 6225 -7738
rect 6289 -7802 6305 -7738
rect 6178 -7818 6305 -7802
rect 6178 -7882 6225 -7818
rect 6289 -7882 6305 -7818
rect 6178 -7898 6305 -7882
rect 6178 -7962 6225 -7898
rect 6289 -7962 6305 -7898
rect 6178 -7978 6305 -7962
rect 6178 -8042 6225 -7978
rect 6289 -8042 6305 -7978
rect 6178 -8058 6305 -8042
rect 6178 -8122 6225 -8058
rect 6289 -8122 6305 -8058
rect 6178 -8138 6305 -8122
rect 6178 -8202 6225 -8138
rect 6289 -8202 6305 -8138
rect 6178 -8218 6305 -8202
rect 6178 -8282 6225 -8218
rect 6289 -8282 6305 -8218
rect 6178 -8298 6305 -8282
rect 6178 -8362 6225 -8298
rect 6289 -8362 6305 -8298
rect 6178 -8378 6305 -8362
rect 6178 -8442 6225 -8378
rect 6289 -8442 6305 -8378
rect 6178 -8458 6305 -8442
rect 6178 -8522 6225 -8458
rect 6289 -8522 6305 -8458
rect 6178 -8538 6305 -8522
rect 6178 -8602 6225 -8538
rect 6289 -8602 6305 -8538
rect 6178 -8618 6305 -8602
rect 6178 -8682 6225 -8618
rect 6289 -8682 6305 -8618
rect 6178 -8698 6305 -8682
rect 6178 -8762 6225 -8698
rect 6289 -8762 6305 -8698
rect 6178 -8778 6305 -8762
rect 6178 -8842 6225 -8778
rect 6289 -8842 6305 -8778
rect 6178 -8858 6305 -8842
rect 6178 -8922 6225 -8858
rect 6289 -8922 6305 -8858
rect 6178 -8938 6305 -8922
rect 6178 -9002 6225 -8938
rect 6289 -9002 6305 -8938
rect 6178 -9018 6305 -9002
rect 6178 -9082 6225 -9018
rect 6289 -9082 6305 -9018
rect 6178 -9098 6305 -9082
rect 6178 -9162 6225 -9098
rect 6289 -9162 6305 -9098
rect 6178 -9178 6305 -9162
rect 6178 -9242 6225 -9178
rect 6289 -9242 6305 -9178
rect 6178 -9258 6305 -9242
rect 6178 -9322 6225 -9258
rect 6289 -9322 6305 -9258
rect 6178 -9338 6305 -9322
rect 6178 -9402 6225 -9338
rect 6289 -9402 6305 -9338
rect 6178 -9418 6305 -9402
rect 6178 -9482 6225 -9418
rect 6289 -9482 6305 -9418
rect 6178 -9498 6305 -9482
rect 6178 -9562 6225 -9498
rect 6289 -9562 6305 -9498
rect 6178 -9578 6305 -9562
rect 6178 -9642 6225 -9578
rect 6289 -9642 6305 -9578
rect 6178 -9658 6305 -9642
rect 6178 -9722 6225 -9658
rect 6289 -9722 6305 -9658
rect 6178 -9738 6305 -9722
rect 6178 -9802 6225 -9738
rect 6289 -9802 6305 -9738
rect 6178 -9818 6305 -9802
rect 6178 -9882 6225 -9818
rect 6289 -9882 6305 -9818
rect 6178 -9898 6305 -9882
rect 6178 -9962 6225 -9898
rect 6289 -9962 6305 -9898
rect 6178 -9978 6305 -9962
rect 6178 -10042 6225 -9978
rect 6289 -10042 6305 -9978
rect 6178 -10058 6305 -10042
rect 6178 -10122 6225 -10058
rect 6289 -10122 6305 -10058
rect 6178 -10138 6305 -10122
rect 6178 -10202 6225 -10138
rect 6289 -10202 6305 -10138
rect 6178 -10218 6305 -10202
rect 6178 -10282 6225 -10218
rect 6289 -10282 6305 -10218
rect 6178 -10298 6305 -10282
rect 6178 -10362 6225 -10298
rect 6289 -10362 6305 -10298
rect 6178 -10378 6305 -10362
rect 6178 -10442 6225 -10378
rect 6289 -10442 6305 -10378
rect 6178 -10458 6305 -10442
rect 6178 -10522 6225 -10458
rect 6289 -10522 6305 -10458
rect 6178 -10538 6305 -10522
rect 6178 -10602 6225 -10538
rect 6289 -10602 6305 -10538
rect 6178 -10618 6305 -10602
rect 6178 -10682 6225 -10618
rect 6289 -10682 6305 -10618
rect 6178 -10698 6305 -10682
rect 6178 -10762 6225 -10698
rect 6289 -10762 6305 -10698
rect 6178 -10778 6305 -10762
rect 6178 -10842 6225 -10778
rect 6289 -10842 6305 -10778
rect 6178 -10858 6305 -10842
rect 6178 -10922 6225 -10858
rect 6289 -10922 6305 -10858
rect 6178 -10938 6305 -10922
rect 6178 -11002 6225 -10938
rect 6289 -11002 6305 -10938
rect 6178 -11018 6305 -11002
rect 6178 -11082 6225 -11018
rect 6289 -11082 6305 -11018
rect 6178 -11098 6305 -11082
rect 6178 -11162 6225 -11098
rect 6289 -11162 6305 -11098
rect 6178 -11178 6305 -11162
rect 6178 -11242 6225 -11178
rect 6289 -11242 6305 -11178
rect 6178 -11258 6305 -11242
rect 6178 -11322 6225 -11258
rect 6289 -11322 6305 -11258
rect 6178 -11338 6305 -11322
rect 6178 -11402 6225 -11338
rect 6289 -11402 6305 -11338
rect 6178 -11418 6305 -11402
rect 6178 -11482 6225 -11418
rect 6289 -11482 6305 -11418
rect 6178 -11498 6305 -11482
rect 6178 -11562 6225 -11498
rect 6289 -11562 6305 -11498
rect 6178 -11578 6305 -11562
rect 6178 -11642 6225 -11578
rect 6289 -11642 6305 -11578
rect 6178 -11658 6305 -11642
rect 6178 -11722 6225 -11658
rect 6289 -11722 6305 -11658
rect 6178 -11738 6305 -11722
rect 6178 -11802 6225 -11738
rect 6289 -11802 6305 -11738
rect 6178 -11818 6305 -11802
rect 6178 -11882 6225 -11818
rect 6289 -11882 6305 -11818
rect 6178 -11898 6305 -11882
rect 6178 -11962 6225 -11898
rect 6289 -11962 6305 -11898
rect 6178 -11978 6305 -11962
rect 6178 -12042 6225 -11978
rect 6289 -12042 6305 -11978
rect 6178 -12058 6305 -12042
rect 6178 -12122 6225 -12058
rect 6289 -12122 6305 -12058
rect 6178 -12138 6305 -12122
rect 6178 -12202 6225 -12138
rect 6289 -12202 6305 -12138
rect 6178 -12218 6305 -12202
rect 6178 -12282 6225 -12218
rect 6289 -12282 6305 -12218
rect 6178 -12298 6305 -12282
rect 6178 -12362 6225 -12298
rect 6289 -12362 6305 -12298
rect 6178 -12378 6305 -12362
rect -141 -12458 -14 -12442
rect -141 -12522 -94 -12458
rect -30 -12522 -14 -12458
rect -141 -12538 -14 -12522
rect -141 -12600 -37 -12538
rect 3058 -12600 3162 -12411
rect 6178 -12442 6225 -12378
rect 6289 -12442 6305 -12378
rect 6468 -6498 12390 -6489
rect 6468 -12402 6477 -6498
rect 12381 -12402 12390 -6498
rect 6468 -12411 12390 -12402
rect 12497 -6522 12544 -6458
rect 12608 -6522 12624 -6458
rect 12497 -6538 12624 -6522
rect 12497 -6602 12544 -6538
rect 12608 -6602 12624 -6538
rect 12497 -6618 12624 -6602
rect 12497 -6682 12544 -6618
rect 12608 -6682 12624 -6618
rect 12497 -6698 12624 -6682
rect 12497 -6762 12544 -6698
rect 12608 -6762 12624 -6698
rect 12497 -6778 12624 -6762
rect 12497 -6842 12544 -6778
rect 12608 -6842 12624 -6778
rect 12497 -6858 12624 -6842
rect 12497 -6922 12544 -6858
rect 12608 -6922 12624 -6858
rect 12497 -6938 12624 -6922
rect 12497 -7002 12544 -6938
rect 12608 -7002 12624 -6938
rect 12497 -7018 12624 -7002
rect 12497 -7082 12544 -7018
rect 12608 -7082 12624 -7018
rect 12497 -7098 12624 -7082
rect 12497 -7162 12544 -7098
rect 12608 -7162 12624 -7098
rect 12497 -7178 12624 -7162
rect 12497 -7242 12544 -7178
rect 12608 -7242 12624 -7178
rect 12497 -7258 12624 -7242
rect 12497 -7322 12544 -7258
rect 12608 -7322 12624 -7258
rect 12497 -7338 12624 -7322
rect 12497 -7402 12544 -7338
rect 12608 -7402 12624 -7338
rect 12497 -7418 12624 -7402
rect 12497 -7482 12544 -7418
rect 12608 -7482 12624 -7418
rect 12497 -7498 12624 -7482
rect 12497 -7562 12544 -7498
rect 12608 -7562 12624 -7498
rect 12497 -7578 12624 -7562
rect 12497 -7642 12544 -7578
rect 12608 -7642 12624 -7578
rect 12497 -7658 12624 -7642
rect 12497 -7722 12544 -7658
rect 12608 -7722 12624 -7658
rect 12497 -7738 12624 -7722
rect 12497 -7802 12544 -7738
rect 12608 -7802 12624 -7738
rect 12497 -7818 12624 -7802
rect 12497 -7882 12544 -7818
rect 12608 -7882 12624 -7818
rect 12497 -7898 12624 -7882
rect 12497 -7962 12544 -7898
rect 12608 -7962 12624 -7898
rect 12497 -7978 12624 -7962
rect 12497 -8042 12544 -7978
rect 12608 -8042 12624 -7978
rect 12497 -8058 12624 -8042
rect 12497 -8122 12544 -8058
rect 12608 -8122 12624 -8058
rect 12497 -8138 12624 -8122
rect 12497 -8202 12544 -8138
rect 12608 -8202 12624 -8138
rect 12497 -8218 12624 -8202
rect 12497 -8282 12544 -8218
rect 12608 -8282 12624 -8218
rect 12497 -8298 12624 -8282
rect 12497 -8362 12544 -8298
rect 12608 -8362 12624 -8298
rect 12497 -8378 12624 -8362
rect 12497 -8442 12544 -8378
rect 12608 -8442 12624 -8378
rect 12497 -8458 12624 -8442
rect 12497 -8522 12544 -8458
rect 12608 -8522 12624 -8458
rect 12497 -8538 12624 -8522
rect 12497 -8602 12544 -8538
rect 12608 -8602 12624 -8538
rect 12497 -8618 12624 -8602
rect 12497 -8682 12544 -8618
rect 12608 -8682 12624 -8618
rect 12497 -8698 12624 -8682
rect 12497 -8762 12544 -8698
rect 12608 -8762 12624 -8698
rect 12497 -8778 12624 -8762
rect 12497 -8842 12544 -8778
rect 12608 -8842 12624 -8778
rect 12497 -8858 12624 -8842
rect 12497 -8922 12544 -8858
rect 12608 -8922 12624 -8858
rect 12497 -8938 12624 -8922
rect 12497 -9002 12544 -8938
rect 12608 -9002 12624 -8938
rect 12497 -9018 12624 -9002
rect 12497 -9082 12544 -9018
rect 12608 -9082 12624 -9018
rect 12497 -9098 12624 -9082
rect 12497 -9162 12544 -9098
rect 12608 -9162 12624 -9098
rect 12497 -9178 12624 -9162
rect 12497 -9242 12544 -9178
rect 12608 -9242 12624 -9178
rect 12497 -9258 12624 -9242
rect 12497 -9322 12544 -9258
rect 12608 -9322 12624 -9258
rect 12497 -9338 12624 -9322
rect 12497 -9402 12544 -9338
rect 12608 -9402 12624 -9338
rect 12497 -9418 12624 -9402
rect 12497 -9482 12544 -9418
rect 12608 -9482 12624 -9418
rect 12497 -9498 12624 -9482
rect 12497 -9562 12544 -9498
rect 12608 -9562 12624 -9498
rect 12497 -9578 12624 -9562
rect 12497 -9642 12544 -9578
rect 12608 -9642 12624 -9578
rect 12497 -9658 12624 -9642
rect 12497 -9722 12544 -9658
rect 12608 -9722 12624 -9658
rect 12497 -9738 12624 -9722
rect 12497 -9802 12544 -9738
rect 12608 -9802 12624 -9738
rect 12497 -9818 12624 -9802
rect 12497 -9882 12544 -9818
rect 12608 -9882 12624 -9818
rect 12497 -9898 12624 -9882
rect 12497 -9962 12544 -9898
rect 12608 -9962 12624 -9898
rect 12497 -9978 12624 -9962
rect 12497 -10042 12544 -9978
rect 12608 -10042 12624 -9978
rect 12497 -10058 12624 -10042
rect 12497 -10122 12544 -10058
rect 12608 -10122 12624 -10058
rect 12497 -10138 12624 -10122
rect 12497 -10202 12544 -10138
rect 12608 -10202 12624 -10138
rect 12497 -10218 12624 -10202
rect 12497 -10282 12544 -10218
rect 12608 -10282 12624 -10218
rect 12497 -10298 12624 -10282
rect 12497 -10362 12544 -10298
rect 12608 -10362 12624 -10298
rect 12497 -10378 12624 -10362
rect 12497 -10442 12544 -10378
rect 12608 -10442 12624 -10378
rect 12497 -10458 12624 -10442
rect 12497 -10522 12544 -10458
rect 12608 -10522 12624 -10458
rect 12497 -10538 12624 -10522
rect 12497 -10602 12544 -10538
rect 12608 -10602 12624 -10538
rect 12497 -10618 12624 -10602
rect 12497 -10682 12544 -10618
rect 12608 -10682 12624 -10618
rect 12497 -10698 12624 -10682
rect 12497 -10762 12544 -10698
rect 12608 -10762 12624 -10698
rect 12497 -10778 12624 -10762
rect 12497 -10842 12544 -10778
rect 12608 -10842 12624 -10778
rect 12497 -10858 12624 -10842
rect 12497 -10922 12544 -10858
rect 12608 -10922 12624 -10858
rect 12497 -10938 12624 -10922
rect 12497 -11002 12544 -10938
rect 12608 -11002 12624 -10938
rect 12497 -11018 12624 -11002
rect 12497 -11082 12544 -11018
rect 12608 -11082 12624 -11018
rect 12497 -11098 12624 -11082
rect 12497 -11162 12544 -11098
rect 12608 -11162 12624 -11098
rect 12497 -11178 12624 -11162
rect 12497 -11242 12544 -11178
rect 12608 -11242 12624 -11178
rect 12497 -11258 12624 -11242
rect 12497 -11322 12544 -11258
rect 12608 -11322 12624 -11258
rect 12497 -11338 12624 -11322
rect 12497 -11402 12544 -11338
rect 12608 -11402 12624 -11338
rect 12497 -11418 12624 -11402
rect 12497 -11482 12544 -11418
rect 12608 -11482 12624 -11418
rect 12497 -11498 12624 -11482
rect 12497 -11562 12544 -11498
rect 12608 -11562 12624 -11498
rect 12497 -11578 12624 -11562
rect 12497 -11642 12544 -11578
rect 12608 -11642 12624 -11578
rect 12497 -11658 12624 -11642
rect 12497 -11722 12544 -11658
rect 12608 -11722 12624 -11658
rect 12497 -11738 12624 -11722
rect 12497 -11802 12544 -11738
rect 12608 -11802 12624 -11738
rect 12497 -11818 12624 -11802
rect 12497 -11882 12544 -11818
rect 12608 -11882 12624 -11818
rect 12497 -11898 12624 -11882
rect 12497 -11962 12544 -11898
rect 12608 -11962 12624 -11898
rect 12497 -11978 12624 -11962
rect 12497 -12042 12544 -11978
rect 12608 -12042 12624 -11978
rect 12497 -12058 12624 -12042
rect 12497 -12122 12544 -12058
rect 12608 -12122 12624 -12058
rect 12497 -12138 12624 -12122
rect 12497 -12202 12544 -12138
rect 12608 -12202 12624 -12138
rect 12497 -12218 12624 -12202
rect 12497 -12282 12544 -12218
rect 12608 -12282 12624 -12218
rect 12497 -12298 12624 -12282
rect 12497 -12362 12544 -12298
rect 12608 -12362 12624 -12298
rect 12497 -12378 12624 -12362
rect 6178 -12458 6305 -12442
rect 6178 -12522 6225 -12458
rect 6289 -12522 6305 -12458
rect 6178 -12538 6305 -12522
rect 6178 -12600 6282 -12538
rect 9377 -12600 9481 -12411
rect 12497 -12442 12544 -12378
rect 12608 -12442 12624 -12378
rect 12497 -12458 12624 -12442
rect 12497 -12522 12544 -12458
rect 12608 -12522 12624 -12458
rect 12497 -12538 12624 -12522
rect 12497 -12600 12601 -12538
<< properties >>
string FIXED_BBOX 6329 6350 12529 12550
<< end >>
