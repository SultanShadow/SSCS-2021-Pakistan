magic
tech sky130A
timestamp 1635939177
<< nwell >>
rect -269 -269 269 269
<< pwell >>
rect -338 269 338 338
rect -338 -269 -269 269
rect 269 -269 338 269
rect -338 -338 338 -269
<< psubdiff >>
rect -320 303 -272 320
rect 272 303 320 320
rect -320 272 -303 303
rect 303 272 320 303
rect -320 -303 -303 -272
rect 303 -303 320 -272
rect -320 -320 -272 -303
rect 272 -320 320 -303
<< nsubdiff >>
rect -251 234 -203 251
rect 203 234 251 251
rect -251 203 -234 234
rect 234 203 251 234
rect -251 -234 -234 -203
rect 234 -234 251 -203
rect -251 -251 -203 -234
rect 203 -251 251 -234
<< psubdiffcont >>
rect -272 303 272 320
rect -320 -272 -303 272
rect 303 -272 320 272
rect -272 -320 272 -303
<< nsubdiffcont >>
rect -203 234 203 251
rect -251 -203 -234 203
rect 234 -203 251 203
rect -203 -251 203 -234
<< pdiode >>
rect -200 194 200 200
rect -200 -194 -194 194
rect 194 -194 200 194
rect -200 -200 200 -194
<< pdiodec >>
rect -194 -194 194 194
<< locali >>
rect -320 303 -272 320
rect 272 303 320 320
rect -320 272 -303 303
rect 303 272 320 303
rect -251 234 -203 251
rect 203 234 251 251
rect -251 203 -234 234
rect 234 203 251 234
rect -202 -194 -194 194
rect 194 -194 202 194
rect -251 -234 -234 -203
rect 234 -234 251 -203
rect -251 -251 -203 -234
rect 203 -251 251 -234
rect -320 -303 -303 -272
rect 303 -303 320 -272
rect -320 -320 -272 -303
rect 272 -320 320 -303
<< viali >>
rect -194 -194 194 194
<< metal1 >>
rect -200 194 200 197
rect -200 -194 -194 194
rect 194 -194 200 194
rect -200 -197 200 -194
<< properties >>
string gencell sky130_fd_pr__diode_pd2nw_05v5
string FIXED_BBOX -242 -242 242 242
string parameters w 4 l 4 area 16.0 peri 16.0 nx 1 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 glc 1 grc 1 gtc 1 gbc 1 doverlap 0 compatible {sky130_fd_pr__diode_pd2nw_05v5 sky130_fd_pr__diode_pd2nw_05v5_lvt  sky130_fd_pr__diode_pd2nw_05v5_hvt sky130_fd_pr__diode_pd2nw_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
string library sky130
<< end >>
